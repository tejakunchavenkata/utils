g7.sv