class board;
  typedef enum {
    AAA=1,
    AAB=2,
    AAC=3,
    AAD=4,
    AAE=5,
    AAF=6,
    AAG=7,
    AAH=8,
    AAI=9,
    AAJ=10,
    AAK=11,
    AAL=12,
    AAM=13,
    AAN=14,
    AAO=15,
    AAP=16,
    AAQ=17,
    AAR=18,
    AAS=19,
    AAT=20,
    AAU=21,
    AAV=22,
    AAW=23,
    AAX=24,
    AAY
  } elements;
  rand elements ele[25][25];
  constraint all {
    ele[0][0] != ele[0][1];
    ele[0][0] != ele[0][10];
    ele[0][0] != ele[0][11];
    ele[0][0] != ele[0][12];
    ele[0][0] != ele[0][13];
    ele[0][0] != ele[0][14];
    ele[0][0] != ele[0][15];
    ele[0][0] != ele[0][16];
    ele[0][0] != ele[0][17];
    ele[0][0] != ele[0][18];
    ele[0][0] != ele[0][19];
    ele[0][0] != ele[0][2];
    ele[0][0] != ele[0][20];
    ele[0][0] != ele[0][21];
    ele[0][0] != ele[0][22];
    ele[0][0] != ele[0][23];
    ele[0][0] != ele[0][24];
    ele[0][0] != ele[0][3];
    ele[0][0] != ele[0][4];
    ele[0][0] != ele[0][5];
    ele[0][0] != ele[0][6];
    ele[0][0] != ele[0][7];
    ele[0][0] != ele[0][8];
    ele[0][0] != ele[0][9];
    ele[0][0] != ele[1][0];
    ele[0][0] != ele[1][1];
    ele[0][0] != ele[1][2];
    ele[0][0] != ele[1][3];
    ele[0][0] != ele[1][4];
    ele[0][0] != ele[10][0];
    ele[0][0] != ele[11][0];
    ele[0][0] != ele[12][0];
    ele[0][0] != ele[13][0];
    ele[0][0] != ele[14][0];
    ele[0][0] != ele[15][0];
    ele[0][0] != ele[16][0];
    ele[0][0] != ele[17][0];
    ele[0][0] != ele[18][0];
    ele[0][0] != ele[19][0];
    ele[0][0] != ele[2][0];
    ele[0][0] != ele[2][1];
    ele[0][0] != ele[2][2];
    ele[0][0] != ele[2][3];
    ele[0][0] != ele[2][4];
    ele[0][0] != ele[20][0];
    ele[0][0] != ele[21][0];
    ele[0][0] != ele[22][0];
    ele[0][0] != ele[23][0];
    ele[0][0] != ele[24][0];
    ele[0][0] != ele[3][0];
    ele[0][0] != ele[3][1];
    ele[0][0] != ele[3][2];
    ele[0][0] != ele[3][3];
    ele[0][0] != ele[3][4];
    ele[0][0] != ele[4][0];
    ele[0][0] != ele[4][1];
    ele[0][0] != ele[4][2];
    ele[0][0] != ele[4][3];
    ele[0][0] != ele[4][4];
    ele[0][0] != ele[5][0];
    ele[0][0] != ele[6][0];
    ele[0][0] != ele[7][0];
    ele[0][0] != ele[8][0];
    ele[0][0] != ele[9][0];
    ele[0][1] != ele[0][10];
    ele[0][1] != ele[0][11];
    ele[0][1] != ele[0][12];
    ele[0][1] != ele[0][13];
    ele[0][1] != ele[0][14];
    ele[0][1] != ele[0][15];
    ele[0][1] != ele[0][16];
    ele[0][1] != ele[0][17];
    ele[0][1] != ele[0][18];
    ele[0][1] != ele[0][19];
    ele[0][1] != ele[0][2];
    ele[0][1] != ele[0][20];
    ele[0][1] != ele[0][21];
    ele[0][1] != ele[0][22];
    ele[0][1] != ele[0][23];
    ele[0][1] != ele[0][24];
    ele[0][1] != ele[0][3];
    ele[0][1] != ele[0][4];
    ele[0][1] != ele[0][5];
    ele[0][1] != ele[0][6];
    ele[0][1] != ele[0][7];
    ele[0][1] != ele[0][8];
    ele[0][1] != ele[0][9];
    ele[0][1] != ele[1][0];
    ele[0][1] != ele[1][1];
    ele[0][1] != ele[1][2];
    ele[0][1] != ele[1][3];
    ele[0][1] != ele[1][4];
    ele[0][1] != ele[10][1];
    ele[0][1] != ele[11][1];
    ele[0][1] != ele[12][1];
    ele[0][1] != ele[13][1];
    ele[0][1] != ele[14][1];
    ele[0][1] != ele[15][1];
    ele[0][1] != ele[16][1];
    ele[0][1] != ele[17][1];
    ele[0][1] != ele[18][1];
    ele[0][1] != ele[19][1];
    ele[0][1] != ele[2][0];
    ele[0][1] != ele[2][1];
    ele[0][1] != ele[2][2];
    ele[0][1] != ele[2][3];
    ele[0][1] != ele[2][4];
    ele[0][1] != ele[20][1];
    ele[0][1] != ele[21][1];
    ele[0][1] != ele[22][1];
    ele[0][1] != ele[23][1];
    ele[0][1] != ele[24][1];
    ele[0][1] != ele[3][0];
    ele[0][1] != ele[3][1];
    ele[0][1] != ele[3][2];
    ele[0][1] != ele[3][3];
    ele[0][1] != ele[3][4];
    ele[0][1] != ele[4][0];
    ele[0][1] != ele[4][1];
    ele[0][1] != ele[4][2];
    ele[0][1] != ele[4][3];
    ele[0][1] != ele[4][4];
    ele[0][1] != ele[5][1];
    ele[0][1] != ele[6][1];
    ele[0][1] != ele[7][1];
    ele[0][1] != ele[8][1];
    ele[0][1] != ele[9][1];
    ele[0][10] != ele[0][11];
    ele[0][10] != ele[0][12];
    ele[0][10] != ele[0][13];
    ele[0][10] != ele[0][14];
    ele[0][10] != ele[0][15];
    ele[0][10] != ele[0][16];
    ele[0][10] != ele[0][17];
    ele[0][10] != ele[0][18];
    ele[0][10] != ele[0][19];
    ele[0][10] != ele[0][20];
    ele[0][10] != ele[0][21];
    ele[0][10] != ele[0][22];
    ele[0][10] != ele[0][23];
    ele[0][10] != ele[0][24];
    ele[0][10] != ele[1][10];
    ele[0][10] != ele[1][11];
    ele[0][10] != ele[1][12];
    ele[0][10] != ele[1][13];
    ele[0][10] != ele[1][14];
    ele[0][10] != ele[10][10];
    ele[0][10] != ele[11][10];
    ele[0][10] != ele[12][10];
    ele[0][10] != ele[13][10];
    ele[0][10] != ele[14][10];
    ele[0][10] != ele[15][10];
    ele[0][10] != ele[16][10];
    ele[0][10] != ele[17][10];
    ele[0][10] != ele[18][10];
    ele[0][10] != ele[19][10];
    ele[0][10] != ele[2][10];
    ele[0][10] != ele[2][11];
    ele[0][10] != ele[2][12];
    ele[0][10] != ele[2][13];
    ele[0][10] != ele[2][14];
    ele[0][10] != ele[20][10];
    ele[0][10] != ele[21][10];
    ele[0][10] != ele[22][10];
    ele[0][10] != ele[23][10];
    ele[0][10] != ele[24][10];
    ele[0][10] != ele[3][10];
    ele[0][10] != ele[3][11];
    ele[0][10] != ele[3][12];
    ele[0][10] != ele[3][13];
    ele[0][10] != ele[3][14];
    ele[0][10] != ele[4][10];
    ele[0][10] != ele[4][11];
    ele[0][10] != ele[4][12];
    ele[0][10] != ele[4][13];
    ele[0][10] != ele[4][14];
    ele[0][10] != ele[5][10];
    ele[0][10] != ele[6][10];
    ele[0][10] != ele[7][10];
    ele[0][10] != ele[8][10];
    ele[0][10] != ele[9][10];
    ele[0][11] != ele[0][12];
    ele[0][11] != ele[0][13];
    ele[0][11] != ele[0][14];
    ele[0][11] != ele[0][15];
    ele[0][11] != ele[0][16];
    ele[0][11] != ele[0][17];
    ele[0][11] != ele[0][18];
    ele[0][11] != ele[0][19];
    ele[0][11] != ele[0][20];
    ele[0][11] != ele[0][21];
    ele[0][11] != ele[0][22];
    ele[0][11] != ele[0][23];
    ele[0][11] != ele[0][24];
    ele[0][11] != ele[1][10];
    ele[0][11] != ele[1][11];
    ele[0][11] != ele[1][12];
    ele[0][11] != ele[1][13];
    ele[0][11] != ele[1][14];
    ele[0][11] != ele[10][11];
    ele[0][11] != ele[11][11];
    ele[0][11] != ele[12][11];
    ele[0][11] != ele[13][11];
    ele[0][11] != ele[14][11];
    ele[0][11] != ele[15][11];
    ele[0][11] != ele[16][11];
    ele[0][11] != ele[17][11];
    ele[0][11] != ele[18][11];
    ele[0][11] != ele[19][11];
    ele[0][11] != ele[2][10];
    ele[0][11] != ele[2][11];
    ele[0][11] != ele[2][12];
    ele[0][11] != ele[2][13];
    ele[0][11] != ele[2][14];
    ele[0][11] != ele[20][11];
    ele[0][11] != ele[21][11];
    ele[0][11] != ele[22][11];
    ele[0][11] != ele[23][11];
    ele[0][11] != ele[24][11];
    ele[0][11] != ele[3][10];
    ele[0][11] != ele[3][11];
    ele[0][11] != ele[3][12];
    ele[0][11] != ele[3][13];
    ele[0][11] != ele[3][14];
    ele[0][11] != ele[4][10];
    ele[0][11] != ele[4][11];
    ele[0][11] != ele[4][12];
    ele[0][11] != ele[4][13];
    ele[0][11] != ele[4][14];
    ele[0][11] != ele[5][11];
    ele[0][11] != ele[6][11];
    ele[0][11] != ele[7][11];
    ele[0][11] != ele[8][11];
    ele[0][11] != ele[9][11];
    ele[0][12] != ele[0][13];
    ele[0][12] != ele[0][14];
    ele[0][12] != ele[0][15];
    ele[0][12] != ele[0][16];
    ele[0][12] != ele[0][17];
    ele[0][12] != ele[0][18];
    ele[0][12] != ele[0][19];
    ele[0][12] != ele[0][20];
    ele[0][12] != ele[0][21];
    ele[0][12] != ele[0][22];
    ele[0][12] != ele[0][23];
    ele[0][12] != ele[0][24];
    ele[0][12] != ele[1][10];
    ele[0][12] != ele[1][11];
    ele[0][12] != ele[1][12];
    ele[0][12] != ele[1][13];
    ele[0][12] != ele[1][14];
    ele[0][12] != ele[10][12];
    ele[0][12] != ele[11][12];
    ele[0][12] != ele[12][12];
    ele[0][12] != ele[13][12];
    ele[0][12] != ele[14][12];
    ele[0][12] != ele[15][12];
    ele[0][12] != ele[16][12];
    ele[0][12] != ele[17][12];
    ele[0][12] != ele[18][12];
    ele[0][12] != ele[19][12];
    ele[0][12] != ele[2][10];
    ele[0][12] != ele[2][11];
    ele[0][12] != ele[2][12];
    ele[0][12] != ele[2][13];
    ele[0][12] != ele[2][14];
    ele[0][12] != ele[20][12];
    ele[0][12] != ele[21][12];
    ele[0][12] != ele[22][12];
    ele[0][12] != ele[23][12];
    ele[0][12] != ele[24][12];
    ele[0][12] != ele[3][10];
    ele[0][12] != ele[3][11];
    ele[0][12] != ele[3][12];
    ele[0][12] != ele[3][13];
    ele[0][12] != ele[3][14];
    ele[0][12] != ele[4][10];
    ele[0][12] != ele[4][11];
    ele[0][12] != ele[4][12];
    ele[0][12] != ele[4][13];
    ele[0][12] != ele[4][14];
    ele[0][12] != ele[5][12];
    ele[0][12] != ele[6][12];
    ele[0][12] != ele[7][12];
    ele[0][12] != ele[8][12];
    ele[0][12] != ele[9][12];
    ele[0][13] != ele[0][14];
    ele[0][13] != ele[0][15];
    ele[0][13] != ele[0][16];
    ele[0][13] != ele[0][17];
    ele[0][13] != ele[0][18];
    ele[0][13] != ele[0][19];
    ele[0][13] != ele[0][20];
    ele[0][13] != ele[0][21];
    ele[0][13] != ele[0][22];
    ele[0][13] != ele[0][23];
    ele[0][13] != ele[0][24];
    ele[0][13] != ele[1][10];
    ele[0][13] != ele[1][11];
    ele[0][13] != ele[1][12];
    ele[0][13] != ele[1][13];
    ele[0][13] != ele[1][14];
    ele[0][13] != ele[10][13];
    ele[0][13] != ele[11][13];
    ele[0][13] != ele[12][13];
    ele[0][13] != ele[13][13];
    ele[0][13] != ele[14][13];
    ele[0][13] != ele[15][13];
    ele[0][13] != ele[16][13];
    ele[0][13] != ele[17][13];
    ele[0][13] != ele[18][13];
    ele[0][13] != ele[19][13];
    ele[0][13] != ele[2][10];
    ele[0][13] != ele[2][11];
    ele[0][13] != ele[2][12];
    ele[0][13] != ele[2][13];
    ele[0][13] != ele[2][14];
    ele[0][13] != ele[20][13];
    ele[0][13] != ele[21][13];
    ele[0][13] != ele[22][13];
    ele[0][13] != ele[23][13];
    ele[0][13] != ele[24][13];
    ele[0][13] != ele[3][10];
    ele[0][13] != ele[3][11];
    ele[0][13] != ele[3][12];
    ele[0][13] != ele[3][13];
    ele[0][13] != ele[3][14];
    ele[0][13] != ele[4][10];
    ele[0][13] != ele[4][11];
    ele[0][13] != ele[4][12];
    ele[0][13] != ele[4][13];
    ele[0][13] != ele[4][14];
    ele[0][13] != ele[5][13];
    ele[0][13] != ele[6][13];
    ele[0][13] != ele[7][13];
    ele[0][13] != ele[8][13];
    ele[0][13] != ele[9][13];
    ele[0][14] != ele[0][15];
    ele[0][14] != ele[0][16];
    ele[0][14] != ele[0][17];
    ele[0][14] != ele[0][18];
    ele[0][14] != ele[0][19];
    ele[0][14] != ele[0][20];
    ele[0][14] != ele[0][21];
    ele[0][14] != ele[0][22];
    ele[0][14] != ele[0][23];
    ele[0][14] != ele[0][24];
    ele[0][14] != ele[1][10];
    ele[0][14] != ele[1][11];
    ele[0][14] != ele[1][12];
    ele[0][14] != ele[1][13];
    ele[0][14] != ele[1][14];
    ele[0][14] != ele[10][14];
    ele[0][14] != ele[11][14];
    ele[0][14] != ele[12][14];
    ele[0][14] != ele[13][14];
    ele[0][14] != ele[14][14];
    ele[0][14] != ele[15][14];
    ele[0][14] != ele[16][14];
    ele[0][14] != ele[17][14];
    ele[0][14] != ele[18][14];
    ele[0][14] != ele[19][14];
    ele[0][14] != ele[2][10];
    ele[0][14] != ele[2][11];
    ele[0][14] != ele[2][12];
    ele[0][14] != ele[2][13];
    ele[0][14] != ele[2][14];
    ele[0][14] != ele[20][14];
    ele[0][14] != ele[21][14];
    ele[0][14] != ele[22][14];
    ele[0][14] != ele[23][14];
    ele[0][14] != ele[24][14];
    ele[0][14] != ele[3][10];
    ele[0][14] != ele[3][11];
    ele[0][14] != ele[3][12];
    ele[0][14] != ele[3][13];
    ele[0][14] != ele[3][14];
    ele[0][14] != ele[4][10];
    ele[0][14] != ele[4][11];
    ele[0][14] != ele[4][12];
    ele[0][14] != ele[4][13];
    ele[0][14] != ele[4][14];
    ele[0][14] != ele[5][14];
    ele[0][14] != ele[6][14];
    ele[0][14] != ele[7][14];
    ele[0][14] != ele[8][14];
    ele[0][14] != ele[9][14];
    ele[0][15] != ele[0][16];
    ele[0][15] != ele[0][17];
    ele[0][15] != ele[0][18];
    ele[0][15] != ele[0][19];
    ele[0][15] != ele[0][20];
    ele[0][15] != ele[0][21];
    ele[0][15] != ele[0][22];
    ele[0][15] != ele[0][23];
    ele[0][15] != ele[0][24];
    ele[0][15] != ele[1][15];
    ele[0][15] != ele[1][16];
    ele[0][15] != ele[1][17];
    ele[0][15] != ele[1][18];
    ele[0][15] != ele[1][19];
    ele[0][15] != ele[10][15];
    ele[0][15] != ele[11][15];
    ele[0][15] != ele[12][15];
    ele[0][15] != ele[13][15];
    ele[0][15] != ele[14][15];
    ele[0][15] != ele[15][15];
    ele[0][15] != ele[16][15];
    ele[0][15] != ele[17][15];
    ele[0][15] != ele[18][15];
    ele[0][15] != ele[19][15];
    ele[0][15] != ele[2][15];
    ele[0][15] != ele[2][16];
    ele[0][15] != ele[2][17];
    ele[0][15] != ele[2][18];
    ele[0][15] != ele[2][19];
    ele[0][15] != ele[20][15];
    ele[0][15] != ele[21][15];
    ele[0][15] != ele[22][15];
    ele[0][15] != ele[23][15];
    ele[0][15] != ele[24][15];
    ele[0][15] != ele[3][15];
    ele[0][15] != ele[3][16];
    ele[0][15] != ele[3][17];
    ele[0][15] != ele[3][18];
    ele[0][15] != ele[3][19];
    ele[0][15] != ele[4][15];
    ele[0][15] != ele[4][16];
    ele[0][15] != ele[4][17];
    ele[0][15] != ele[4][18];
    ele[0][15] != ele[4][19];
    ele[0][15] != ele[5][15];
    ele[0][15] != ele[6][15];
    ele[0][15] != ele[7][15];
    ele[0][15] != ele[8][15];
    ele[0][15] != ele[9][15];
    ele[0][16] != ele[0][17];
    ele[0][16] != ele[0][18];
    ele[0][16] != ele[0][19];
    ele[0][16] != ele[0][20];
    ele[0][16] != ele[0][21];
    ele[0][16] != ele[0][22];
    ele[0][16] != ele[0][23];
    ele[0][16] != ele[0][24];
    ele[0][16] != ele[1][15];
    ele[0][16] != ele[1][16];
    ele[0][16] != ele[1][17];
    ele[0][16] != ele[1][18];
    ele[0][16] != ele[1][19];
    ele[0][16] != ele[10][16];
    ele[0][16] != ele[11][16];
    ele[0][16] != ele[12][16];
    ele[0][16] != ele[13][16];
    ele[0][16] != ele[14][16];
    ele[0][16] != ele[15][16];
    ele[0][16] != ele[16][16];
    ele[0][16] != ele[17][16];
    ele[0][16] != ele[18][16];
    ele[0][16] != ele[19][16];
    ele[0][16] != ele[2][15];
    ele[0][16] != ele[2][16];
    ele[0][16] != ele[2][17];
    ele[0][16] != ele[2][18];
    ele[0][16] != ele[2][19];
    ele[0][16] != ele[20][16];
    ele[0][16] != ele[21][16];
    ele[0][16] != ele[22][16];
    ele[0][16] != ele[23][16];
    ele[0][16] != ele[24][16];
    ele[0][16] != ele[3][15];
    ele[0][16] != ele[3][16];
    ele[0][16] != ele[3][17];
    ele[0][16] != ele[3][18];
    ele[0][16] != ele[3][19];
    ele[0][16] != ele[4][15];
    ele[0][16] != ele[4][16];
    ele[0][16] != ele[4][17];
    ele[0][16] != ele[4][18];
    ele[0][16] != ele[4][19];
    ele[0][16] != ele[5][16];
    ele[0][16] != ele[6][16];
    ele[0][16] != ele[7][16];
    ele[0][16] != ele[8][16];
    ele[0][16] != ele[9][16];
    ele[0][17] != ele[0][18];
    ele[0][17] != ele[0][19];
    ele[0][17] != ele[0][20];
    ele[0][17] != ele[0][21];
    ele[0][17] != ele[0][22];
    ele[0][17] != ele[0][23];
    ele[0][17] != ele[0][24];
    ele[0][17] != ele[1][15];
    ele[0][17] != ele[1][16];
    ele[0][17] != ele[1][17];
    ele[0][17] != ele[1][18];
    ele[0][17] != ele[1][19];
    ele[0][17] != ele[10][17];
    ele[0][17] != ele[11][17];
    ele[0][17] != ele[12][17];
    ele[0][17] != ele[13][17];
    ele[0][17] != ele[14][17];
    ele[0][17] != ele[15][17];
    ele[0][17] != ele[16][17];
    ele[0][17] != ele[17][17];
    ele[0][17] != ele[18][17];
    ele[0][17] != ele[19][17];
    ele[0][17] != ele[2][15];
    ele[0][17] != ele[2][16];
    ele[0][17] != ele[2][17];
    ele[0][17] != ele[2][18];
    ele[0][17] != ele[2][19];
    ele[0][17] != ele[20][17];
    ele[0][17] != ele[21][17];
    ele[0][17] != ele[22][17];
    ele[0][17] != ele[23][17];
    ele[0][17] != ele[24][17];
    ele[0][17] != ele[3][15];
    ele[0][17] != ele[3][16];
    ele[0][17] != ele[3][17];
    ele[0][17] != ele[3][18];
    ele[0][17] != ele[3][19];
    ele[0][17] != ele[4][15];
    ele[0][17] != ele[4][16];
    ele[0][17] != ele[4][17];
    ele[0][17] != ele[4][18];
    ele[0][17] != ele[4][19];
    ele[0][17] != ele[5][17];
    ele[0][17] != ele[6][17];
    ele[0][17] != ele[7][17];
    ele[0][17] != ele[8][17];
    ele[0][17] != ele[9][17];
    ele[0][18] != ele[0][19];
    ele[0][18] != ele[0][20];
    ele[0][18] != ele[0][21];
    ele[0][18] != ele[0][22];
    ele[0][18] != ele[0][23];
    ele[0][18] != ele[0][24];
    ele[0][18] != ele[1][15];
    ele[0][18] != ele[1][16];
    ele[0][18] != ele[1][17];
    ele[0][18] != ele[1][18];
    ele[0][18] != ele[1][19];
    ele[0][18] != ele[10][18];
    ele[0][18] != ele[11][18];
    ele[0][18] != ele[12][18];
    ele[0][18] != ele[13][18];
    ele[0][18] != ele[14][18];
    ele[0][18] != ele[15][18];
    ele[0][18] != ele[16][18];
    ele[0][18] != ele[17][18];
    ele[0][18] != ele[18][18];
    ele[0][18] != ele[19][18];
    ele[0][18] != ele[2][15];
    ele[0][18] != ele[2][16];
    ele[0][18] != ele[2][17];
    ele[0][18] != ele[2][18];
    ele[0][18] != ele[2][19];
    ele[0][18] != ele[20][18];
    ele[0][18] != ele[21][18];
    ele[0][18] != ele[22][18];
    ele[0][18] != ele[23][18];
    ele[0][18] != ele[24][18];
    ele[0][18] != ele[3][15];
    ele[0][18] != ele[3][16];
    ele[0][18] != ele[3][17];
    ele[0][18] != ele[3][18];
    ele[0][18] != ele[3][19];
    ele[0][18] != ele[4][15];
    ele[0][18] != ele[4][16];
    ele[0][18] != ele[4][17];
    ele[0][18] != ele[4][18];
    ele[0][18] != ele[4][19];
    ele[0][18] != ele[5][18];
    ele[0][18] != ele[6][18];
    ele[0][18] != ele[7][18];
    ele[0][18] != ele[8][18];
    ele[0][18] != ele[9][18];
    ele[0][19] != ele[0][20];
    ele[0][19] != ele[0][21];
    ele[0][19] != ele[0][22];
    ele[0][19] != ele[0][23];
    ele[0][19] != ele[0][24];
    ele[0][19] != ele[1][15];
    ele[0][19] != ele[1][16];
    ele[0][19] != ele[1][17];
    ele[0][19] != ele[1][18];
    ele[0][19] != ele[1][19];
    ele[0][19] != ele[10][19];
    ele[0][19] != ele[11][19];
    ele[0][19] != ele[12][19];
    ele[0][19] != ele[13][19];
    ele[0][19] != ele[14][19];
    ele[0][19] != ele[15][19];
    ele[0][19] != ele[16][19];
    ele[0][19] != ele[17][19];
    ele[0][19] != ele[18][19];
    ele[0][19] != ele[19][19];
    ele[0][19] != ele[2][15];
    ele[0][19] != ele[2][16];
    ele[0][19] != ele[2][17];
    ele[0][19] != ele[2][18];
    ele[0][19] != ele[2][19];
    ele[0][19] != ele[20][19];
    ele[0][19] != ele[21][19];
    ele[0][19] != ele[22][19];
    ele[0][19] != ele[23][19];
    ele[0][19] != ele[24][19];
    ele[0][19] != ele[3][15];
    ele[0][19] != ele[3][16];
    ele[0][19] != ele[3][17];
    ele[0][19] != ele[3][18];
    ele[0][19] != ele[3][19];
    ele[0][19] != ele[4][15];
    ele[0][19] != ele[4][16];
    ele[0][19] != ele[4][17];
    ele[0][19] != ele[4][18];
    ele[0][19] != ele[4][19];
    ele[0][19] != ele[5][19];
    ele[0][19] != ele[6][19];
    ele[0][19] != ele[7][19];
    ele[0][19] != ele[8][19];
    ele[0][19] != ele[9][19];
    ele[0][2] != ele[0][10];
    ele[0][2] != ele[0][11];
    ele[0][2] != ele[0][12];
    ele[0][2] != ele[0][13];
    ele[0][2] != ele[0][14];
    ele[0][2] != ele[0][15];
    ele[0][2] != ele[0][16];
    ele[0][2] != ele[0][17];
    ele[0][2] != ele[0][18];
    ele[0][2] != ele[0][19];
    ele[0][2] != ele[0][20];
    ele[0][2] != ele[0][21];
    ele[0][2] != ele[0][22];
    ele[0][2] != ele[0][23];
    ele[0][2] != ele[0][24];
    ele[0][2] != ele[0][3];
    ele[0][2] != ele[0][4];
    ele[0][2] != ele[0][5];
    ele[0][2] != ele[0][6];
    ele[0][2] != ele[0][7];
    ele[0][2] != ele[0][8];
    ele[0][2] != ele[0][9];
    ele[0][2] != ele[1][0];
    ele[0][2] != ele[1][1];
    ele[0][2] != ele[1][2];
    ele[0][2] != ele[1][3];
    ele[0][2] != ele[1][4];
    ele[0][2] != ele[10][2];
    ele[0][2] != ele[11][2];
    ele[0][2] != ele[12][2];
    ele[0][2] != ele[13][2];
    ele[0][2] != ele[14][2];
    ele[0][2] != ele[15][2];
    ele[0][2] != ele[16][2];
    ele[0][2] != ele[17][2];
    ele[0][2] != ele[18][2];
    ele[0][2] != ele[19][2];
    ele[0][2] != ele[2][0];
    ele[0][2] != ele[2][1];
    ele[0][2] != ele[2][2];
    ele[0][2] != ele[2][3];
    ele[0][2] != ele[2][4];
    ele[0][2] != ele[20][2];
    ele[0][2] != ele[21][2];
    ele[0][2] != ele[22][2];
    ele[0][2] != ele[23][2];
    ele[0][2] != ele[24][2];
    ele[0][2] != ele[3][0];
    ele[0][2] != ele[3][1];
    ele[0][2] != ele[3][2];
    ele[0][2] != ele[3][3];
    ele[0][2] != ele[3][4];
    ele[0][2] != ele[4][0];
    ele[0][2] != ele[4][1];
    ele[0][2] != ele[4][2];
    ele[0][2] != ele[4][3];
    ele[0][2] != ele[4][4];
    ele[0][2] != ele[5][2];
    ele[0][2] != ele[6][2];
    ele[0][2] != ele[7][2];
    ele[0][2] != ele[8][2];
    ele[0][2] != ele[9][2];
    ele[0][20] != ele[0][21];
    ele[0][20] != ele[0][22];
    ele[0][20] != ele[0][23];
    ele[0][20] != ele[0][24];
    ele[0][20] != ele[1][20];
    ele[0][20] != ele[1][21];
    ele[0][20] != ele[1][22];
    ele[0][20] != ele[1][23];
    ele[0][20] != ele[1][24];
    ele[0][20] != ele[10][20];
    ele[0][20] != ele[11][20];
    ele[0][20] != ele[12][20];
    ele[0][20] != ele[13][20];
    ele[0][20] != ele[14][20];
    ele[0][20] != ele[15][20];
    ele[0][20] != ele[16][20];
    ele[0][20] != ele[17][20];
    ele[0][20] != ele[18][20];
    ele[0][20] != ele[19][20];
    ele[0][20] != ele[2][20];
    ele[0][20] != ele[2][21];
    ele[0][20] != ele[2][22];
    ele[0][20] != ele[2][23];
    ele[0][20] != ele[2][24];
    ele[0][20] != ele[20][20];
    ele[0][20] != ele[21][20];
    ele[0][20] != ele[22][20];
    ele[0][20] != ele[23][20];
    ele[0][20] != ele[24][20];
    ele[0][20] != ele[3][20];
    ele[0][20] != ele[3][21];
    ele[0][20] != ele[3][22];
    ele[0][20] != ele[3][23];
    ele[0][20] != ele[3][24];
    ele[0][20] != ele[4][20];
    ele[0][20] != ele[4][21];
    ele[0][20] != ele[4][22];
    ele[0][20] != ele[4][23];
    ele[0][20] != ele[4][24];
    ele[0][20] != ele[5][20];
    ele[0][20] != ele[6][20];
    ele[0][20] != ele[7][20];
    ele[0][20] != ele[8][20];
    ele[0][20] != ele[9][20];
    ele[0][21] != ele[0][22];
    ele[0][21] != ele[0][23];
    ele[0][21] != ele[0][24];
    ele[0][21] != ele[1][20];
    ele[0][21] != ele[1][21];
    ele[0][21] != ele[1][22];
    ele[0][21] != ele[1][23];
    ele[0][21] != ele[1][24];
    ele[0][21] != ele[10][21];
    ele[0][21] != ele[11][21];
    ele[0][21] != ele[12][21];
    ele[0][21] != ele[13][21];
    ele[0][21] != ele[14][21];
    ele[0][21] != ele[15][21];
    ele[0][21] != ele[16][21];
    ele[0][21] != ele[17][21];
    ele[0][21] != ele[18][21];
    ele[0][21] != ele[19][21];
    ele[0][21] != ele[2][20];
    ele[0][21] != ele[2][21];
    ele[0][21] != ele[2][22];
    ele[0][21] != ele[2][23];
    ele[0][21] != ele[2][24];
    ele[0][21] != ele[20][21];
    ele[0][21] != ele[21][21];
    ele[0][21] != ele[22][21];
    ele[0][21] != ele[23][21];
    ele[0][21] != ele[24][21];
    ele[0][21] != ele[3][20];
    ele[0][21] != ele[3][21];
    ele[0][21] != ele[3][22];
    ele[0][21] != ele[3][23];
    ele[0][21] != ele[3][24];
    ele[0][21] != ele[4][20];
    ele[0][21] != ele[4][21];
    ele[0][21] != ele[4][22];
    ele[0][21] != ele[4][23];
    ele[0][21] != ele[4][24];
    ele[0][21] != ele[5][21];
    ele[0][21] != ele[6][21];
    ele[0][21] != ele[7][21];
    ele[0][21] != ele[8][21];
    ele[0][21] != ele[9][21];
    ele[0][22] != ele[0][23];
    ele[0][22] != ele[0][24];
    ele[0][22] != ele[1][20];
    ele[0][22] != ele[1][21];
    ele[0][22] != ele[1][22];
    ele[0][22] != ele[1][23];
    ele[0][22] != ele[1][24];
    ele[0][22] != ele[10][22];
    ele[0][22] != ele[11][22];
    ele[0][22] != ele[12][22];
    ele[0][22] != ele[13][22];
    ele[0][22] != ele[14][22];
    ele[0][22] != ele[15][22];
    ele[0][22] != ele[16][22];
    ele[0][22] != ele[17][22];
    ele[0][22] != ele[18][22];
    ele[0][22] != ele[19][22];
    ele[0][22] != ele[2][20];
    ele[0][22] != ele[2][21];
    ele[0][22] != ele[2][22];
    ele[0][22] != ele[2][23];
    ele[0][22] != ele[2][24];
    ele[0][22] != ele[20][22];
    ele[0][22] != ele[21][22];
    ele[0][22] != ele[22][22];
    ele[0][22] != ele[23][22];
    ele[0][22] != ele[24][22];
    ele[0][22] != ele[3][20];
    ele[0][22] != ele[3][21];
    ele[0][22] != ele[3][22];
    ele[0][22] != ele[3][23];
    ele[0][22] != ele[3][24];
    ele[0][22] != ele[4][20];
    ele[0][22] != ele[4][21];
    ele[0][22] != ele[4][22];
    ele[0][22] != ele[4][23];
    ele[0][22] != ele[4][24];
    ele[0][22] != ele[5][22];
    ele[0][22] != ele[6][22];
    ele[0][22] != ele[7][22];
    ele[0][22] != ele[8][22];
    ele[0][22] != ele[9][22];
    ele[0][23] != ele[0][24];
    ele[0][23] != ele[1][20];
    ele[0][23] != ele[1][21];
    ele[0][23] != ele[1][22];
    ele[0][23] != ele[1][23];
    ele[0][23] != ele[1][24];
    ele[0][23] != ele[10][23];
    ele[0][23] != ele[11][23];
    ele[0][23] != ele[12][23];
    ele[0][23] != ele[13][23];
    ele[0][23] != ele[14][23];
    ele[0][23] != ele[15][23];
    ele[0][23] != ele[16][23];
    ele[0][23] != ele[17][23];
    ele[0][23] != ele[18][23];
    ele[0][23] != ele[19][23];
    ele[0][23] != ele[2][20];
    ele[0][23] != ele[2][21];
    ele[0][23] != ele[2][22];
    ele[0][23] != ele[2][23];
    ele[0][23] != ele[2][24];
    ele[0][23] != ele[20][23];
    ele[0][23] != ele[21][23];
    ele[0][23] != ele[22][23];
    ele[0][23] != ele[23][23];
    ele[0][23] != ele[24][23];
    ele[0][23] != ele[3][20];
    ele[0][23] != ele[3][21];
    ele[0][23] != ele[3][22];
    ele[0][23] != ele[3][23];
    ele[0][23] != ele[3][24];
    ele[0][23] != ele[4][20];
    ele[0][23] != ele[4][21];
    ele[0][23] != ele[4][22];
    ele[0][23] != ele[4][23];
    ele[0][23] != ele[4][24];
    ele[0][23] != ele[5][23];
    ele[0][23] != ele[6][23];
    ele[0][23] != ele[7][23];
    ele[0][23] != ele[8][23];
    ele[0][23] != ele[9][23];
    ele[0][24] != ele[1][20];
    ele[0][24] != ele[1][21];
    ele[0][24] != ele[1][22];
    ele[0][24] != ele[1][23];
    ele[0][24] != ele[1][24];
    ele[0][24] != ele[10][24];
    ele[0][24] != ele[11][24];
    ele[0][24] != ele[12][24];
    ele[0][24] != ele[13][24];
    ele[0][24] != ele[14][24];
    ele[0][24] != ele[15][24];
    ele[0][24] != ele[16][24];
    ele[0][24] != ele[17][24];
    ele[0][24] != ele[18][24];
    ele[0][24] != ele[19][24];
    ele[0][24] != ele[2][20];
    ele[0][24] != ele[2][21];
    ele[0][24] != ele[2][22];
    ele[0][24] != ele[2][23];
    ele[0][24] != ele[2][24];
    ele[0][24] != ele[20][24];
    ele[0][24] != ele[21][24];
    ele[0][24] != ele[22][24];
    ele[0][24] != ele[23][24];
    ele[0][24] != ele[24][24];
    ele[0][24] != ele[3][20];
    ele[0][24] != ele[3][21];
    ele[0][24] != ele[3][22];
    ele[0][24] != ele[3][23];
    ele[0][24] != ele[3][24];
    ele[0][24] != ele[4][20];
    ele[0][24] != ele[4][21];
    ele[0][24] != ele[4][22];
    ele[0][24] != ele[4][23];
    ele[0][24] != ele[4][24];
    ele[0][24] != ele[5][24];
    ele[0][24] != ele[6][24];
    ele[0][24] != ele[7][24];
    ele[0][24] != ele[8][24];
    ele[0][24] != ele[9][24];
    ele[0][3] != ele[0][10];
    ele[0][3] != ele[0][11];
    ele[0][3] != ele[0][12];
    ele[0][3] != ele[0][13];
    ele[0][3] != ele[0][14];
    ele[0][3] != ele[0][15];
    ele[0][3] != ele[0][16];
    ele[0][3] != ele[0][17];
    ele[0][3] != ele[0][18];
    ele[0][3] != ele[0][19];
    ele[0][3] != ele[0][20];
    ele[0][3] != ele[0][21];
    ele[0][3] != ele[0][22];
    ele[0][3] != ele[0][23];
    ele[0][3] != ele[0][24];
    ele[0][3] != ele[0][4];
    ele[0][3] != ele[0][5];
    ele[0][3] != ele[0][6];
    ele[0][3] != ele[0][7];
    ele[0][3] != ele[0][8];
    ele[0][3] != ele[0][9];
    ele[0][3] != ele[1][0];
    ele[0][3] != ele[1][1];
    ele[0][3] != ele[1][2];
    ele[0][3] != ele[1][3];
    ele[0][3] != ele[1][4];
    ele[0][3] != ele[10][3];
    ele[0][3] != ele[11][3];
    ele[0][3] != ele[12][3];
    ele[0][3] != ele[13][3];
    ele[0][3] != ele[14][3];
    ele[0][3] != ele[15][3];
    ele[0][3] != ele[16][3];
    ele[0][3] != ele[17][3];
    ele[0][3] != ele[18][3];
    ele[0][3] != ele[19][3];
    ele[0][3] != ele[2][0];
    ele[0][3] != ele[2][1];
    ele[0][3] != ele[2][2];
    ele[0][3] != ele[2][3];
    ele[0][3] != ele[2][4];
    ele[0][3] != ele[20][3];
    ele[0][3] != ele[21][3];
    ele[0][3] != ele[22][3];
    ele[0][3] != ele[23][3];
    ele[0][3] != ele[24][3];
    ele[0][3] != ele[3][0];
    ele[0][3] != ele[3][1];
    ele[0][3] != ele[3][2];
    ele[0][3] != ele[3][3];
    ele[0][3] != ele[3][4];
    ele[0][3] != ele[4][0];
    ele[0][3] != ele[4][1];
    ele[0][3] != ele[4][2];
    ele[0][3] != ele[4][3];
    ele[0][3] != ele[4][4];
    ele[0][3] != ele[5][3];
    ele[0][3] != ele[6][3];
    ele[0][3] != ele[7][3];
    ele[0][3] != ele[8][3];
    ele[0][3] != ele[9][3];
    ele[0][4] != ele[0][10];
    ele[0][4] != ele[0][11];
    ele[0][4] != ele[0][12];
    ele[0][4] != ele[0][13];
    ele[0][4] != ele[0][14];
    ele[0][4] != ele[0][15];
    ele[0][4] != ele[0][16];
    ele[0][4] != ele[0][17];
    ele[0][4] != ele[0][18];
    ele[0][4] != ele[0][19];
    ele[0][4] != ele[0][20];
    ele[0][4] != ele[0][21];
    ele[0][4] != ele[0][22];
    ele[0][4] != ele[0][23];
    ele[0][4] != ele[0][24];
    ele[0][4] != ele[0][5];
    ele[0][4] != ele[0][6];
    ele[0][4] != ele[0][7];
    ele[0][4] != ele[0][8];
    ele[0][4] != ele[0][9];
    ele[0][4] != ele[1][0];
    ele[0][4] != ele[1][1];
    ele[0][4] != ele[1][2];
    ele[0][4] != ele[1][3];
    ele[0][4] != ele[1][4];
    ele[0][4] != ele[10][4];
    ele[0][4] != ele[11][4];
    ele[0][4] != ele[12][4];
    ele[0][4] != ele[13][4];
    ele[0][4] != ele[14][4];
    ele[0][4] != ele[15][4];
    ele[0][4] != ele[16][4];
    ele[0][4] != ele[17][4];
    ele[0][4] != ele[18][4];
    ele[0][4] != ele[19][4];
    ele[0][4] != ele[2][0];
    ele[0][4] != ele[2][1];
    ele[0][4] != ele[2][2];
    ele[0][4] != ele[2][3];
    ele[0][4] != ele[2][4];
    ele[0][4] != ele[20][4];
    ele[0][4] != ele[21][4];
    ele[0][4] != ele[22][4];
    ele[0][4] != ele[23][4];
    ele[0][4] != ele[24][4];
    ele[0][4] != ele[3][0];
    ele[0][4] != ele[3][1];
    ele[0][4] != ele[3][2];
    ele[0][4] != ele[3][3];
    ele[0][4] != ele[3][4];
    ele[0][4] != ele[4][0];
    ele[0][4] != ele[4][1];
    ele[0][4] != ele[4][2];
    ele[0][4] != ele[4][3];
    ele[0][4] != ele[4][4];
    ele[0][4] != ele[5][4];
    ele[0][4] != ele[6][4];
    ele[0][4] != ele[7][4];
    ele[0][4] != ele[8][4];
    ele[0][4] != ele[9][4];
    ele[0][5] != ele[0][10];
    ele[0][5] != ele[0][11];
    ele[0][5] != ele[0][12];
    ele[0][5] != ele[0][13];
    ele[0][5] != ele[0][14];
    ele[0][5] != ele[0][15];
    ele[0][5] != ele[0][16];
    ele[0][5] != ele[0][17];
    ele[0][5] != ele[0][18];
    ele[0][5] != ele[0][19];
    ele[0][5] != ele[0][20];
    ele[0][5] != ele[0][21];
    ele[0][5] != ele[0][22];
    ele[0][5] != ele[0][23];
    ele[0][5] != ele[0][24];
    ele[0][5] != ele[0][6];
    ele[0][5] != ele[0][7];
    ele[0][5] != ele[0][8];
    ele[0][5] != ele[0][9];
    ele[0][5] != ele[1][5];
    ele[0][5] != ele[1][6];
    ele[0][5] != ele[1][7];
    ele[0][5] != ele[1][8];
    ele[0][5] != ele[1][9];
    ele[0][5] != ele[10][5];
    ele[0][5] != ele[11][5];
    ele[0][5] != ele[12][5];
    ele[0][5] != ele[13][5];
    ele[0][5] != ele[14][5];
    ele[0][5] != ele[15][5];
    ele[0][5] != ele[16][5];
    ele[0][5] != ele[17][5];
    ele[0][5] != ele[18][5];
    ele[0][5] != ele[19][5];
    ele[0][5] != ele[2][5];
    ele[0][5] != ele[2][6];
    ele[0][5] != ele[2][7];
    ele[0][5] != ele[2][8];
    ele[0][5] != ele[2][9];
    ele[0][5] != ele[20][5];
    ele[0][5] != ele[21][5];
    ele[0][5] != ele[22][5];
    ele[0][5] != ele[23][5];
    ele[0][5] != ele[24][5];
    ele[0][5] != ele[3][5];
    ele[0][5] != ele[3][6];
    ele[0][5] != ele[3][7];
    ele[0][5] != ele[3][8];
    ele[0][5] != ele[3][9];
    ele[0][5] != ele[4][5];
    ele[0][5] != ele[4][6];
    ele[0][5] != ele[4][7];
    ele[0][5] != ele[4][8];
    ele[0][5] != ele[4][9];
    ele[0][5] != ele[5][5];
    ele[0][5] != ele[6][5];
    ele[0][5] != ele[7][5];
    ele[0][5] != ele[8][5];
    ele[0][5] != ele[9][5];
    ele[0][6] != ele[0][10];
    ele[0][6] != ele[0][11];
    ele[0][6] != ele[0][12];
    ele[0][6] != ele[0][13];
    ele[0][6] != ele[0][14];
    ele[0][6] != ele[0][15];
    ele[0][6] != ele[0][16];
    ele[0][6] != ele[0][17];
    ele[0][6] != ele[0][18];
    ele[0][6] != ele[0][19];
    ele[0][6] != ele[0][20];
    ele[0][6] != ele[0][21];
    ele[0][6] != ele[0][22];
    ele[0][6] != ele[0][23];
    ele[0][6] != ele[0][24];
    ele[0][6] != ele[0][7];
    ele[0][6] != ele[0][8];
    ele[0][6] != ele[0][9];
    ele[0][6] != ele[1][5];
    ele[0][6] != ele[1][6];
    ele[0][6] != ele[1][7];
    ele[0][6] != ele[1][8];
    ele[0][6] != ele[1][9];
    ele[0][6] != ele[10][6];
    ele[0][6] != ele[11][6];
    ele[0][6] != ele[12][6];
    ele[0][6] != ele[13][6];
    ele[0][6] != ele[14][6];
    ele[0][6] != ele[15][6];
    ele[0][6] != ele[16][6];
    ele[0][6] != ele[17][6];
    ele[0][6] != ele[18][6];
    ele[0][6] != ele[19][6];
    ele[0][6] != ele[2][5];
    ele[0][6] != ele[2][6];
    ele[0][6] != ele[2][7];
    ele[0][6] != ele[2][8];
    ele[0][6] != ele[2][9];
    ele[0][6] != ele[20][6];
    ele[0][6] != ele[21][6];
    ele[0][6] != ele[22][6];
    ele[0][6] != ele[23][6];
    ele[0][6] != ele[24][6];
    ele[0][6] != ele[3][5];
    ele[0][6] != ele[3][6];
    ele[0][6] != ele[3][7];
    ele[0][6] != ele[3][8];
    ele[0][6] != ele[3][9];
    ele[0][6] != ele[4][5];
    ele[0][6] != ele[4][6];
    ele[0][6] != ele[4][7];
    ele[0][6] != ele[4][8];
    ele[0][6] != ele[4][9];
    ele[0][6] != ele[5][6];
    ele[0][6] != ele[6][6];
    ele[0][6] != ele[7][6];
    ele[0][6] != ele[8][6];
    ele[0][6] != ele[9][6];
    ele[0][7] != ele[0][10];
    ele[0][7] != ele[0][11];
    ele[0][7] != ele[0][12];
    ele[0][7] != ele[0][13];
    ele[0][7] != ele[0][14];
    ele[0][7] != ele[0][15];
    ele[0][7] != ele[0][16];
    ele[0][7] != ele[0][17];
    ele[0][7] != ele[0][18];
    ele[0][7] != ele[0][19];
    ele[0][7] != ele[0][20];
    ele[0][7] != ele[0][21];
    ele[0][7] != ele[0][22];
    ele[0][7] != ele[0][23];
    ele[0][7] != ele[0][24];
    ele[0][7] != ele[0][8];
    ele[0][7] != ele[0][9];
    ele[0][7] != ele[1][5];
    ele[0][7] != ele[1][6];
    ele[0][7] != ele[1][7];
    ele[0][7] != ele[1][8];
    ele[0][7] != ele[1][9];
    ele[0][7] != ele[10][7];
    ele[0][7] != ele[11][7];
    ele[0][7] != ele[12][7];
    ele[0][7] != ele[13][7];
    ele[0][7] != ele[14][7];
    ele[0][7] != ele[15][7];
    ele[0][7] != ele[16][7];
    ele[0][7] != ele[17][7];
    ele[0][7] != ele[18][7];
    ele[0][7] != ele[19][7];
    ele[0][7] != ele[2][5];
    ele[0][7] != ele[2][6];
    ele[0][7] != ele[2][7];
    ele[0][7] != ele[2][8];
    ele[0][7] != ele[2][9];
    ele[0][7] != ele[20][7];
    ele[0][7] != ele[21][7];
    ele[0][7] != ele[22][7];
    ele[0][7] != ele[23][7];
    ele[0][7] != ele[24][7];
    ele[0][7] != ele[3][5];
    ele[0][7] != ele[3][6];
    ele[0][7] != ele[3][7];
    ele[0][7] != ele[3][8];
    ele[0][7] != ele[3][9];
    ele[0][7] != ele[4][5];
    ele[0][7] != ele[4][6];
    ele[0][7] != ele[4][7];
    ele[0][7] != ele[4][8];
    ele[0][7] != ele[4][9];
    ele[0][7] != ele[5][7];
    ele[0][7] != ele[6][7];
    ele[0][7] != ele[7][7];
    ele[0][7] != ele[8][7];
    ele[0][7] != ele[9][7];
    ele[0][8] != ele[0][10];
    ele[0][8] != ele[0][11];
    ele[0][8] != ele[0][12];
    ele[0][8] != ele[0][13];
    ele[0][8] != ele[0][14];
    ele[0][8] != ele[0][15];
    ele[0][8] != ele[0][16];
    ele[0][8] != ele[0][17];
    ele[0][8] != ele[0][18];
    ele[0][8] != ele[0][19];
    ele[0][8] != ele[0][20];
    ele[0][8] != ele[0][21];
    ele[0][8] != ele[0][22];
    ele[0][8] != ele[0][23];
    ele[0][8] != ele[0][24];
    ele[0][8] != ele[0][9];
    ele[0][8] != ele[1][5];
    ele[0][8] != ele[1][6];
    ele[0][8] != ele[1][7];
    ele[0][8] != ele[1][8];
    ele[0][8] != ele[1][9];
    ele[0][8] != ele[10][8];
    ele[0][8] != ele[11][8];
    ele[0][8] != ele[12][8];
    ele[0][8] != ele[13][8];
    ele[0][8] != ele[14][8];
    ele[0][8] != ele[15][8];
    ele[0][8] != ele[16][8];
    ele[0][8] != ele[17][8];
    ele[0][8] != ele[18][8];
    ele[0][8] != ele[19][8];
    ele[0][8] != ele[2][5];
    ele[0][8] != ele[2][6];
    ele[0][8] != ele[2][7];
    ele[0][8] != ele[2][8];
    ele[0][8] != ele[2][9];
    ele[0][8] != ele[20][8];
    ele[0][8] != ele[21][8];
    ele[0][8] != ele[22][8];
    ele[0][8] != ele[23][8];
    ele[0][8] != ele[24][8];
    ele[0][8] != ele[3][5];
    ele[0][8] != ele[3][6];
    ele[0][8] != ele[3][7];
    ele[0][8] != ele[3][8];
    ele[0][8] != ele[3][9];
    ele[0][8] != ele[4][5];
    ele[0][8] != ele[4][6];
    ele[0][8] != ele[4][7];
    ele[0][8] != ele[4][8];
    ele[0][8] != ele[4][9];
    ele[0][8] != ele[5][8];
    ele[0][8] != ele[6][8];
    ele[0][8] != ele[7][8];
    ele[0][8] != ele[8][8];
    ele[0][8] != ele[9][8];
    ele[0][9] != ele[0][10];
    ele[0][9] != ele[0][11];
    ele[0][9] != ele[0][12];
    ele[0][9] != ele[0][13];
    ele[0][9] != ele[0][14];
    ele[0][9] != ele[0][15];
    ele[0][9] != ele[0][16];
    ele[0][9] != ele[0][17];
    ele[0][9] != ele[0][18];
    ele[0][9] != ele[0][19];
    ele[0][9] != ele[0][20];
    ele[0][9] != ele[0][21];
    ele[0][9] != ele[0][22];
    ele[0][9] != ele[0][23];
    ele[0][9] != ele[0][24];
    ele[0][9] != ele[1][5];
    ele[0][9] != ele[1][6];
    ele[0][9] != ele[1][7];
    ele[0][9] != ele[1][8];
    ele[0][9] != ele[1][9];
    ele[0][9] != ele[10][9];
    ele[0][9] != ele[11][9];
    ele[0][9] != ele[12][9];
    ele[0][9] != ele[13][9];
    ele[0][9] != ele[14][9];
    ele[0][9] != ele[15][9];
    ele[0][9] != ele[16][9];
    ele[0][9] != ele[17][9];
    ele[0][9] != ele[18][9];
    ele[0][9] != ele[19][9];
    ele[0][9] != ele[2][5];
    ele[0][9] != ele[2][6];
    ele[0][9] != ele[2][7];
    ele[0][9] != ele[2][8];
    ele[0][9] != ele[2][9];
    ele[0][9] != ele[20][9];
    ele[0][9] != ele[21][9];
    ele[0][9] != ele[22][9];
    ele[0][9] != ele[23][9];
    ele[0][9] != ele[24][9];
    ele[0][9] != ele[3][5];
    ele[0][9] != ele[3][6];
    ele[0][9] != ele[3][7];
    ele[0][9] != ele[3][8];
    ele[0][9] != ele[3][9];
    ele[0][9] != ele[4][5];
    ele[0][9] != ele[4][6];
    ele[0][9] != ele[4][7];
    ele[0][9] != ele[4][8];
    ele[0][9] != ele[4][9];
    ele[0][9] != ele[5][9];
    ele[0][9] != ele[6][9];
    ele[0][9] != ele[7][9];
    ele[0][9] != ele[8][9];
    ele[0][9] != ele[9][9];
    ele[1][0] != ele[1][1];
    ele[1][0] != ele[1][10];
    ele[1][0] != ele[1][11];
    ele[1][0] != ele[1][12];
    ele[1][0] != ele[1][13];
    ele[1][0] != ele[1][14];
    ele[1][0] != ele[1][15];
    ele[1][0] != ele[1][16];
    ele[1][0] != ele[1][17];
    ele[1][0] != ele[1][18];
    ele[1][0] != ele[1][19];
    ele[1][0] != ele[1][2];
    ele[1][0] != ele[1][20];
    ele[1][0] != ele[1][21];
    ele[1][0] != ele[1][22];
    ele[1][0] != ele[1][23];
    ele[1][0] != ele[1][24];
    ele[1][0] != ele[1][3];
    ele[1][0] != ele[1][4];
    ele[1][0] != ele[1][5];
    ele[1][0] != ele[1][6];
    ele[1][0] != ele[1][7];
    ele[1][0] != ele[1][8];
    ele[1][0] != ele[1][9];
    ele[1][0] != ele[10][0];
    ele[1][0] != ele[11][0];
    ele[1][0] != ele[12][0];
    ele[1][0] != ele[13][0];
    ele[1][0] != ele[14][0];
    ele[1][0] != ele[15][0];
    ele[1][0] != ele[16][0];
    ele[1][0] != ele[17][0];
    ele[1][0] != ele[18][0];
    ele[1][0] != ele[19][0];
    ele[1][0] != ele[2][0];
    ele[1][0] != ele[2][1];
    ele[1][0] != ele[2][2];
    ele[1][0] != ele[2][3];
    ele[1][0] != ele[2][4];
    ele[1][0] != ele[20][0];
    ele[1][0] != ele[21][0];
    ele[1][0] != ele[22][0];
    ele[1][0] != ele[23][0];
    ele[1][0] != ele[24][0];
    ele[1][0] != ele[3][0];
    ele[1][0] != ele[3][1];
    ele[1][0] != ele[3][2];
    ele[1][0] != ele[3][3];
    ele[1][0] != ele[3][4];
    ele[1][0] != ele[4][0];
    ele[1][0] != ele[4][1];
    ele[1][0] != ele[4][2];
    ele[1][0] != ele[4][3];
    ele[1][0] != ele[4][4];
    ele[1][0] != ele[5][0];
    ele[1][0] != ele[6][0];
    ele[1][0] != ele[7][0];
    ele[1][0] != ele[8][0];
    ele[1][0] != ele[9][0];
    ele[1][1] != ele[1][10];
    ele[1][1] != ele[1][11];
    ele[1][1] != ele[1][12];
    ele[1][1] != ele[1][13];
    ele[1][1] != ele[1][14];
    ele[1][1] != ele[1][15];
    ele[1][1] != ele[1][16];
    ele[1][1] != ele[1][17];
    ele[1][1] != ele[1][18];
    ele[1][1] != ele[1][19];
    ele[1][1] != ele[1][2];
    ele[1][1] != ele[1][20];
    ele[1][1] != ele[1][21];
    ele[1][1] != ele[1][22];
    ele[1][1] != ele[1][23];
    ele[1][1] != ele[1][24];
    ele[1][1] != ele[1][3];
    ele[1][1] != ele[1][4];
    ele[1][1] != ele[1][5];
    ele[1][1] != ele[1][6];
    ele[1][1] != ele[1][7];
    ele[1][1] != ele[1][8];
    ele[1][1] != ele[1][9];
    ele[1][1] != ele[10][1];
    ele[1][1] != ele[11][1];
    ele[1][1] != ele[12][1];
    ele[1][1] != ele[13][1];
    ele[1][1] != ele[14][1];
    ele[1][1] != ele[15][1];
    ele[1][1] != ele[16][1];
    ele[1][1] != ele[17][1];
    ele[1][1] != ele[18][1];
    ele[1][1] != ele[19][1];
    ele[1][1] != ele[2][0];
    ele[1][1] != ele[2][1];
    ele[1][1] != ele[2][2];
    ele[1][1] != ele[2][3];
    ele[1][1] != ele[2][4];
    ele[1][1] != ele[20][1];
    ele[1][1] != ele[21][1];
    ele[1][1] != ele[22][1];
    ele[1][1] != ele[23][1];
    ele[1][1] != ele[24][1];
    ele[1][1] != ele[3][0];
    ele[1][1] != ele[3][1];
    ele[1][1] != ele[3][2];
    ele[1][1] != ele[3][3];
    ele[1][1] != ele[3][4];
    ele[1][1] != ele[4][0];
    ele[1][1] != ele[4][1];
    ele[1][1] != ele[4][2];
    ele[1][1] != ele[4][3];
    ele[1][1] != ele[4][4];
    ele[1][1] != ele[5][1];
    ele[1][1] != ele[6][1];
    ele[1][1] != ele[7][1];
    ele[1][1] != ele[8][1];
    ele[1][1] != ele[9][1];
    ele[1][10] != ele[1][11];
    ele[1][10] != ele[1][12];
    ele[1][10] != ele[1][13];
    ele[1][10] != ele[1][14];
    ele[1][10] != ele[1][15];
    ele[1][10] != ele[1][16];
    ele[1][10] != ele[1][17];
    ele[1][10] != ele[1][18];
    ele[1][10] != ele[1][19];
    ele[1][10] != ele[1][20];
    ele[1][10] != ele[1][21];
    ele[1][10] != ele[1][22];
    ele[1][10] != ele[1][23];
    ele[1][10] != ele[1][24];
    ele[1][10] != ele[10][10];
    ele[1][10] != ele[11][10];
    ele[1][10] != ele[12][10];
    ele[1][10] != ele[13][10];
    ele[1][10] != ele[14][10];
    ele[1][10] != ele[15][10];
    ele[1][10] != ele[16][10];
    ele[1][10] != ele[17][10];
    ele[1][10] != ele[18][10];
    ele[1][10] != ele[19][10];
    ele[1][10] != ele[2][10];
    ele[1][10] != ele[2][11];
    ele[1][10] != ele[2][12];
    ele[1][10] != ele[2][13];
    ele[1][10] != ele[2][14];
    ele[1][10] != ele[20][10];
    ele[1][10] != ele[21][10];
    ele[1][10] != ele[22][10];
    ele[1][10] != ele[23][10];
    ele[1][10] != ele[24][10];
    ele[1][10] != ele[3][10];
    ele[1][10] != ele[3][11];
    ele[1][10] != ele[3][12];
    ele[1][10] != ele[3][13];
    ele[1][10] != ele[3][14];
    ele[1][10] != ele[4][10];
    ele[1][10] != ele[4][11];
    ele[1][10] != ele[4][12];
    ele[1][10] != ele[4][13];
    ele[1][10] != ele[4][14];
    ele[1][10] != ele[5][10];
    ele[1][10] != ele[6][10];
    ele[1][10] != ele[7][10];
    ele[1][10] != ele[8][10];
    ele[1][10] != ele[9][10];
    ele[1][11] != ele[1][12];
    ele[1][11] != ele[1][13];
    ele[1][11] != ele[1][14];
    ele[1][11] != ele[1][15];
    ele[1][11] != ele[1][16];
    ele[1][11] != ele[1][17];
    ele[1][11] != ele[1][18];
    ele[1][11] != ele[1][19];
    ele[1][11] != ele[1][20];
    ele[1][11] != ele[1][21];
    ele[1][11] != ele[1][22];
    ele[1][11] != ele[1][23];
    ele[1][11] != ele[1][24];
    ele[1][11] != ele[10][11];
    ele[1][11] != ele[11][11];
    ele[1][11] != ele[12][11];
    ele[1][11] != ele[13][11];
    ele[1][11] != ele[14][11];
    ele[1][11] != ele[15][11];
    ele[1][11] != ele[16][11];
    ele[1][11] != ele[17][11];
    ele[1][11] != ele[18][11];
    ele[1][11] != ele[19][11];
    ele[1][11] != ele[2][10];
    ele[1][11] != ele[2][11];
    ele[1][11] != ele[2][12];
    ele[1][11] != ele[2][13];
    ele[1][11] != ele[2][14];
    ele[1][11] != ele[20][11];
    ele[1][11] != ele[21][11];
    ele[1][11] != ele[22][11];
    ele[1][11] != ele[23][11];
    ele[1][11] != ele[24][11];
    ele[1][11] != ele[3][10];
    ele[1][11] != ele[3][11];
    ele[1][11] != ele[3][12];
    ele[1][11] != ele[3][13];
    ele[1][11] != ele[3][14];
    ele[1][11] != ele[4][10];
    ele[1][11] != ele[4][11];
    ele[1][11] != ele[4][12];
    ele[1][11] != ele[4][13];
    ele[1][11] != ele[4][14];
    ele[1][11] != ele[5][11];
    ele[1][11] != ele[6][11];
    ele[1][11] != ele[7][11];
    ele[1][11] != ele[8][11];
    ele[1][11] != ele[9][11];
    ele[1][12] != ele[1][13];
    ele[1][12] != ele[1][14];
    ele[1][12] != ele[1][15];
    ele[1][12] != ele[1][16];
    ele[1][12] != ele[1][17];
    ele[1][12] != ele[1][18];
    ele[1][12] != ele[1][19];
    ele[1][12] != ele[1][20];
    ele[1][12] != ele[1][21];
    ele[1][12] != ele[1][22];
    ele[1][12] != ele[1][23];
    ele[1][12] != ele[1][24];
    ele[1][12] != ele[10][12];
    ele[1][12] != ele[11][12];
    ele[1][12] != ele[12][12];
    ele[1][12] != ele[13][12];
    ele[1][12] != ele[14][12];
    ele[1][12] != ele[15][12];
    ele[1][12] != ele[16][12];
    ele[1][12] != ele[17][12];
    ele[1][12] != ele[18][12];
    ele[1][12] != ele[19][12];
    ele[1][12] != ele[2][10];
    ele[1][12] != ele[2][11];
    ele[1][12] != ele[2][12];
    ele[1][12] != ele[2][13];
    ele[1][12] != ele[2][14];
    ele[1][12] != ele[20][12];
    ele[1][12] != ele[21][12];
    ele[1][12] != ele[22][12];
    ele[1][12] != ele[23][12];
    ele[1][12] != ele[24][12];
    ele[1][12] != ele[3][10];
    ele[1][12] != ele[3][11];
    ele[1][12] != ele[3][12];
    ele[1][12] != ele[3][13];
    ele[1][12] != ele[3][14];
    ele[1][12] != ele[4][10];
    ele[1][12] != ele[4][11];
    ele[1][12] != ele[4][12];
    ele[1][12] != ele[4][13];
    ele[1][12] != ele[4][14];
    ele[1][12] != ele[5][12];
    ele[1][12] != ele[6][12];
    ele[1][12] != ele[7][12];
    ele[1][12] != ele[8][12];
    ele[1][12] != ele[9][12];
    ele[1][13] != ele[1][14];
    ele[1][13] != ele[1][15];
    ele[1][13] != ele[1][16];
    ele[1][13] != ele[1][17];
    ele[1][13] != ele[1][18];
    ele[1][13] != ele[1][19];
    ele[1][13] != ele[1][20];
    ele[1][13] != ele[1][21];
    ele[1][13] != ele[1][22];
    ele[1][13] != ele[1][23];
    ele[1][13] != ele[1][24];
    ele[1][13] != ele[10][13];
    ele[1][13] != ele[11][13];
    ele[1][13] != ele[12][13];
    ele[1][13] != ele[13][13];
    ele[1][13] != ele[14][13];
    ele[1][13] != ele[15][13];
    ele[1][13] != ele[16][13];
    ele[1][13] != ele[17][13];
    ele[1][13] != ele[18][13];
    ele[1][13] != ele[19][13];
    ele[1][13] != ele[2][10];
    ele[1][13] != ele[2][11];
    ele[1][13] != ele[2][12];
    ele[1][13] != ele[2][13];
    ele[1][13] != ele[2][14];
    ele[1][13] != ele[20][13];
    ele[1][13] != ele[21][13];
    ele[1][13] != ele[22][13];
    ele[1][13] != ele[23][13];
    ele[1][13] != ele[24][13];
    ele[1][13] != ele[3][10];
    ele[1][13] != ele[3][11];
    ele[1][13] != ele[3][12];
    ele[1][13] != ele[3][13];
    ele[1][13] != ele[3][14];
    ele[1][13] != ele[4][10];
    ele[1][13] != ele[4][11];
    ele[1][13] != ele[4][12];
    ele[1][13] != ele[4][13];
    ele[1][13] != ele[4][14];
    ele[1][13] != ele[5][13];
    ele[1][13] != ele[6][13];
    ele[1][13] != ele[7][13];
    ele[1][13] != ele[8][13];
    ele[1][13] != ele[9][13];
    ele[1][14] != ele[1][15];
    ele[1][14] != ele[1][16];
    ele[1][14] != ele[1][17];
    ele[1][14] != ele[1][18];
    ele[1][14] != ele[1][19];
    ele[1][14] != ele[1][20];
    ele[1][14] != ele[1][21];
    ele[1][14] != ele[1][22];
    ele[1][14] != ele[1][23];
    ele[1][14] != ele[1][24];
    ele[1][14] != ele[10][14];
    ele[1][14] != ele[11][14];
    ele[1][14] != ele[12][14];
    ele[1][14] != ele[13][14];
    ele[1][14] != ele[14][14];
    ele[1][14] != ele[15][14];
    ele[1][14] != ele[16][14];
    ele[1][14] != ele[17][14];
    ele[1][14] != ele[18][14];
    ele[1][14] != ele[19][14];
    ele[1][14] != ele[2][10];
    ele[1][14] != ele[2][11];
    ele[1][14] != ele[2][12];
    ele[1][14] != ele[2][13];
    ele[1][14] != ele[2][14];
    ele[1][14] != ele[20][14];
    ele[1][14] != ele[21][14];
    ele[1][14] != ele[22][14];
    ele[1][14] != ele[23][14];
    ele[1][14] != ele[24][14];
    ele[1][14] != ele[3][10];
    ele[1][14] != ele[3][11];
    ele[1][14] != ele[3][12];
    ele[1][14] != ele[3][13];
    ele[1][14] != ele[3][14];
    ele[1][14] != ele[4][10];
    ele[1][14] != ele[4][11];
    ele[1][14] != ele[4][12];
    ele[1][14] != ele[4][13];
    ele[1][14] != ele[4][14];
    ele[1][14] != ele[5][14];
    ele[1][14] != ele[6][14];
    ele[1][14] != ele[7][14];
    ele[1][14] != ele[8][14];
    ele[1][14] != ele[9][14];
    ele[1][15] != ele[1][16];
    ele[1][15] != ele[1][17];
    ele[1][15] != ele[1][18];
    ele[1][15] != ele[1][19];
    ele[1][15] != ele[1][20];
    ele[1][15] != ele[1][21];
    ele[1][15] != ele[1][22];
    ele[1][15] != ele[1][23];
    ele[1][15] != ele[1][24];
    ele[1][15] != ele[10][15];
    ele[1][15] != ele[11][15];
    ele[1][15] != ele[12][15];
    ele[1][15] != ele[13][15];
    ele[1][15] != ele[14][15];
    ele[1][15] != ele[15][15];
    ele[1][15] != ele[16][15];
    ele[1][15] != ele[17][15];
    ele[1][15] != ele[18][15];
    ele[1][15] != ele[19][15];
    ele[1][15] != ele[2][15];
    ele[1][15] != ele[2][16];
    ele[1][15] != ele[2][17];
    ele[1][15] != ele[2][18];
    ele[1][15] != ele[2][19];
    ele[1][15] != ele[20][15];
    ele[1][15] != ele[21][15];
    ele[1][15] != ele[22][15];
    ele[1][15] != ele[23][15];
    ele[1][15] != ele[24][15];
    ele[1][15] != ele[3][15];
    ele[1][15] != ele[3][16];
    ele[1][15] != ele[3][17];
    ele[1][15] != ele[3][18];
    ele[1][15] != ele[3][19];
    ele[1][15] != ele[4][15];
    ele[1][15] != ele[4][16];
    ele[1][15] != ele[4][17];
    ele[1][15] != ele[4][18];
    ele[1][15] != ele[4][19];
    ele[1][15] != ele[5][15];
    ele[1][15] != ele[6][15];
    ele[1][15] != ele[7][15];
    ele[1][15] != ele[8][15];
    ele[1][15] != ele[9][15];
    ele[1][16] != ele[1][17];
    ele[1][16] != ele[1][18];
    ele[1][16] != ele[1][19];
    ele[1][16] != ele[1][20];
    ele[1][16] != ele[1][21];
    ele[1][16] != ele[1][22];
    ele[1][16] != ele[1][23];
    ele[1][16] != ele[1][24];
    ele[1][16] != ele[10][16];
    ele[1][16] != ele[11][16];
    ele[1][16] != ele[12][16];
    ele[1][16] != ele[13][16];
    ele[1][16] != ele[14][16];
    ele[1][16] != ele[15][16];
    ele[1][16] != ele[16][16];
    ele[1][16] != ele[17][16];
    ele[1][16] != ele[18][16];
    ele[1][16] != ele[19][16];
    ele[1][16] != ele[2][15];
    ele[1][16] != ele[2][16];
    ele[1][16] != ele[2][17];
    ele[1][16] != ele[2][18];
    ele[1][16] != ele[2][19];
    ele[1][16] != ele[20][16];
    ele[1][16] != ele[21][16];
    ele[1][16] != ele[22][16];
    ele[1][16] != ele[23][16];
    ele[1][16] != ele[24][16];
    ele[1][16] != ele[3][15];
    ele[1][16] != ele[3][16];
    ele[1][16] != ele[3][17];
    ele[1][16] != ele[3][18];
    ele[1][16] != ele[3][19];
    ele[1][16] != ele[4][15];
    ele[1][16] != ele[4][16];
    ele[1][16] != ele[4][17];
    ele[1][16] != ele[4][18];
    ele[1][16] != ele[4][19];
    ele[1][16] != ele[5][16];
    ele[1][16] != ele[6][16];
    ele[1][16] != ele[7][16];
    ele[1][16] != ele[8][16];
    ele[1][16] != ele[9][16];
    ele[1][17] != ele[1][18];
    ele[1][17] != ele[1][19];
    ele[1][17] != ele[1][20];
    ele[1][17] != ele[1][21];
    ele[1][17] != ele[1][22];
    ele[1][17] != ele[1][23];
    ele[1][17] != ele[1][24];
    ele[1][17] != ele[10][17];
    ele[1][17] != ele[11][17];
    ele[1][17] != ele[12][17];
    ele[1][17] != ele[13][17];
    ele[1][17] != ele[14][17];
    ele[1][17] != ele[15][17];
    ele[1][17] != ele[16][17];
    ele[1][17] != ele[17][17];
    ele[1][17] != ele[18][17];
    ele[1][17] != ele[19][17];
    ele[1][17] != ele[2][15];
    ele[1][17] != ele[2][16];
    ele[1][17] != ele[2][17];
    ele[1][17] != ele[2][18];
    ele[1][17] != ele[2][19];
    ele[1][17] != ele[20][17];
    ele[1][17] != ele[21][17];
    ele[1][17] != ele[22][17];
    ele[1][17] != ele[23][17];
    ele[1][17] != ele[24][17];
    ele[1][17] != ele[3][15];
    ele[1][17] != ele[3][16];
    ele[1][17] != ele[3][17];
    ele[1][17] != ele[3][18];
    ele[1][17] != ele[3][19];
    ele[1][17] != ele[4][15];
    ele[1][17] != ele[4][16];
    ele[1][17] != ele[4][17];
    ele[1][17] != ele[4][18];
    ele[1][17] != ele[4][19];
    ele[1][17] != ele[5][17];
    ele[1][17] != ele[6][17];
    ele[1][17] != ele[7][17];
    ele[1][17] != ele[8][17];
    ele[1][17] != ele[9][17];
    ele[1][18] != ele[1][19];
    ele[1][18] != ele[1][20];
    ele[1][18] != ele[1][21];
    ele[1][18] != ele[1][22];
    ele[1][18] != ele[1][23];
    ele[1][18] != ele[1][24];
    ele[1][18] != ele[10][18];
    ele[1][18] != ele[11][18];
    ele[1][18] != ele[12][18];
    ele[1][18] != ele[13][18];
    ele[1][18] != ele[14][18];
    ele[1][18] != ele[15][18];
    ele[1][18] != ele[16][18];
    ele[1][18] != ele[17][18];
    ele[1][18] != ele[18][18];
    ele[1][18] != ele[19][18];
    ele[1][18] != ele[2][15];
    ele[1][18] != ele[2][16];
    ele[1][18] != ele[2][17];
    ele[1][18] != ele[2][18];
    ele[1][18] != ele[2][19];
    ele[1][18] != ele[20][18];
    ele[1][18] != ele[21][18];
    ele[1][18] != ele[22][18];
    ele[1][18] != ele[23][18];
    ele[1][18] != ele[24][18];
    ele[1][18] != ele[3][15];
    ele[1][18] != ele[3][16];
    ele[1][18] != ele[3][17];
    ele[1][18] != ele[3][18];
    ele[1][18] != ele[3][19];
    ele[1][18] != ele[4][15];
    ele[1][18] != ele[4][16];
    ele[1][18] != ele[4][17];
    ele[1][18] != ele[4][18];
    ele[1][18] != ele[4][19];
    ele[1][18] != ele[5][18];
    ele[1][18] != ele[6][18];
    ele[1][18] != ele[7][18];
    ele[1][18] != ele[8][18];
    ele[1][18] != ele[9][18];
    ele[1][19] != ele[1][20];
    ele[1][19] != ele[1][21];
    ele[1][19] != ele[1][22];
    ele[1][19] != ele[1][23];
    ele[1][19] != ele[1][24];
    ele[1][19] != ele[10][19];
    ele[1][19] != ele[11][19];
    ele[1][19] != ele[12][19];
    ele[1][19] != ele[13][19];
    ele[1][19] != ele[14][19];
    ele[1][19] != ele[15][19];
    ele[1][19] != ele[16][19];
    ele[1][19] != ele[17][19];
    ele[1][19] != ele[18][19];
    ele[1][19] != ele[19][19];
    ele[1][19] != ele[2][15];
    ele[1][19] != ele[2][16];
    ele[1][19] != ele[2][17];
    ele[1][19] != ele[2][18];
    ele[1][19] != ele[2][19];
    ele[1][19] != ele[20][19];
    ele[1][19] != ele[21][19];
    ele[1][19] != ele[22][19];
    ele[1][19] != ele[23][19];
    ele[1][19] != ele[24][19];
    ele[1][19] != ele[3][15];
    ele[1][19] != ele[3][16];
    ele[1][19] != ele[3][17];
    ele[1][19] != ele[3][18];
    ele[1][19] != ele[3][19];
    ele[1][19] != ele[4][15];
    ele[1][19] != ele[4][16];
    ele[1][19] != ele[4][17];
    ele[1][19] != ele[4][18];
    ele[1][19] != ele[4][19];
    ele[1][19] != ele[5][19];
    ele[1][19] != ele[6][19];
    ele[1][19] != ele[7][19];
    ele[1][19] != ele[8][19];
    ele[1][19] != ele[9][19];
    ele[1][2] != ele[1][10];
    ele[1][2] != ele[1][11];
    ele[1][2] != ele[1][12];
    ele[1][2] != ele[1][13];
    ele[1][2] != ele[1][14];
    ele[1][2] != ele[1][15];
    ele[1][2] != ele[1][16];
    ele[1][2] != ele[1][17];
    ele[1][2] != ele[1][18];
    ele[1][2] != ele[1][19];
    ele[1][2] != ele[1][20];
    ele[1][2] != ele[1][21];
    ele[1][2] != ele[1][22];
    ele[1][2] != ele[1][23];
    ele[1][2] != ele[1][24];
    ele[1][2] != ele[1][3];
    ele[1][2] != ele[1][4];
    ele[1][2] != ele[1][5];
    ele[1][2] != ele[1][6];
    ele[1][2] != ele[1][7];
    ele[1][2] != ele[1][8];
    ele[1][2] != ele[1][9];
    ele[1][2] != ele[10][2];
    ele[1][2] != ele[11][2];
    ele[1][2] != ele[12][2];
    ele[1][2] != ele[13][2];
    ele[1][2] != ele[14][2];
    ele[1][2] != ele[15][2];
    ele[1][2] != ele[16][2];
    ele[1][2] != ele[17][2];
    ele[1][2] != ele[18][2];
    ele[1][2] != ele[19][2];
    ele[1][2] != ele[2][0];
    ele[1][2] != ele[2][1];
    ele[1][2] != ele[2][2];
    ele[1][2] != ele[2][3];
    ele[1][2] != ele[2][4];
    ele[1][2] != ele[20][2];
    ele[1][2] != ele[21][2];
    ele[1][2] != ele[22][2];
    ele[1][2] != ele[23][2];
    ele[1][2] != ele[24][2];
    ele[1][2] != ele[3][0];
    ele[1][2] != ele[3][1];
    ele[1][2] != ele[3][2];
    ele[1][2] != ele[3][3];
    ele[1][2] != ele[3][4];
    ele[1][2] != ele[4][0];
    ele[1][2] != ele[4][1];
    ele[1][2] != ele[4][2];
    ele[1][2] != ele[4][3];
    ele[1][2] != ele[4][4];
    ele[1][2] != ele[5][2];
    ele[1][2] != ele[6][2];
    ele[1][2] != ele[7][2];
    ele[1][2] != ele[8][2];
    ele[1][2] != ele[9][2];
    ele[1][20] != ele[1][21];
    ele[1][20] != ele[1][22];
    ele[1][20] != ele[1][23];
    ele[1][20] != ele[1][24];
    ele[1][20] != ele[10][20];
    ele[1][20] != ele[11][20];
    ele[1][20] != ele[12][20];
    ele[1][20] != ele[13][20];
    ele[1][20] != ele[14][20];
    ele[1][20] != ele[15][20];
    ele[1][20] != ele[16][20];
    ele[1][20] != ele[17][20];
    ele[1][20] != ele[18][20];
    ele[1][20] != ele[19][20];
    ele[1][20] != ele[2][20];
    ele[1][20] != ele[2][21];
    ele[1][20] != ele[2][22];
    ele[1][20] != ele[2][23];
    ele[1][20] != ele[2][24];
    ele[1][20] != ele[20][20];
    ele[1][20] != ele[21][20];
    ele[1][20] != ele[22][20];
    ele[1][20] != ele[23][20];
    ele[1][20] != ele[24][20];
    ele[1][20] != ele[3][20];
    ele[1][20] != ele[3][21];
    ele[1][20] != ele[3][22];
    ele[1][20] != ele[3][23];
    ele[1][20] != ele[3][24];
    ele[1][20] != ele[4][20];
    ele[1][20] != ele[4][21];
    ele[1][20] != ele[4][22];
    ele[1][20] != ele[4][23];
    ele[1][20] != ele[4][24];
    ele[1][20] != ele[5][20];
    ele[1][20] != ele[6][20];
    ele[1][20] != ele[7][20];
    ele[1][20] != ele[8][20];
    ele[1][20] != ele[9][20];
    ele[1][21] != ele[1][22];
    ele[1][21] != ele[1][23];
    ele[1][21] != ele[1][24];
    ele[1][21] != ele[10][21];
    ele[1][21] != ele[11][21];
    ele[1][21] != ele[12][21];
    ele[1][21] != ele[13][21];
    ele[1][21] != ele[14][21];
    ele[1][21] != ele[15][21];
    ele[1][21] != ele[16][21];
    ele[1][21] != ele[17][21];
    ele[1][21] != ele[18][21];
    ele[1][21] != ele[19][21];
    ele[1][21] != ele[2][20];
    ele[1][21] != ele[2][21];
    ele[1][21] != ele[2][22];
    ele[1][21] != ele[2][23];
    ele[1][21] != ele[2][24];
    ele[1][21] != ele[20][21];
    ele[1][21] != ele[21][21];
    ele[1][21] != ele[22][21];
    ele[1][21] != ele[23][21];
    ele[1][21] != ele[24][21];
    ele[1][21] != ele[3][20];
    ele[1][21] != ele[3][21];
    ele[1][21] != ele[3][22];
    ele[1][21] != ele[3][23];
    ele[1][21] != ele[3][24];
    ele[1][21] != ele[4][20];
    ele[1][21] != ele[4][21];
    ele[1][21] != ele[4][22];
    ele[1][21] != ele[4][23];
    ele[1][21] != ele[4][24];
    ele[1][21] != ele[5][21];
    ele[1][21] != ele[6][21];
    ele[1][21] != ele[7][21];
    ele[1][21] != ele[8][21];
    ele[1][21] != ele[9][21];
    ele[1][22] != ele[1][23];
    ele[1][22] != ele[1][24];
    ele[1][22] != ele[10][22];
    ele[1][22] != ele[11][22];
    ele[1][22] != ele[12][22];
    ele[1][22] != ele[13][22];
    ele[1][22] != ele[14][22];
    ele[1][22] != ele[15][22];
    ele[1][22] != ele[16][22];
    ele[1][22] != ele[17][22];
    ele[1][22] != ele[18][22];
    ele[1][22] != ele[19][22];
    ele[1][22] != ele[2][20];
    ele[1][22] != ele[2][21];
    ele[1][22] != ele[2][22];
    ele[1][22] != ele[2][23];
    ele[1][22] != ele[2][24];
    ele[1][22] != ele[20][22];
    ele[1][22] != ele[21][22];
    ele[1][22] != ele[22][22];
    ele[1][22] != ele[23][22];
    ele[1][22] != ele[24][22];
    ele[1][22] != ele[3][20];
    ele[1][22] != ele[3][21];
    ele[1][22] != ele[3][22];
    ele[1][22] != ele[3][23];
    ele[1][22] != ele[3][24];
    ele[1][22] != ele[4][20];
    ele[1][22] != ele[4][21];
    ele[1][22] != ele[4][22];
    ele[1][22] != ele[4][23];
    ele[1][22] != ele[4][24];
    ele[1][22] != ele[5][22];
    ele[1][22] != ele[6][22];
    ele[1][22] != ele[7][22];
    ele[1][22] != ele[8][22];
    ele[1][22] != ele[9][22];
    ele[1][23] != ele[1][24];
    ele[1][23] != ele[10][23];
    ele[1][23] != ele[11][23];
    ele[1][23] != ele[12][23];
    ele[1][23] != ele[13][23];
    ele[1][23] != ele[14][23];
    ele[1][23] != ele[15][23];
    ele[1][23] != ele[16][23];
    ele[1][23] != ele[17][23];
    ele[1][23] != ele[18][23];
    ele[1][23] != ele[19][23];
    ele[1][23] != ele[2][20];
    ele[1][23] != ele[2][21];
    ele[1][23] != ele[2][22];
    ele[1][23] != ele[2][23];
    ele[1][23] != ele[2][24];
    ele[1][23] != ele[20][23];
    ele[1][23] != ele[21][23];
    ele[1][23] != ele[22][23];
    ele[1][23] != ele[23][23];
    ele[1][23] != ele[24][23];
    ele[1][23] != ele[3][20];
    ele[1][23] != ele[3][21];
    ele[1][23] != ele[3][22];
    ele[1][23] != ele[3][23];
    ele[1][23] != ele[3][24];
    ele[1][23] != ele[4][20];
    ele[1][23] != ele[4][21];
    ele[1][23] != ele[4][22];
    ele[1][23] != ele[4][23];
    ele[1][23] != ele[4][24];
    ele[1][23] != ele[5][23];
    ele[1][23] != ele[6][23];
    ele[1][23] != ele[7][23];
    ele[1][23] != ele[8][23];
    ele[1][23] != ele[9][23];
    ele[1][24] != ele[10][24];
    ele[1][24] != ele[11][24];
    ele[1][24] != ele[12][24];
    ele[1][24] != ele[13][24];
    ele[1][24] != ele[14][24];
    ele[1][24] != ele[15][24];
    ele[1][24] != ele[16][24];
    ele[1][24] != ele[17][24];
    ele[1][24] != ele[18][24];
    ele[1][24] != ele[19][24];
    ele[1][24] != ele[2][20];
    ele[1][24] != ele[2][21];
    ele[1][24] != ele[2][22];
    ele[1][24] != ele[2][23];
    ele[1][24] != ele[2][24];
    ele[1][24] != ele[20][24];
    ele[1][24] != ele[21][24];
    ele[1][24] != ele[22][24];
    ele[1][24] != ele[23][24];
    ele[1][24] != ele[24][24];
    ele[1][24] != ele[3][20];
    ele[1][24] != ele[3][21];
    ele[1][24] != ele[3][22];
    ele[1][24] != ele[3][23];
    ele[1][24] != ele[3][24];
    ele[1][24] != ele[4][20];
    ele[1][24] != ele[4][21];
    ele[1][24] != ele[4][22];
    ele[1][24] != ele[4][23];
    ele[1][24] != ele[4][24];
    ele[1][24] != ele[5][24];
    ele[1][24] != ele[6][24];
    ele[1][24] != ele[7][24];
    ele[1][24] != ele[8][24];
    ele[1][24] != ele[9][24];
    ele[1][3] != ele[1][10];
    ele[1][3] != ele[1][11];
    ele[1][3] != ele[1][12];
    ele[1][3] != ele[1][13];
    ele[1][3] != ele[1][14];
    ele[1][3] != ele[1][15];
    ele[1][3] != ele[1][16];
    ele[1][3] != ele[1][17];
    ele[1][3] != ele[1][18];
    ele[1][3] != ele[1][19];
    ele[1][3] != ele[1][20];
    ele[1][3] != ele[1][21];
    ele[1][3] != ele[1][22];
    ele[1][3] != ele[1][23];
    ele[1][3] != ele[1][24];
    ele[1][3] != ele[1][4];
    ele[1][3] != ele[1][5];
    ele[1][3] != ele[1][6];
    ele[1][3] != ele[1][7];
    ele[1][3] != ele[1][8];
    ele[1][3] != ele[1][9];
    ele[1][3] != ele[10][3];
    ele[1][3] != ele[11][3];
    ele[1][3] != ele[12][3];
    ele[1][3] != ele[13][3];
    ele[1][3] != ele[14][3];
    ele[1][3] != ele[15][3];
    ele[1][3] != ele[16][3];
    ele[1][3] != ele[17][3];
    ele[1][3] != ele[18][3];
    ele[1][3] != ele[19][3];
    ele[1][3] != ele[2][0];
    ele[1][3] != ele[2][1];
    ele[1][3] != ele[2][2];
    ele[1][3] != ele[2][3];
    ele[1][3] != ele[2][4];
    ele[1][3] != ele[20][3];
    ele[1][3] != ele[21][3];
    ele[1][3] != ele[22][3];
    ele[1][3] != ele[23][3];
    ele[1][3] != ele[24][3];
    ele[1][3] != ele[3][0];
    ele[1][3] != ele[3][1];
    ele[1][3] != ele[3][2];
    ele[1][3] != ele[3][3];
    ele[1][3] != ele[3][4];
    ele[1][3] != ele[4][0];
    ele[1][3] != ele[4][1];
    ele[1][3] != ele[4][2];
    ele[1][3] != ele[4][3];
    ele[1][3] != ele[4][4];
    ele[1][3] != ele[5][3];
    ele[1][3] != ele[6][3];
    ele[1][3] != ele[7][3];
    ele[1][3] != ele[8][3];
    ele[1][3] != ele[9][3];
    ele[1][4] != ele[1][10];
    ele[1][4] != ele[1][11];
    ele[1][4] != ele[1][12];
    ele[1][4] != ele[1][13];
    ele[1][4] != ele[1][14];
    ele[1][4] != ele[1][15];
    ele[1][4] != ele[1][16];
    ele[1][4] != ele[1][17];
    ele[1][4] != ele[1][18];
    ele[1][4] != ele[1][19];
    ele[1][4] != ele[1][20];
    ele[1][4] != ele[1][21];
    ele[1][4] != ele[1][22];
    ele[1][4] != ele[1][23];
    ele[1][4] != ele[1][24];
    ele[1][4] != ele[1][5];
    ele[1][4] != ele[1][6];
    ele[1][4] != ele[1][7];
    ele[1][4] != ele[1][8];
    ele[1][4] != ele[1][9];
    ele[1][4] != ele[10][4];
    ele[1][4] != ele[11][4];
    ele[1][4] != ele[12][4];
    ele[1][4] != ele[13][4];
    ele[1][4] != ele[14][4];
    ele[1][4] != ele[15][4];
    ele[1][4] != ele[16][4];
    ele[1][4] != ele[17][4];
    ele[1][4] != ele[18][4];
    ele[1][4] != ele[19][4];
    ele[1][4] != ele[2][0];
    ele[1][4] != ele[2][1];
    ele[1][4] != ele[2][2];
    ele[1][4] != ele[2][3];
    ele[1][4] != ele[2][4];
    ele[1][4] != ele[20][4];
    ele[1][4] != ele[21][4];
    ele[1][4] != ele[22][4];
    ele[1][4] != ele[23][4];
    ele[1][4] != ele[24][4];
    ele[1][4] != ele[3][0];
    ele[1][4] != ele[3][1];
    ele[1][4] != ele[3][2];
    ele[1][4] != ele[3][3];
    ele[1][4] != ele[3][4];
    ele[1][4] != ele[4][0];
    ele[1][4] != ele[4][1];
    ele[1][4] != ele[4][2];
    ele[1][4] != ele[4][3];
    ele[1][4] != ele[4][4];
    ele[1][4] != ele[5][4];
    ele[1][4] != ele[6][4];
    ele[1][4] != ele[7][4];
    ele[1][4] != ele[8][4];
    ele[1][4] != ele[9][4];
    ele[1][5] != ele[1][10];
    ele[1][5] != ele[1][11];
    ele[1][5] != ele[1][12];
    ele[1][5] != ele[1][13];
    ele[1][5] != ele[1][14];
    ele[1][5] != ele[1][15];
    ele[1][5] != ele[1][16];
    ele[1][5] != ele[1][17];
    ele[1][5] != ele[1][18];
    ele[1][5] != ele[1][19];
    ele[1][5] != ele[1][20];
    ele[1][5] != ele[1][21];
    ele[1][5] != ele[1][22];
    ele[1][5] != ele[1][23];
    ele[1][5] != ele[1][24];
    ele[1][5] != ele[1][6];
    ele[1][5] != ele[1][7];
    ele[1][5] != ele[1][8];
    ele[1][5] != ele[1][9];
    ele[1][5] != ele[10][5];
    ele[1][5] != ele[11][5];
    ele[1][5] != ele[12][5];
    ele[1][5] != ele[13][5];
    ele[1][5] != ele[14][5];
    ele[1][5] != ele[15][5];
    ele[1][5] != ele[16][5];
    ele[1][5] != ele[17][5];
    ele[1][5] != ele[18][5];
    ele[1][5] != ele[19][5];
    ele[1][5] != ele[2][5];
    ele[1][5] != ele[2][6];
    ele[1][5] != ele[2][7];
    ele[1][5] != ele[2][8];
    ele[1][5] != ele[2][9];
    ele[1][5] != ele[20][5];
    ele[1][5] != ele[21][5];
    ele[1][5] != ele[22][5];
    ele[1][5] != ele[23][5];
    ele[1][5] != ele[24][5];
    ele[1][5] != ele[3][5];
    ele[1][5] != ele[3][6];
    ele[1][5] != ele[3][7];
    ele[1][5] != ele[3][8];
    ele[1][5] != ele[3][9];
    ele[1][5] != ele[4][5];
    ele[1][5] != ele[4][6];
    ele[1][5] != ele[4][7];
    ele[1][5] != ele[4][8];
    ele[1][5] != ele[4][9];
    ele[1][5] != ele[5][5];
    ele[1][5] != ele[6][5];
    ele[1][5] != ele[7][5];
    ele[1][5] != ele[8][5];
    ele[1][5] != ele[9][5];
    ele[1][6] != ele[1][10];
    ele[1][6] != ele[1][11];
    ele[1][6] != ele[1][12];
    ele[1][6] != ele[1][13];
    ele[1][6] != ele[1][14];
    ele[1][6] != ele[1][15];
    ele[1][6] != ele[1][16];
    ele[1][6] != ele[1][17];
    ele[1][6] != ele[1][18];
    ele[1][6] != ele[1][19];
    ele[1][6] != ele[1][20];
    ele[1][6] != ele[1][21];
    ele[1][6] != ele[1][22];
    ele[1][6] != ele[1][23];
    ele[1][6] != ele[1][24];
    ele[1][6] != ele[1][7];
    ele[1][6] != ele[1][8];
    ele[1][6] != ele[1][9];
    ele[1][6] != ele[10][6];
    ele[1][6] != ele[11][6];
    ele[1][6] != ele[12][6];
    ele[1][6] != ele[13][6];
    ele[1][6] != ele[14][6];
    ele[1][6] != ele[15][6];
    ele[1][6] != ele[16][6];
    ele[1][6] != ele[17][6];
    ele[1][6] != ele[18][6];
    ele[1][6] != ele[19][6];
    ele[1][6] != ele[2][5];
    ele[1][6] != ele[2][6];
    ele[1][6] != ele[2][7];
    ele[1][6] != ele[2][8];
    ele[1][6] != ele[2][9];
    ele[1][6] != ele[20][6];
    ele[1][6] != ele[21][6];
    ele[1][6] != ele[22][6];
    ele[1][6] != ele[23][6];
    ele[1][6] != ele[24][6];
    ele[1][6] != ele[3][5];
    ele[1][6] != ele[3][6];
    ele[1][6] != ele[3][7];
    ele[1][6] != ele[3][8];
    ele[1][6] != ele[3][9];
    ele[1][6] != ele[4][5];
    ele[1][6] != ele[4][6];
    ele[1][6] != ele[4][7];
    ele[1][6] != ele[4][8];
    ele[1][6] != ele[4][9];
    ele[1][6] != ele[5][6];
    ele[1][6] != ele[6][6];
    ele[1][6] != ele[7][6];
    ele[1][6] != ele[8][6];
    ele[1][6] != ele[9][6];
    ele[1][7] != ele[1][10];
    ele[1][7] != ele[1][11];
    ele[1][7] != ele[1][12];
    ele[1][7] != ele[1][13];
    ele[1][7] != ele[1][14];
    ele[1][7] != ele[1][15];
    ele[1][7] != ele[1][16];
    ele[1][7] != ele[1][17];
    ele[1][7] != ele[1][18];
    ele[1][7] != ele[1][19];
    ele[1][7] != ele[1][20];
    ele[1][7] != ele[1][21];
    ele[1][7] != ele[1][22];
    ele[1][7] != ele[1][23];
    ele[1][7] != ele[1][24];
    ele[1][7] != ele[1][8];
    ele[1][7] != ele[1][9];
    ele[1][7] != ele[10][7];
    ele[1][7] != ele[11][7];
    ele[1][7] != ele[12][7];
    ele[1][7] != ele[13][7];
    ele[1][7] != ele[14][7];
    ele[1][7] != ele[15][7];
    ele[1][7] != ele[16][7];
    ele[1][7] != ele[17][7];
    ele[1][7] != ele[18][7];
    ele[1][7] != ele[19][7];
    ele[1][7] != ele[2][5];
    ele[1][7] != ele[2][6];
    ele[1][7] != ele[2][7];
    ele[1][7] != ele[2][8];
    ele[1][7] != ele[2][9];
    ele[1][7] != ele[20][7];
    ele[1][7] != ele[21][7];
    ele[1][7] != ele[22][7];
    ele[1][7] != ele[23][7];
    ele[1][7] != ele[24][7];
    ele[1][7] != ele[3][5];
    ele[1][7] != ele[3][6];
    ele[1][7] != ele[3][7];
    ele[1][7] != ele[3][8];
    ele[1][7] != ele[3][9];
    ele[1][7] != ele[4][5];
    ele[1][7] != ele[4][6];
    ele[1][7] != ele[4][7];
    ele[1][7] != ele[4][8];
    ele[1][7] != ele[4][9];
    ele[1][7] != ele[5][7];
    ele[1][7] != ele[6][7];
    ele[1][7] != ele[7][7];
    ele[1][7] != ele[8][7];
    ele[1][7] != ele[9][7];
    ele[1][8] != ele[1][10];
    ele[1][8] != ele[1][11];
    ele[1][8] != ele[1][12];
    ele[1][8] != ele[1][13];
    ele[1][8] != ele[1][14];
    ele[1][8] != ele[1][15];
    ele[1][8] != ele[1][16];
    ele[1][8] != ele[1][17];
    ele[1][8] != ele[1][18];
    ele[1][8] != ele[1][19];
    ele[1][8] != ele[1][20];
    ele[1][8] != ele[1][21];
    ele[1][8] != ele[1][22];
    ele[1][8] != ele[1][23];
    ele[1][8] != ele[1][24];
    ele[1][8] != ele[1][9];
    ele[1][8] != ele[10][8];
    ele[1][8] != ele[11][8];
    ele[1][8] != ele[12][8];
    ele[1][8] != ele[13][8];
    ele[1][8] != ele[14][8];
    ele[1][8] != ele[15][8];
    ele[1][8] != ele[16][8];
    ele[1][8] != ele[17][8];
    ele[1][8] != ele[18][8];
    ele[1][8] != ele[19][8];
    ele[1][8] != ele[2][5];
    ele[1][8] != ele[2][6];
    ele[1][8] != ele[2][7];
    ele[1][8] != ele[2][8];
    ele[1][8] != ele[2][9];
    ele[1][8] != ele[20][8];
    ele[1][8] != ele[21][8];
    ele[1][8] != ele[22][8];
    ele[1][8] != ele[23][8];
    ele[1][8] != ele[24][8];
    ele[1][8] != ele[3][5];
    ele[1][8] != ele[3][6];
    ele[1][8] != ele[3][7];
    ele[1][8] != ele[3][8];
    ele[1][8] != ele[3][9];
    ele[1][8] != ele[4][5];
    ele[1][8] != ele[4][6];
    ele[1][8] != ele[4][7];
    ele[1][8] != ele[4][8];
    ele[1][8] != ele[4][9];
    ele[1][8] != ele[5][8];
    ele[1][8] != ele[6][8];
    ele[1][8] != ele[7][8];
    ele[1][8] != ele[8][8];
    ele[1][8] != ele[9][8];
    ele[1][9] != ele[1][10];
    ele[1][9] != ele[1][11];
    ele[1][9] != ele[1][12];
    ele[1][9] != ele[1][13];
    ele[1][9] != ele[1][14];
    ele[1][9] != ele[1][15];
    ele[1][9] != ele[1][16];
    ele[1][9] != ele[1][17];
    ele[1][9] != ele[1][18];
    ele[1][9] != ele[1][19];
    ele[1][9] != ele[1][20];
    ele[1][9] != ele[1][21];
    ele[1][9] != ele[1][22];
    ele[1][9] != ele[1][23];
    ele[1][9] != ele[1][24];
    ele[1][9] != ele[10][9];
    ele[1][9] != ele[11][9];
    ele[1][9] != ele[12][9];
    ele[1][9] != ele[13][9];
    ele[1][9] != ele[14][9];
    ele[1][9] != ele[15][9];
    ele[1][9] != ele[16][9];
    ele[1][9] != ele[17][9];
    ele[1][9] != ele[18][9];
    ele[1][9] != ele[19][9];
    ele[1][9] != ele[2][5];
    ele[1][9] != ele[2][6];
    ele[1][9] != ele[2][7];
    ele[1][9] != ele[2][8];
    ele[1][9] != ele[2][9];
    ele[1][9] != ele[20][9];
    ele[1][9] != ele[21][9];
    ele[1][9] != ele[22][9];
    ele[1][9] != ele[23][9];
    ele[1][9] != ele[24][9];
    ele[1][9] != ele[3][5];
    ele[1][9] != ele[3][6];
    ele[1][9] != ele[3][7];
    ele[1][9] != ele[3][8];
    ele[1][9] != ele[3][9];
    ele[1][9] != ele[4][5];
    ele[1][9] != ele[4][6];
    ele[1][9] != ele[4][7];
    ele[1][9] != ele[4][8];
    ele[1][9] != ele[4][9];
    ele[1][9] != ele[5][9];
    ele[1][9] != ele[6][9];
    ele[1][9] != ele[7][9];
    ele[1][9] != ele[8][9];
    ele[1][9] != ele[9][9];
    ele[10][0] != ele[10][1];
    ele[10][0] != ele[10][10];
    ele[10][0] != ele[10][11];
    ele[10][0] != ele[10][12];
    ele[10][0] != ele[10][13];
    ele[10][0] != ele[10][14];
    ele[10][0] != ele[10][15];
    ele[10][0] != ele[10][16];
    ele[10][0] != ele[10][17];
    ele[10][0] != ele[10][18];
    ele[10][0] != ele[10][19];
    ele[10][0] != ele[10][2];
    ele[10][0] != ele[10][20];
    ele[10][0] != ele[10][21];
    ele[10][0] != ele[10][22];
    ele[10][0] != ele[10][23];
    ele[10][0] != ele[10][24];
    ele[10][0] != ele[10][3];
    ele[10][0] != ele[10][4];
    ele[10][0] != ele[10][5];
    ele[10][0] != ele[10][6];
    ele[10][0] != ele[10][7];
    ele[10][0] != ele[10][8];
    ele[10][0] != ele[10][9];
    ele[10][0] != ele[11][0];
    ele[10][0] != ele[11][1];
    ele[10][0] != ele[11][2];
    ele[10][0] != ele[11][3];
    ele[10][0] != ele[11][4];
    ele[10][0] != ele[12][0];
    ele[10][0] != ele[12][1];
    ele[10][0] != ele[12][2];
    ele[10][0] != ele[12][3];
    ele[10][0] != ele[12][4];
    ele[10][0] != ele[13][0];
    ele[10][0] != ele[13][1];
    ele[10][0] != ele[13][2];
    ele[10][0] != ele[13][3];
    ele[10][0] != ele[13][4];
    ele[10][0] != ele[14][0];
    ele[10][0] != ele[14][1];
    ele[10][0] != ele[14][2];
    ele[10][0] != ele[14][3];
    ele[10][0] != ele[14][4];
    ele[10][0] != ele[15][0];
    ele[10][0] != ele[16][0];
    ele[10][0] != ele[17][0];
    ele[10][0] != ele[18][0];
    ele[10][0] != ele[19][0];
    ele[10][0] != ele[20][0];
    ele[10][0] != ele[21][0];
    ele[10][0] != ele[22][0];
    ele[10][0] != ele[23][0];
    ele[10][0] != ele[24][0];
    ele[10][1] != ele[10][10];
    ele[10][1] != ele[10][11];
    ele[10][1] != ele[10][12];
    ele[10][1] != ele[10][13];
    ele[10][1] != ele[10][14];
    ele[10][1] != ele[10][15];
    ele[10][1] != ele[10][16];
    ele[10][1] != ele[10][17];
    ele[10][1] != ele[10][18];
    ele[10][1] != ele[10][19];
    ele[10][1] != ele[10][2];
    ele[10][1] != ele[10][20];
    ele[10][1] != ele[10][21];
    ele[10][1] != ele[10][22];
    ele[10][1] != ele[10][23];
    ele[10][1] != ele[10][24];
    ele[10][1] != ele[10][3];
    ele[10][1] != ele[10][4];
    ele[10][1] != ele[10][5];
    ele[10][1] != ele[10][6];
    ele[10][1] != ele[10][7];
    ele[10][1] != ele[10][8];
    ele[10][1] != ele[10][9];
    ele[10][1] != ele[11][0];
    ele[10][1] != ele[11][1];
    ele[10][1] != ele[11][2];
    ele[10][1] != ele[11][3];
    ele[10][1] != ele[11][4];
    ele[10][1] != ele[12][0];
    ele[10][1] != ele[12][1];
    ele[10][1] != ele[12][2];
    ele[10][1] != ele[12][3];
    ele[10][1] != ele[12][4];
    ele[10][1] != ele[13][0];
    ele[10][1] != ele[13][1];
    ele[10][1] != ele[13][2];
    ele[10][1] != ele[13][3];
    ele[10][1] != ele[13][4];
    ele[10][1] != ele[14][0];
    ele[10][1] != ele[14][1];
    ele[10][1] != ele[14][2];
    ele[10][1] != ele[14][3];
    ele[10][1] != ele[14][4];
    ele[10][1] != ele[15][1];
    ele[10][1] != ele[16][1];
    ele[10][1] != ele[17][1];
    ele[10][1] != ele[18][1];
    ele[10][1] != ele[19][1];
    ele[10][1] != ele[20][1];
    ele[10][1] != ele[21][1];
    ele[10][1] != ele[22][1];
    ele[10][1] != ele[23][1];
    ele[10][1] != ele[24][1];
    ele[10][10] != ele[10][11];
    ele[10][10] != ele[10][12];
    ele[10][10] != ele[10][13];
    ele[10][10] != ele[10][14];
    ele[10][10] != ele[10][15];
    ele[10][10] != ele[10][16];
    ele[10][10] != ele[10][17];
    ele[10][10] != ele[10][18];
    ele[10][10] != ele[10][19];
    ele[10][10] != ele[10][20];
    ele[10][10] != ele[10][21];
    ele[10][10] != ele[10][22];
    ele[10][10] != ele[10][23];
    ele[10][10] != ele[10][24];
    ele[10][10] != ele[11][10];
    ele[10][10] != ele[11][11];
    ele[10][10] != ele[11][12];
    ele[10][10] != ele[11][13];
    ele[10][10] != ele[11][14];
    ele[10][10] != ele[12][10];
    ele[10][10] != ele[12][11];
    ele[10][10] != ele[12][12];
    ele[10][10] != ele[12][13];
    ele[10][10] != ele[12][14];
    ele[10][10] != ele[13][10];
    ele[10][10] != ele[13][11];
    ele[10][10] != ele[13][12];
    ele[10][10] != ele[13][13];
    ele[10][10] != ele[13][14];
    ele[10][10] != ele[14][10];
    ele[10][10] != ele[14][11];
    ele[10][10] != ele[14][12];
    ele[10][10] != ele[14][13];
    ele[10][10] != ele[14][14];
    ele[10][10] != ele[15][10];
    ele[10][10] != ele[16][10];
    ele[10][10] != ele[17][10];
    ele[10][10] != ele[18][10];
    ele[10][10] != ele[19][10];
    ele[10][10] != ele[20][10];
    ele[10][10] != ele[21][10];
    ele[10][10] != ele[22][10];
    ele[10][10] != ele[23][10];
    ele[10][10] != ele[24][10];
    ele[10][11] != ele[10][12];
    ele[10][11] != ele[10][13];
    ele[10][11] != ele[10][14];
    ele[10][11] != ele[10][15];
    ele[10][11] != ele[10][16];
    ele[10][11] != ele[10][17];
    ele[10][11] != ele[10][18];
    ele[10][11] != ele[10][19];
    ele[10][11] != ele[10][20];
    ele[10][11] != ele[10][21];
    ele[10][11] != ele[10][22];
    ele[10][11] != ele[10][23];
    ele[10][11] != ele[10][24];
    ele[10][11] != ele[11][10];
    ele[10][11] != ele[11][11];
    ele[10][11] != ele[11][12];
    ele[10][11] != ele[11][13];
    ele[10][11] != ele[11][14];
    ele[10][11] != ele[12][10];
    ele[10][11] != ele[12][11];
    ele[10][11] != ele[12][12];
    ele[10][11] != ele[12][13];
    ele[10][11] != ele[12][14];
    ele[10][11] != ele[13][10];
    ele[10][11] != ele[13][11];
    ele[10][11] != ele[13][12];
    ele[10][11] != ele[13][13];
    ele[10][11] != ele[13][14];
    ele[10][11] != ele[14][10];
    ele[10][11] != ele[14][11];
    ele[10][11] != ele[14][12];
    ele[10][11] != ele[14][13];
    ele[10][11] != ele[14][14];
    ele[10][11] != ele[15][11];
    ele[10][11] != ele[16][11];
    ele[10][11] != ele[17][11];
    ele[10][11] != ele[18][11];
    ele[10][11] != ele[19][11];
    ele[10][11] != ele[20][11];
    ele[10][11] != ele[21][11];
    ele[10][11] != ele[22][11];
    ele[10][11] != ele[23][11];
    ele[10][11] != ele[24][11];
    ele[10][12] != ele[10][13];
    ele[10][12] != ele[10][14];
    ele[10][12] != ele[10][15];
    ele[10][12] != ele[10][16];
    ele[10][12] != ele[10][17];
    ele[10][12] != ele[10][18];
    ele[10][12] != ele[10][19];
    ele[10][12] != ele[10][20];
    ele[10][12] != ele[10][21];
    ele[10][12] != ele[10][22];
    ele[10][12] != ele[10][23];
    ele[10][12] != ele[10][24];
    ele[10][12] != ele[11][10];
    ele[10][12] != ele[11][11];
    ele[10][12] != ele[11][12];
    ele[10][12] != ele[11][13];
    ele[10][12] != ele[11][14];
    ele[10][12] != ele[12][10];
    ele[10][12] != ele[12][11];
    ele[10][12] != ele[12][12];
    ele[10][12] != ele[12][13];
    ele[10][12] != ele[12][14];
    ele[10][12] != ele[13][10];
    ele[10][12] != ele[13][11];
    ele[10][12] != ele[13][12];
    ele[10][12] != ele[13][13];
    ele[10][12] != ele[13][14];
    ele[10][12] != ele[14][10];
    ele[10][12] != ele[14][11];
    ele[10][12] != ele[14][12];
    ele[10][12] != ele[14][13];
    ele[10][12] != ele[14][14];
    ele[10][12] != ele[15][12];
    ele[10][12] != ele[16][12];
    ele[10][12] != ele[17][12];
    ele[10][12] != ele[18][12];
    ele[10][12] != ele[19][12];
    ele[10][12] != ele[20][12];
    ele[10][12] != ele[21][12];
    ele[10][12] != ele[22][12];
    ele[10][12] != ele[23][12];
    ele[10][12] != ele[24][12];
    ele[10][13] != ele[10][14];
    ele[10][13] != ele[10][15];
    ele[10][13] != ele[10][16];
    ele[10][13] != ele[10][17];
    ele[10][13] != ele[10][18];
    ele[10][13] != ele[10][19];
    ele[10][13] != ele[10][20];
    ele[10][13] != ele[10][21];
    ele[10][13] != ele[10][22];
    ele[10][13] != ele[10][23];
    ele[10][13] != ele[10][24];
    ele[10][13] != ele[11][10];
    ele[10][13] != ele[11][11];
    ele[10][13] != ele[11][12];
    ele[10][13] != ele[11][13];
    ele[10][13] != ele[11][14];
    ele[10][13] != ele[12][10];
    ele[10][13] != ele[12][11];
    ele[10][13] != ele[12][12];
    ele[10][13] != ele[12][13];
    ele[10][13] != ele[12][14];
    ele[10][13] != ele[13][10];
    ele[10][13] != ele[13][11];
    ele[10][13] != ele[13][12];
    ele[10][13] != ele[13][13];
    ele[10][13] != ele[13][14];
    ele[10][13] != ele[14][10];
    ele[10][13] != ele[14][11];
    ele[10][13] != ele[14][12];
    ele[10][13] != ele[14][13];
    ele[10][13] != ele[14][14];
    ele[10][13] != ele[15][13];
    ele[10][13] != ele[16][13];
    ele[10][13] != ele[17][13];
    ele[10][13] != ele[18][13];
    ele[10][13] != ele[19][13];
    ele[10][13] != ele[20][13];
    ele[10][13] != ele[21][13];
    ele[10][13] != ele[22][13];
    ele[10][13] != ele[23][13];
    ele[10][13] != ele[24][13];
    ele[10][14] != ele[10][15];
    ele[10][14] != ele[10][16];
    ele[10][14] != ele[10][17];
    ele[10][14] != ele[10][18];
    ele[10][14] != ele[10][19];
    ele[10][14] != ele[10][20];
    ele[10][14] != ele[10][21];
    ele[10][14] != ele[10][22];
    ele[10][14] != ele[10][23];
    ele[10][14] != ele[10][24];
    ele[10][14] != ele[11][10];
    ele[10][14] != ele[11][11];
    ele[10][14] != ele[11][12];
    ele[10][14] != ele[11][13];
    ele[10][14] != ele[11][14];
    ele[10][14] != ele[12][10];
    ele[10][14] != ele[12][11];
    ele[10][14] != ele[12][12];
    ele[10][14] != ele[12][13];
    ele[10][14] != ele[12][14];
    ele[10][14] != ele[13][10];
    ele[10][14] != ele[13][11];
    ele[10][14] != ele[13][12];
    ele[10][14] != ele[13][13];
    ele[10][14] != ele[13][14];
    ele[10][14] != ele[14][10];
    ele[10][14] != ele[14][11];
    ele[10][14] != ele[14][12];
    ele[10][14] != ele[14][13];
    ele[10][14] != ele[14][14];
    ele[10][14] != ele[15][14];
    ele[10][14] != ele[16][14];
    ele[10][14] != ele[17][14];
    ele[10][14] != ele[18][14];
    ele[10][14] != ele[19][14];
    ele[10][14] != ele[20][14];
    ele[10][14] != ele[21][14];
    ele[10][14] != ele[22][14];
    ele[10][14] != ele[23][14];
    ele[10][14] != ele[24][14];
    ele[10][15] != ele[10][16];
    ele[10][15] != ele[10][17];
    ele[10][15] != ele[10][18];
    ele[10][15] != ele[10][19];
    ele[10][15] != ele[10][20];
    ele[10][15] != ele[10][21];
    ele[10][15] != ele[10][22];
    ele[10][15] != ele[10][23];
    ele[10][15] != ele[10][24];
    ele[10][15] != ele[11][15];
    ele[10][15] != ele[11][16];
    ele[10][15] != ele[11][17];
    ele[10][15] != ele[11][18];
    ele[10][15] != ele[11][19];
    ele[10][15] != ele[12][15];
    ele[10][15] != ele[12][16];
    ele[10][15] != ele[12][17];
    ele[10][15] != ele[12][18];
    ele[10][15] != ele[12][19];
    ele[10][15] != ele[13][15];
    ele[10][15] != ele[13][16];
    ele[10][15] != ele[13][17];
    ele[10][15] != ele[13][18];
    ele[10][15] != ele[13][19];
    ele[10][15] != ele[14][15];
    ele[10][15] != ele[14][16];
    ele[10][15] != ele[14][17];
    ele[10][15] != ele[14][18];
    ele[10][15] != ele[14][19];
    ele[10][15] != ele[15][15];
    ele[10][15] != ele[16][15];
    ele[10][15] != ele[17][15];
    ele[10][15] != ele[18][15];
    ele[10][15] != ele[19][15];
    ele[10][15] != ele[20][15];
    ele[10][15] != ele[21][15];
    ele[10][15] != ele[22][15];
    ele[10][15] != ele[23][15];
    ele[10][15] != ele[24][15];
    ele[10][16] != ele[10][17];
    ele[10][16] != ele[10][18];
    ele[10][16] != ele[10][19];
    ele[10][16] != ele[10][20];
    ele[10][16] != ele[10][21];
    ele[10][16] != ele[10][22];
    ele[10][16] != ele[10][23];
    ele[10][16] != ele[10][24];
    ele[10][16] != ele[11][15];
    ele[10][16] != ele[11][16];
    ele[10][16] != ele[11][17];
    ele[10][16] != ele[11][18];
    ele[10][16] != ele[11][19];
    ele[10][16] != ele[12][15];
    ele[10][16] != ele[12][16];
    ele[10][16] != ele[12][17];
    ele[10][16] != ele[12][18];
    ele[10][16] != ele[12][19];
    ele[10][16] != ele[13][15];
    ele[10][16] != ele[13][16];
    ele[10][16] != ele[13][17];
    ele[10][16] != ele[13][18];
    ele[10][16] != ele[13][19];
    ele[10][16] != ele[14][15];
    ele[10][16] != ele[14][16];
    ele[10][16] != ele[14][17];
    ele[10][16] != ele[14][18];
    ele[10][16] != ele[14][19];
    ele[10][16] != ele[15][16];
    ele[10][16] != ele[16][16];
    ele[10][16] != ele[17][16];
    ele[10][16] != ele[18][16];
    ele[10][16] != ele[19][16];
    ele[10][16] != ele[20][16];
    ele[10][16] != ele[21][16];
    ele[10][16] != ele[22][16];
    ele[10][16] != ele[23][16];
    ele[10][16] != ele[24][16];
    ele[10][17] != ele[10][18];
    ele[10][17] != ele[10][19];
    ele[10][17] != ele[10][20];
    ele[10][17] != ele[10][21];
    ele[10][17] != ele[10][22];
    ele[10][17] != ele[10][23];
    ele[10][17] != ele[10][24];
    ele[10][17] != ele[11][15];
    ele[10][17] != ele[11][16];
    ele[10][17] != ele[11][17];
    ele[10][17] != ele[11][18];
    ele[10][17] != ele[11][19];
    ele[10][17] != ele[12][15];
    ele[10][17] != ele[12][16];
    ele[10][17] != ele[12][17];
    ele[10][17] != ele[12][18];
    ele[10][17] != ele[12][19];
    ele[10][17] != ele[13][15];
    ele[10][17] != ele[13][16];
    ele[10][17] != ele[13][17];
    ele[10][17] != ele[13][18];
    ele[10][17] != ele[13][19];
    ele[10][17] != ele[14][15];
    ele[10][17] != ele[14][16];
    ele[10][17] != ele[14][17];
    ele[10][17] != ele[14][18];
    ele[10][17] != ele[14][19];
    ele[10][17] != ele[15][17];
    ele[10][17] != ele[16][17];
    ele[10][17] != ele[17][17];
    ele[10][17] != ele[18][17];
    ele[10][17] != ele[19][17];
    ele[10][17] != ele[20][17];
    ele[10][17] != ele[21][17];
    ele[10][17] != ele[22][17];
    ele[10][17] != ele[23][17];
    ele[10][17] != ele[24][17];
    ele[10][18] != ele[10][19];
    ele[10][18] != ele[10][20];
    ele[10][18] != ele[10][21];
    ele[10][18] != ele[10][22];
    ele[10][18] != ele[10][23];
    ele[10][18] != ele[10][24];
    ele[10][18] != ele[11][15];
    ele[10][18] != ele[11][16];
    ele[10][18] != ele[11][17];
    ele[10][18] != ele[11][18];
    ele[10][18] != ele[11][19];
    ele[10][18] != ele[12][15];
    ele[10][18] != ele[12][16];
    ele[10][18] != ele[12][17];
    ele[10][18] != ele[12][18];
    ele[10][18] != ele[12][19];
    ele[10][18] != ele[13][15];
    ele[10][18] != ele[13][16];
    ele[10][18] != ele[13][17];
    ele[10][18] != ele[13][18];
    ele[10][18] != ele[13][19];
    ele[10][18] != ele[14][15];
    ele[10][18] != ele[14][16];
    ele[10][18] != ele[14][17];
    ele[10][18] != ele[14][18];
    ele[10][18] != ele[14][19];
    ele[10][18] != ele[15][18];
    ele[10][18] != ele[16][18];
    ele[10][18] != ele[17][18];
    ele[10][18] != ele[18][18];
    ele[10][18] != ele[19][18];
    ele[10][18] != ele[20][18];
    ele[10][18] != ele[21][18];
    ele[10][18] != ele[22][18];
    ele[10][18] != ele[23][18];
    ele[10][18] != ele[24][18];
    ele[10][19] != ele[10][20];
    ele[10][19] != ele[10][21];
    ele[10][19] != ele[10][22];
    ele[10][19] != ele[10][23];
    ele[10][19] != ele[10][24];
    ele[10][19] != ele[11][15];
    ele[10][19] != ele[11][16];
    ele[10][19] != ele[11][17];
    ele[10][19] != ele[11][18];
    ele[10][19] != ele[11][19];
    ele[10][19] != ele[12][15];
    ele[10][19] != ele[12][16];
    ele[10][19] != ele[12][17];
    ele[10][19] != ele[12][18];
    ele[10][19] != ele[12][19];
    ele[10][19] != ele[13][15];
    ele[10][19] != ele[13][16];
    ele[10][19] != ele[13][17];
    ele[10][19] != ele[13][18];
    ele[10][19] != ele[13][19];
    ele[10][19] != ele[14][15];
    ele[10][19] != ele[14][16];
    ele[10][19] != ele[14][17];
    ele[10][19] != ele[14][18];
    ele[10][19] != ele[14][19];
    ele[10][19] != ele[15][19];
    ele[10][19] != ele[16][19];
    ele[10][19] != ele[17][19];
    ele[10][19] != ele[18][19];
    ele[10][19] != ele[19][19];
    ele[10][19] != ele[20][19];
    ele[10][19] != ele[21][19];
    ele[10][19] != ele[22][19];
    ele[10][19] != ele[23][19];
    ele[10][19] != ele[24][19];
    ele[10][2] != ele[10][10];
    ele[10][2] != ele[10][11];
    ele[10][2] != ele[10][12];
    ele[10][2] != ele[10][13];
    ele[10][2] != ele[10][14];
    ele[10][2] != ele[10][15];
    ele[10][2] != ele[10][16];
    ele[10][2] != ele[10][17];
    ele[10][2] != ele[10][18];
    ele[10][2] != ele[10][19];
    ele[10][2] != ele[10][20];
    ele[10][2] != ele[10][21];
    ele[10][2] != ele[10][22];
    ele[10][2] != ele[10][23];
    ele[10][2] != ele[10][24];
    ele[10][2] != ele[10][3];
    ele[10][2] != ele[10][4];
    ele[10][2] != ele[10][5];
    ele[10][2] != ele[10][6];
    ele[10][2] != ele[10][7];
    ele[10][2] != ele[10][8];
    ele[10][2] != ele[10][9];
    ele[10][2] != ele[11][0];
    ele[10][2] != ele[11][1];
    ele[10][2] != ele[11][2];
    ele[10][2] != ele[11][3];
    ele[10][2] != ele[11][4];
    ele[10][2] != ele[12][0];
    ele[10][2] != ele[12][1];
    ele[10][2] != ele[12][2];
    ele[10][2] != ele[12][3];
    ele[10][2] != ele[12][4];
    ele[10][2] != ele[13][0];
    ele[10][2] != ele[13][1];
    ele[10][2] != ele[13][2];
    ele[10][2] != ele[13][3];
    ele[10][2] != ele[13][4];
    ele[10][2] != ele[14][0];
    ele[10][2] != ele[14][1];
    ele[10][2] != ele[14][2];
    ele[10][2] != ele[14][3];
    ele[10][2] != ele[14][4];
    ele[10][2] != ele[15][2];
    ele[10][2] != ele[16][2];
    ele[10][2] != ele[17][2];
    ele[10][2] != ele[18][2];
    ele[10][2] != ele[19][2];
    ele[10][2] != ele[20][2];
    ele[10][2] != ele[21][2];
    ele[10][2] != ele[22][2];
    ele[10][2] != ele[23][2];
    ele[10][2] != ele[24][2];
    ele[10][20] != ele[10][21];
    ele[10][20] != ele[10][22];
    ele[10][20] != ele[10][23];
    ele[10][20] != ele[10][24];
    ele[10][20] != ele[11][20];
    ele[10][20] != ele[11][21];
    ele[10][20] != ele[11][22];
    ele[10][20] != ele[11][23];
    ele[10][20] != ele[11][24];
    ele[10][20] != ele[12][20];
    ele[10][20] != ele[12][21];
    ele[10][20] != ele[12][22];
    ele[10][20] != ele[12][23];
    ele[10][20] != ele[12][24];
    ele[10][20] != ele[13][20];
    ele[10][20] != ele[13][21];
    ele[10][20] != ele[13][22];
    ele[10][20] != ele[13][23];
    ele[10][20] != ele[13][24];
    ele[10][20] != ele[14][20];
    ele[10][20] != ele[14][21];
    ele[10][20] != ele[14][22];
    ele[10][20] != ele[14][23];
    ele[10][20] != ele[14][24];
    ele[10][20] != ele[15][20];
    ele[10][20] != ele[16][20];
    ele[10][20] != ele[17][20];
    ele[10][20] != ele[18][20];
    ele[10][20] != ele[19][20];
    ele[10][20] != ele[20][20];
    ele[10][20] != ele[21][20];
    ele[10][20] != ele[22][20];
    ele[10][20] != ele[23][20];
    ele[10][20] != ele[24][20];
    ele[10][21] != ele[10][22];
    ele[10][21] != ele[10][23];
    ele[10][21] != ele[10][24];
    ele[10][21] != ele[11][20];
    ele[10][21] != ele[11][21];
    ele[10][21] != ele[11][22];
    ele[10][21] != ele[11][23];
    ele[10][21] != ele[11][24];
    ele[10][21] != ele[12][20];
    ele[10][21] != ele[12][21];
    ele[10][21] != ele[12][22];
    ele[10][21] != ele[12][23];
    ele[10][21] != ele[12][24];
    ele[10][21] != ele[13][20];
    ele[10][21] != ele[13][21];
    ele[10][21] != ele[13][22];
    ele[10][21] != ele[13][23];
    ele[10][21] != ele[13][24];
    ele[10][21] != ele[14][20];
    ele[10][21] != ele[14][21];
    ele[10][21] != ele[14][22];
    ele[10][21] != ele[14][23];
    ele[10][21] != ele[14][24];
    ele[10][21] != ele[15][21];
    ele[10][21] != ele[16][21];
    ele[10][21] != ele[17][21];
    ele[10][21] != ele[18][21];
    ele[10][21] != ele[19][21];
    ele[10][21] != ele[20][21];
    ele[10][21] != ele[21][21];
    ele[10][21] != ele[22][21];
    ele[10][21] != ele[23][21];
    ele[10][21] != ele[24][21];
    ele[10][22] != ele[10][23];
    ele[10][22] != ele[10][24];
    ele[10][22] != ele[11][20];
    ele[10][22] != ele[11][21];
    ele[10][22] != ele[11][22];
    ele[10][22] != ele[11][23];
    ele[10][22] != ele[11][24];
    ele[10][22] != ele[12][20];
    ele[10][22] != ele[12][21];
    ele[10][22] != ele[12][22];
    ele[10][22] != ele[12][23];
    ele[10][22] != ele[12][24];
    ele[10][22] != ele[13][20];
    ele[10][22] != ele[13][21];
    ele[10][22] != ele[13][22];
    ele[10][22] != ele[13][23];
    ele[10][22] != ele[13][24];
    ele[10][22] != ele[14][20];
    ele[10][22] != ele[14][21];
    ele[10][22] != ele[14][22];
    ele[10][22] != ele[14][23];
    ele[10][22] != ele[14][24];
    ele[10][22] != ele[15][22];
    ele[10][22] != ele[16][22];
    ele[10][22] != ele[17][22];
    ele[10][22] != ele[18][22];
    ele[10][22] != ele[19][22];
    ele[10][22] != ele[20][22];
    ele[10][22] != ele[21][22];
    ele[10][22] != ele[22][22];
    ele[10][22] != ele[23][22];
    ele[10][22] != ele[24][22];
    ele[10][23] != ele[10][24];
    ele[10][23] != ele[11][20];
    ele[10][23] != ele[11][21];
    ele[10][23] != ele[11][22];
    ele[10][23] != ele[11][23];
    ele[10][23] != ele[11][24];
    ele[10][23] != ele[12][20];
    ele[10][23] != ele[12][21];
    ele[10][23] != ele[12][22];
    ele[10][23] != ele[12][23];
    ele[10][23] != ele[12][24];
    ele[10][23] != ele[13][20];
    ele[10][23] != ele[13][21];
    ele[10][23] != ele[13][22];
    ele[10][23] != ele[13][23];
    ele[10][23] != ele[13][24];
    ele[10][23] != ele[14][20];
    ele[10][23] != ele[14][21];
    ele[10][23] != ele[14][22];
    ele[10][23] != ele[14][23];
    ele[10][23] != ele[14][24];
    ele[10][23] != ele[15][23];
    ele[10][23] != ele[16][23];
    ele[10][23] != ele[17][23];
    ele[10][23] != ele[18][23];
    ele[10][23] != ele[19][23];
    ele[10][23] != ele[20][23];
    ele[10][23] != ele[21][23];
    ele[10][23] != ele[22][23];
    ele[10][23] != ele[23][23];
    ele[10][23] != ele[24][23];
    ele[10][24] != ele[11][20];
    ele[10][24] != ele[11][21];
    ele[10][24] != ele[11][22];
    ele[10][24] != ele[11][23];
    ele[10][24] != ele[11][24];
    ele[10][24] != ele[12][20];
    ele[10][24] != ele[12][21];
    ele[10][24] != ele[12][22];
    ele[10][24] != ele[12][23];
    ele[10][24] != ele[12][24];
    ele[10][24] != ele[13][20];
    ele[10][24] != ele[13][21];
    ele[10][24] != ele[13][22];
    ele[10][24] != ele[13][23];
    ele[10][24] != ele[13][24];
    ele[10][24] != ele[14][20];
    ele[10][24] != ele[14][21];
    ele[10][24] != ele[14][22];
    ele[10][24] != ele[14][23];
    ele[10][24] != ele[14][24];
    ele[10][24] != ele[15][24];
    ele[10][24] != ele[16][24];
    ele[10][24] != ele[17][24];
    ele[10][24] != ele[18][24];
    ele[10][24] != ele[19][24];
    ele[10][24] != ele[20][24];
    ele[10][24] != ele[21][24];
    ele[10][24] != ele[22][24];
    ele[10][24] != ele[23][24];
    ele[10][24] != ele[24][24];
    ele[10][3] != ele[10][10];
    ele[10][3] != ele[10][11];
    ele[10][3] != ele[10][12];
    ele[10][3] != ele[10][13];
    ele[10][3] != ele[10][14];
    ele[10][3] != ele[10][15];
    ele[10][3] != ele[10][16];
    ele[10][3] != ele[10][17];
    ele[10][3] != ele[10][18];
    ele[10][3] != ele[10][19];
    ele[10][3] != ele[10][20];
    ele[10][3] != ele[10][21];
    ele[10][3] != ele[10][22];
    ele[10][3] != ele[10][23];
    ele[10][3] != ele[10][24];
    ele[10][3] != ele[10][4];
    ele[10][3] != ele[10][5];
    ele[10][3] != ele[10][6];
    ele[10][3] != ele[10][7];
    ele[10][3] != ele[10][8];
    ele[10][3] != ele[10][9];
    ele[10][3] != ele[11][0];
    ele[10][3] != ele[11][1];
    ele[10][3] != ele[11][2];
    ele[10][3] != ele[11][3];
    ele[10][3] != ele[11][4];
    ele[10][3] != ele[12][0];
    ele[10][3] != ele[12][1];
    ele[10][3] != ele[12][2];
    ele[10][3] != ele[12][3];
    ele[10][3] != ele[12][4];
    ele[10][3] != ele[13][0];
    ele[10][3] != ele[13][1];
    ele[10][3] != ele[13][2];
    ele[10][3] != ele[13][3];
    ele[10][3] != ele[13][4];
    ele[10][3] != ele[14][0];
    ele[10][3] != ele[14][1];
    ele[10][3] != ele[14][2];
    ele[10][3] != ele[14][3];
    ele[10][3] != ele[14][4];
    ele[10][3] != ele[15][3];
    ele[10][3] != ele[16][3];
    ele[10][3] != ele[17][3];
    ele[10][3] != ele[18][3];
    ele[10][3] != ele[19][3];
    ele[10][3] != ele[20][3];
    ele[10][3] != ele[21][3];
    ele[10][3] != ele[22][3];
    ele[10][3] != ele[23][3];
    ele[10][3] != ele[24][3];
    ele[10][4] != ele[10][10];
    ele[10][4] != ele[10][11];
    ele[10][4] != ele[10][12];
    ele[10][4] != ele[10][13];
    ele[10][4] != ele[10][14];
    ele[10][4] != ele[10][15];
    ele[10][4] != ele[10][16];
    ele[10][4] != ele[10][17];
    ele[10][4] != ele[10][18];
    ele[10][4] != ele[10][19];
    ele[10][4] != ele[10][20];
    ele[10][4] != ele[10][21];
    ele[10][4] != ele[10][22];
    ele[10][4] != ele[10][23];
    ele[10][4] != ele[10][24];
    ele[10][4] != ele[10][5];
    ele[10][4] != ele[10][6];
    ele[10][4] != ele[10][7];
    ele[10][4] != ele[10][8];
    ele[10][4] != ele[10][9];
    ele[10][4] != ele[11][0];
    ele[10][4] != ele[11][1];
    ele[10][4] != ele[11][2];
    ele[10][4] != ele[11][3];
    ele[10][4] != ele[11][4];
    ele[10][4] != ele[12][0];
    ele[10][4] != ele[12][1];
    ele[10][4] != ele[12][2];
    ele[10][4] != ele[12][3];
    ele[10][4] != ele[12][4];
    ele[10][4] != ele[13][0];
    ele[10][4] != ele[13][1];
    ele[10][4] != ele[13][2];
    ele[10][4] != ele[13][3];
    ele[10][4] != ele[13][4];
    ele[10][4] != ele[14][0];
    ele[10][4] != ele[14][1];
    ele[10][4] != ele[14][2];
    ele[10][4] != ele[14][3];
    ele[10][4] != ele[14][4];
    ele[10][4] != ele[15][4];
    ele[10][4] != ele[16][4];
    ele[10][4] != ele[17][4];
    ele[10][4] != ele[18][4];
    ele[10][4] != ele[19][4];
    ele[10][4] != ele[20][4];
    ele[10][4] != ele[21][4];
    ele[10][4] != ele[22][4];
    ele[10][4] != ele[23][4];
    ele[10][4] != ele[24][4];
    ele[10][5] != ele[10][10];
    ele[10][5] != ele[10][11];
    ele[10][5] != ele[10][12];
    ele[10][5] != ele[10][13];
    ele[10][5] != ele[10][14];
    ele[10][5] != ele[10][15];
    ele[10][5] != ele[10][16];
    ele[10][5] != ele[10][17];
    ele[10][5] != ele[10][18];
    ele[10][5] != ele[10][19];
    ele[10][5] != ele[10][20];
    ele[10][5] != ele[10][21];
    ele[10][5] != ele[10][22];
    ele[10][5] != ele[10][23];
    ele[10][5] != ele[10][24];
    ele[10][5] != ele[10][6];
    ele[10][5] != ele[10][7];
    ele[10][5] != ele[10][8];
    ele[10][5] != ele[10][9];
    ele[10][5] != ele[11][5];
    ele[10][5] != ele[11][6];
    ele[10][5] != ele[11][7];
    ele[10][5] != ele[11][8];
    ele[10][5] != ele[11][9];
    ele[10][5] != ele[12][5];
    ele[10][5] != ele[12][6];
    ele[10][5] != ele[12][7];
    ele[10][5] != ele[12][8];
    ele[10][5] != ele[12][9];
    ele[10][5] != ele[13][5];
    ele[10][5] != ele[13][6];
    ele[10][5] != ele[13][7];
    ele[10][5] != ele[13][8];
    ele[10][5] != ele[13][9];
    ele[10][5] != ele[14][5];
    ele[10][5] != ele[14][6];
    ele[10][5] != ele[14][7];
    ele[10][5] != ele[14][8];
    ele[10][5] != ele[14][9];
    ele[10][5] != ele[15][5];
    ele[10][5] != ele[16][5];
    ele[10][5] != ele[17][5];
    ele[10][5] != ele[18][5];
    ele[10][5] != ele[19][5];
    ele[10][5] != ele[20][5];
    ele[10][5] != ele[21][5];
    ele[10][5] != ele[22][5];
    ele[10][5] != ele[23][5];
    ele[10][5] != ele[24][5];
    ele[10][6] != ele[10][10];
    ele[10][6] != ele[10][11];
    ele[10][6] != ele[10][12];
    ele[10][6] != ele[10][13];
    ele[10][6] != ele[10][14];
    ele[10][6] != ele[10][15];
    ele[10][6] != ele[10][16];
    ele[10][6] != ele[10][17];
    ele[10][6] != ele[10][18];
    ele[10][6] != ele[10][19];
    ele[10][6] != ele[10][20];
    ele[10][6] != ele[10][21];
    ele[10][6] != ele[10][22];
    ele[10][6] != ele[10][23];
    ele[10][6] != ele[10][24];
    ele[10][6] != ele[10][7];
    ele[10][6] != ele[10][8];
    ele[10][6] != ele[10][9];
    ele[10][6] != ele[11][5];
    ele[10][6] != ele[11][6];
    ele[10][6] != ele[11][7];
    ele[10][6] != ele[11][8];
    ele[10][6] != ele[11][9];
    ele[10][6] != ele[12][5];
    ele[10][6] != ele[12][6];
    ele[10][6] != ele[12][7];
    ele[10][6] != ele[12][8];
    ele[10][6] != ele[12][9];
    ele[10][6] != ele[13][5];
    ele[10][6] != ele[13][6];
    ele[10][6] != ele[13][7];
    ele[10][6] != ele[13][8];
    ele[10][6] != ele[13][9];
    ele[10][6] != ele[14][5];
    ele[10][6] != ele[14][6];
    ele[10][6] != ele[14][7];
    ele[10][6] != ele[14][8];
    ele[10][6] != ele[14][9];
    ele[10][6] != ele[15][6];
    ele[10][6] != ele[16][6];
    ele[10][6] != ele[17][6];
    ele[10][6] != ele[18][6];
    ele[10][6] != ele[19][6];
    ele[10][6] != ele[20][6];
    ele[10][6] != ele[21][6];
    ele[10][6] != ele[22][6];
    ele[10][6] != ele[23][6];
    ele[10][6] != ele[24][6];
    ele[10][7] != ele[10][10];
    ele[10][7] != ele[10][11];
    ele[10][7] != ele[10][12];
    ele[10][7] != ele[10][13];
    ele[10][7] != ele[10][14];
    ele[10][7] != ele[10][15];
    ele[10][7] != ele[10][16];
    ele[10][7] != ele[10][17];
    ele[10][7] != ele[10][18];
    ele[10][7] != ele[10][19];
    ele[10][7] != ele[10][20];
    ele[10][7] != ele[10][21];
    ele[10][7] != ele[10][22];
    ele[10][7] != ele[10][23];
    ele[10][7] != ele[10][24];
    ele[10][7] != ele[10][8];
    ele[10][7] != ele[10][9];
    ele[10][7] != ele[11][5];
    ele[10][7] != ele[11][6];
    ele[10][7] != ele[11][7];
    ele[10][7] != ele[11][8];
    ele[10][7] != ele[11][9];
    ele[10][7] != ele[12][5];
    ele[10][7] != ele[12][6];
    ele[10][7] != ele[12][7];
    ele[10][7] != ele[12][8];
    ele[10][7] != ele[12][9];
    ele[10][7] != ele[13][5];
    ele[10][7] != ele[13][6];
    ele[10][7] != ele[13][7];
    ele[10][7] != ele[13][8];
    ele[10][7] != ele[13][9];
    ele[10][7] != ele[14][5];
    ele[10][7] != ele[14][6];
    ele[10][7] != ele[14][7];
    ele[10][7] != ele[14][8];
    ele[10][7] != ele[14][9];
    ele[10][7] != ele[15][7];
    ele[10][7] != ele[16][7];
    ele[10][7] != ele[17][7];
    ele[10][7] != ele[18][7];
    ele[10][7] != ele[19][7];
    ele[10][7] != ele[20][7];
    ele[10][7] != ele[21][7];
    ele[10][7] != ele[22][7];
    ele[10][7] != ele[23][7];
    ele[10][7] != ele[24][7];
    ele[10][8] != ele[10][10];
    ele[10][8] != ele[10][11];
    ele[10][8] != ele[10][12];
    ele[10][8] != ele[10][13];
    ele[10][8] != ele[10][14];
    ele[10][8] != ele[10][15];
    ele[10][8] != ele[10][16];
    ele[10][8] != ele[10][17];
    ele[10][8] != ele[10][18];
    ele[10][8] != ele[10][19];
    ele[10][8] != ele[10][20];
    ele[10][8] != ele[10][21];
    ele[10][8] != ele[10][22];
    ele[10][8] != ele[10][23];
    ele[10][8] != ele[10][24];
    ele[10][8] != ele[10][9];
    ele[10][8] != ele[11][5];
    ele[10][8] != ele[11][6];
    ele[10][8] != ele[11][7];
    ele[10][8] != ele[11][8];
    ele[10][8] != ele[11][9];
    ele[10][8] != ele[12][5];
    ele[10][8] != ele[12][6];
    ele[10][8] != ele[12][7];
    ele[10][8] != ele[12][8];
    ele[10][8] != ele[12][9];
    ele[10][8] != ele[13][5];
    ele[10][8] != ele[13][6];
    ele[10][8] != ele[13][7];
    ele[10][8] != ele[13][8];
    ele[10][8] != ele[13][9];
    ele[10][8] != ele[14][5];
    ele[10][8] != ele[14][6];
    ele[10][8] != ele[14][7];
    ele[10][8] != ele[14][8];
    ele[10][8] != ele[14][9];
    ele[10][8] != ele[15][8];
    ele[10][8] != ele[16][8];
    ele[10][8] != ele[17][8];
    ele[10][8] != ele[18][8];
    ele[10][8] != ele[19][8];
    ele[10][8] != ele[20][8];
    ele[10][8] != ele[21][8];
    ele[10][8] != ele[22][8];
    ele[10][8] != ele[23][8];
    ele[10][8] != ele[24][8];
    ele[10][9] != ele[10][10];
    ele[10][9] != ele[10][11];
    ele[10][9] != ele[10][12];
    ele[10][9] != ele[10][13];
    ele[10][9] != ele[10][14];
    ele[10][9] != ele[10][15];
    ele[10][9] != ele[10][16];
    ele[10][9] != ele[10][17];
    ele[10][9] != ele[10][18];
    ele[10][9] != ele[10][19];
    ele[10][9] != ele[10][20];
    ele[10][9] != ele[10][21];
    ele[10][9] != ele[10][22];
    ele[10][9] != ele[10][23];
    ele[10][9] != ele[10][24];
    ele[10][9] != ele[11][5];
    ele[10][9] != ele[11][6];
    ele[10][9] != ele[11][7];
    ele[10][9] != ele[11][8];
    ele[10][9] != ele[11][9];
    ele[10][9] != ele[12][5];
    ele[10][9] != ele[12][6];
    ele[10][9] != ele[12][7];
    ele[10][9] != ele[12][8];
    ele[10][9] != ele[12][9];
    ele[10][9] != ele[13][5];
    ele[10][9] != ele[13][6];
    ele[10][9] != ele[13][7];
    ele[10][9] != ele[13][8];
    ele[10][9] != ele[13][9];
    ele[10][9] != ele[14][5];
    ele[10][9] != ele[14][6];
    ele[10][9] != ele[14][7];
    ele[10][9] != ele[14][8];
    ele[10][9] != ele[14][9];
    ele[10][9] != ele[15][9];
    ele[10][9] != ele[16][9];
    ele[10][9] != ele[17][9];
    ele[10][9] != ele[18][9];
    ele[10][9] != ele[19][9];
    ele[10][9] != ele[20][9];
    ele[10][9] != ele[21][9];
    ele[10][9] != ele[22][9];
    ele[10][9] != ele[23][9];
    ele[10][9] != ele[24][9];
    ele[11][0] != ele[11][1];
    ele[11][0] != ele[11][10];
    ele[11][0] != ele[11][11];
    ele[11][0] != ele[11][12];
    ele[11][0] != ele[11][13];
    ele[11][0] != ele[11][14];
    ele[11][0] != ele[11][15];
    ele[11][0] != ele[11][16];
    ele[11][0] != ele[11][17];
    ele[11][0] != ele[11][18];
    ele[11][0] != ele[11][19];
    ele[11][0] != ele[11][2];
    ele[11][0] != ele[11][20];
    ele[11][0] != ele[11][21];
    ele[11][0] != ele[11][22];
    ele[11][0] != ele[11][23];
    ele[11][0] != ele[11][24];
    ele[11][0] != ele[11][3];
    ele[11][0] != ele[11][4];
    ele[11][0] != ele[11][5];
    ele[11][0] != ele[11][6];
    ele[11][0] != ele[11][7];
    ele[11][0] != ele[11][8];
    ele[11][0] != ele[11][9];
    ele[11][0] != ele[12][0];
    ele[11][0] != ele[12][1];
    ele[11][0] != ele[12][2];
    ele[11][0] != ele[12][3];
    ele[11][0] != ele[12][4];
    ele[11][0] != ele[13][0];
    ele[11][0] != ele[13][1];
    ele[11][0] != ele[13][2];
    ele[11][0] != ele[13][3];
    ele[11][0] != ele[13][4];
    ele[11][0] != ele[14][0];
    ele[11][0] != ele[14][1];
    ele[11][0] != ele[14][2];
    ele[11][0] != ele[14][3];
    ele[11][0] != ele[14][4];
    ele[11][0] != ele[15][0];
    ele[11][0] != ele[16][0];
    ele[11][0] != ele[17][0];
    ele[11][0] != ele[18][0];
    ele[11][0] != ele[19][0];
    ele[11][0] != ele[20][0];
    ele[11][0] != ele[21][0];
    ele[11][0] != ele[22][0];
    ele[11][0] != ele[23][0];
    ele[11][0] != ele[24][0];
    ele[11][1] != ele[11][10];
    ele[11][1] != ele[11][11];
    ele[11][1] != ele[11][12];
    ele[11][1] != ele[11][13];
    ele[11][1] != ele[11][14];
    ele[11][1] != ele[11][15];
    ele[11][1] != ele[11][16];
    ele[11][1] != ele[11][17];
    ele[11][1] != ele[11][18];
    ele[11][1] != ele[11][19];
    ele[11][1] != ele[11][2];
    ele[11][1] != ele[11][20];
    ele[11][1] != ele[11][21];
    ele[11][1] != ele[11][22];
    ele[11][1] != ele[11][23];
    ele[11][1] != ele[11][24];
    ele[11][1] != ele[11][3];
    ele[11][1] != ele[11][4];
    ele[11][1] != ele[11][5];
    ele[11][1] != ele[11][6];
    ele[11][1] != ele[11][7];
    ele[11][1] != ele[11][8];
    ele[11][1] != ele[11][9];
    ele[11][1] != ele[12][0];
    ele[11][1] != ele[12][1];
    ele[11][1] != ele[12][2];
    ele[11][1] != ele[12][3];
    ele[11][1] != ele[12][4];
    ele[11][1] != ele[13][0];
    ele[11][1] != ele[13][1];
    ele[11][1] != ele[13][2];
    ele[11][1] != ele[13][3];
    ele[11][1] != ele[13][4];
    ele[11][1] != ele[14][0];
    ele[11][1] != ele[14][1];
    ele[11][1] != ele[14][2];
    ele[11][1] != ele[14][3];
    ele[11][1] != ele[14][4];
    ele[11][1] != ele[15][1];
    ele[11][1] != ele[16][1];
    ele[11][1] != ele[17][1];
    ele[11][1] != ele[18][1];
    ele[11][1] != ele[19][1];
    ele[11][1] != ele[20][1];
    ele[11][1] != ele[21][1];
    ele[11][1] != ele[22][1];
    ele[11][1] != ele[23][1];
    ele[11][1] != ele[24][1];
    ele[11][10] != ele[11][11];
    ele[11][10] != ele[11][12];
    ele[11][10] != ele[11][13];
    ele[11][10] != ele[11][14];
    ele[11][10] != ele[11][15];
    ele[11][10] != ele[11][16];
    ele[11][10] != ele[11][17];
    ele[11][10] != ele[11][18];
    ele[11][10] != ele[11][19];
    ele[11][10] != ele[11][20];
    ele[11][10] != ele[11][21];
    ele[11][10] != ele[11][22];
    ele[11][10] != ele[11][23];
    ele[11][10] != ele[11][24];
    ele[11][10] != ele[12][10];
    ele[11][10] != ele[12][11];
    ele[11][10] != ele[12][12];
    ele[11][10] != ele[12][13];
    ele[11][10] != ele[12][14];
    ele[11][10] != ele[13][10];
    ele[11][10] != ele[13][11];
    ele[11][10] != ele[13][12];
    ele[11][10] != ele[13][13];
    ele[11][10] != ele[13][14];
    ele[11][10] != ele[14][10];
    ele[11][10] != ele[14][11];
    ele[11][10] != ele[14][12];
    ele[11][10] != ele[14][13];
    ele[11][10] != ele[14][14];
    ele[11][10] != ele[15][10];
    ele[11][10] != ele[16][10];
    ele[11][10] != ele[17][10];
    ele[11][10] != ele[18][10];
    ele[11][10] != ele[19][10];
    ele[11][10] != ele[20][10];
    ele[11][10] != ele[21][10];
    ele[11][10] != ele[22][10];
    ele[11][10] != ele[23][10];
    ele[11][10] != ele[24][10];
    ele[11][11] != ele[11][12];
    ele[11][11] != ele[11][13];
    ele[11][11] != ele[11][14];
    ele[11][11] != ele[11][15];
    ele[11][11] != ele[11][16];
    ele[11][11] != ele[11][17];
    ele[11][11] != ele[11][18];
    ele[11][11] != ele[11][19];
    ele[11][11] != ele[11][20];
    ele[11][11] != ele[11][21];
    ele[11][11] != ele[11][22];
    ele[11][11] != ele[11][23];
    ele[11][11] != ele[11][24];
    ele[11][11] != ele[12][10];
    ele[11][11] != ele[12][11];
    ele[11][11] != ele[12][12];
    ele[11][11] != ele[12][13];
    ele[11][11] != ele[12][14];
    ele[11][11] != ele[13][10];
    ele[11][11] != ele[13][11];
    ele[11][11] != ele[13][12];
    ele[11][11] != ele[13][13];
    ele[11][11] != ele[13][14];
    ele[11][11] != ele[14][10];
    ele[11][11] != ele[14][11];
    ele[11][11] != ele[14][12];
    ele[11][11] != ele[14][13];
    ele[11][11] != ele[14][14];
    ele[11][11] != ele[15][11];
    ele[11][11] != ele[16][11];
    ele[11][11] != ele[17][11];
    ele[11][11] != ele[18][11];
    ele[11][11] != ele[19][11];
    ele[11][11] != ele[20][11];
    ele[11][11] != ele[21][11];
    ele[11][11] != ele[22][11];
    ele[11][11] != ele[23][11];
    ele[11][11] != ele[24][11];
    ele[11][12] != ele[11][13];
    ele[11][12] != ele[11][14];
    ele[11][12] != ele[11][15];
    ele[11][12] != ele[11][16];
    ele[11][12] != ele[11][17];
    ele[11][12] != ele[11][18];
    ele[11][12] != ele[11][19];
    ele[11][12] != ele[11][20];
    ele[11][12] != ele[11][21];
    ele[11][12] != ele[11][22];
    ele[11][12] != ele[11][23];
    ele[11][12] != ele[11][24];
    ele[11][12] != ele[12][10];
    ele[11][12] != ele[12][11];
    ele[11][12] != ele[12][12];
    ele[11][12] != ele[12][13];
    ele[11][12] != ele[12][14];
    ele[11][12] != ele[13][10];
    ele[11][12] != ele[13][11];
    ele[11][12] != ele[13][12];
    ele[11][12] != ele[13][13];
    ele[11][12] != ele[13][14];
    ele[11][12] != ele[14][10];
    ele[11][12] != ele[14][11];
    ele[11][12] != ele[14][12];
    ele[11][12] != ele[14][13];
    ele[11][12] != ele[14][14];
    ele[11][12] != ele[15][12];
    ele[11][12] != ele[16][12];
    ele[11][12] != ele[17][12];
    ele[11][12] != ele[18][12];
    ele[11][12] != ele[19][12];
    ele[11][12] != ele[20][12];
    ele[11][12] != ele[21][12];
    ele[11][12] != ele[22][12];
    ele[11][12] != ele[23][12];
    ele[11][12] != ele[24][12];
    ele[11][13] != ele[11][14];
    ele[11][13] != ele[11][15];
    ele[11][13] != ele[11][16];
    ele[11][13] != ele[11][17];
    ele[11][13] != ele[11][18];
    ele[11][13] != ele[11][19];
    ele[11][13] != ele[11][20];
    ele[11][13] != ele[11][21];
    ele[11][13] != ele[11][22];
    ele[11][13] != ele[11][23];
    ele[11][13] != ele[11][24];
    ele[11][13] != ele[12][10];
    ele[11][13] != ele[12][11];
    ele[11][13] != ele[12][12];
    ele[11][13] != ele[12][13];
    ele[11][13] != ele[12][14];
    ele[11][13] != ele[13][10];
    ele[11][13] != ele[13][11];
    ele[11][13] != ele[13][12];
    ele[11][13] != ele[13][13];
    ele[11][13] != ele[13][14];
    ele[11][13] != ele[14][10];
    ele[11][13] != ele[14][11];
    ele[11][13] != ele[14][12];
    ele[11][13] != ele[14][13];
    ele[11][13] != ele[14][14];
    ele[11][13] != ele[15][13];
    ele[11][13] != ele[16][13];
    ele[11][13] != ele[17][13];
    ele[11][13] != ele[18][13];
    ele[11][13] != ele[19][13];
    ele[11][13] != ele[20][13];
    ele[11][13] != ele[21][13];
    ele[11][13] != ele[22][13];
    ele[11][13] != ele[23][13];
    ele[11][13] != ele[24][13];
    ele[11][14] != ele[11][15];
    ele[11][14] != ele[11][16];
    ele[11][14] != ele[11][17];
    ele[11][14] != ele[11][18];
    ele[11][14] != ele[11][19];
    ele[11][14] != ele[11][20];
    ele[11][14] != ele[11][21];
    ele[11][14] != ele[11][22];
    ele[11][14] != ele[11][23];
    ele[11][14] != ele[11][24];
    ele[11][14] != ele[12][10];
    ele[11][14] != ele[12][11];
    ele[11][14] != ele[12][12];
    ele[11][14] != ele[12][13];
    ele[11][14] != ele[12][14];
    ele[11][14] != ele[13][10];
    ele[11][14] != ele[13][11];
    ele[11][14] != ele[13][12];
    ele[11][14] != ele[13][13];
    ele[11][14] != ele[13][14];
    ele[11][14] != ele[14][10];
    ele[11][14] != ele[14][11];
    ele[11][14] != ele[14][12];
    ele[11][14] != ele[14][13];
    ele[11][14] != ele[14][14];
    ele[11][14] != ele[15][14];
    ele[11][14] != ele[16][14];
    ele[11][14] != ele[17][14];
    ele[11][14] != ele[18][14];
    ele[11][14] != ele[19][14];
    ele[11][14] != ele[20][14];
    ele[11][14] != ele[21][14];
    ele[11][14] != ele[22][14];
    ele[11][14] != ele[23][14];
    ele[11][14] != ele[24][14];
    ele[11][15] != ele[11][16];
    ele[11][15] != ele[11][17];
    ele[11][15] != ele[11][18];
    ele[11][15] != ele[11][19];
    ele[11][15] != ele[11][20];
    ele[11][15] != ele[11][21];
    ele[11][15] != ele[11][22];
    ele[11][15] != ele[11][23];
    ele[11][15] != ele[11][24];
    ele[11][15] != ele[12][15];
    ele[11][15] != ele[12][16];
    ele[11][15] != ele[12][17];
    ele[11][15] != ele[12][18];
    ele[11][15] != ele[12][19];
    ele[11][15] != ele[13][15];
    ele[11][15] != ele[13][16];
    ele[11][15] != ele[13][17];
    ele[11][15] != ele[13][18];
    ele[11][15] != ele[13][19];
    ele[11][15] != ele[14][15];
    ele[11][15] != ele[14][16];
    ele[11][15] != ele[14][17];
    ele[11][15] != ele[14][18];
    ele[11][15] != ele[14][19];
    ele[11][15] != ele[15][15];
    ele[11][15] != ele[16][15];
    ele[11][15] != ele[17][15];
    ele[11][15] != ele[18][15];
    ele[11][15] != ele[19][15];
    ele[11][15] != ele[20][15];
    ele[11][15] != ele[21][15];
    ele[11][15] != ele[22][15];
    ele[11][15] != ele[23][15];
    ele[11][15] != ele[24][15];
    ele[11][16] != ele[11][17];
    ele[11][16] != ele[11][18];
    ele[11][16] != ele[11][19];
    ele[11][16] != ele[11][20];
    ele[11][16] != ele[11][21];
    ele[11][16] != ele[11][22];
    ele[11][16] != ele[11][23];
    ele[11][16] != ele[11][24];
    ele[11][16] != ele[12][15];
    ele[11][16] != ele[12][16];
    ele[11][16] != ele[12][17];
    ele[11][16] != ele[12][18];
    ele[11][16] != ele[12][19];
    ele[11][16] != ele[13][15];
    ele[11][16] != ele[13][16];
    ele[11][16] != ele[13][17];
    ele[11][16] != ele[13][18];
    ele[11][16] != ele[13][19];
    ele[11][16] != ele[14][15];
    ele[11][16] != ele[14][16];
    ele[11][16] != ele[14][17];
    ele[11][16] != ele[14][18];
    ele[11][16] != ele[14][19];
    ele[11][16] != ele[15][16];
    ele[11][16] != ele[16][16];
    ele[11][16] != ele[17][16];
    ele[11][16] != ele[18][16];
    ele[11][16] != ele[19][16];
    ele[11][16] != ele[20][16];
    ele[11][16] != ele[21][16];
    ele[11][16] != ele[22][16];
    ele[11][16] != ele[23][16];
    ele[11][16] != ele[24][16];
    ele[11][17] != ele[11][18];
    ele[11][17] != ele[11][19];
    ele[11][17] != ele[11][20];
    ele[11][17] != ele[11][21];
    ele[11][17] != ele[11][22];
    ele[11][17] != ele[11][23];
    ele[11][17] != ele[11][24];
    ele[11][17] != ele[12][15];
    ele[11][17] != ele[12][16];
    ele[11][17] != ele[12][17];
    ele[11][17] != ele[12][18];
    ele[11][17] != ele[12][19];
    ele[11][17] != ele[13][15];
    ele[11][17] != ele[13][16];
    ele[11][17] != ele[13][17];
    ele[11][17] != ele[13][18];
    ele[11][17] != ele[13][19];
    ele[11][17] != ele[14][15];
    ele[11][17] != ele[14][16];
    ele[11][17] != ele[14][17];
    ele[11][17] != ele[14][18];
    ele[11][17] != ele[14][19];
    ele[11][17] != ele[15][17];
    ele[11][17] != ele[16][17];
    ele[11][17] != ele[17][17];
    ele[11][17] != ele[18][17];
    ele[11][17] != ele[19][17];
    ele[11][17] != ele[20][17];
    ele[11][17] != ele[21][17];
    ele[11][17] != ele[22][17];
    ele[11][17] != ele[23][17];
    ele[11][17] != ele[24][17];
    ele[11][18] != ele[11][19];
    ele[11][18] != ele[11][20];
    ele[11][18] != ele[11][21];
    ele[11][18] != ele[11][22];
    ele[11][18] != ele[11][23];
    ele[11][18] != ele[11][24];
    ele[11][18] != ele[12][15];
    ele[11][18] != ele[12][16];
    ele[11][18] != ele[12][17];
    ele[11][18] != ele[12][18];
    ele[11][18] != ele[12][19];
    ele[11][18] != ele[13][15];
    ele[11][18] != ele[13][16];
    ele[11][18] != ele[13][17];
    ele[11][18] != ele[13][18];
    ele[11][18] != ele[13][19];
    ele[11][18] != ele[14][15];
    ele[11][18] != ele[14][16];
    ele[11][18] != ele[14][17];
    ele[11][18] != ele[14][18];
    ele[11][18] != ele[14][19];
    ele[11][18] != ele[15][18];
    ele[11][18] != ele[16][18];
    ele[11][18] != ele[17][18];
    ele[11][18] != ele[18][18];
    ele[11][18] != ele[19][18];
    ele[11][18] != ele[20][18];
    ele[11][18] != ele[21][18];
    ele[11][18] != ele[22][18];
    ele[11][18] != ele[23][18];
    ele[11][18] != ele[24][18];
    ele[11][19] != ele[11][20];
    ele[11][19] != ele[11][21];
    ele[11][19] != ele[11][22];
    ele[11][19] != ele[11][23];
    ele[11][19] != ele[11][24];
    ele[11][19] != ele[12][15];
    ele[11][19] != ele[12][16];
    ele[11][19] != ele[12][17];
    ele[11][19] != ele[12][18];
    ele[11][19] != ele[12][19];
    ele[11][19] != ele[13][15];
    ele[11][19] != ele[13][16];
    ele[11][19] != ele[13][17];
    ele[11][19] != ele[13][18];
    ele[11][19] != ele[13][19];
    ele[11][19] != ele[14][15];
    ele[11][19] != ele[14][16];
    ele[11][19] != ele[14][17];
    ele[11][19] != ele[14][18];
    ele[11][19] != ele[14][19];
    ele[11][19] != ele[15][19];
    ele[11][19] != ele[16][19];
    ele[11][19] != ele[17][19];
    ele[11][19] != ele[18][19];
    ele[11][19] != ele[19][19];
    ele[11][19] != ele[20][19];
    ele[11][19] != ele[21][19];
    ele[11][19] != ele[22][19];
    ele[11][19] != ele[23][19];
    ele[11][19] != ele[24][19];
    ele[11][2] != ele[11][10];
    ele[11][2] != ele[11][11];
    ele[11][2] != ele[11][12];
    ele[11][2] != ele[11][13];
    ele[11][2] != ele[11][14];
    ele[11][2] != ele[11][15];
    ele[11][2] != ele[11][16];
    ele[11][2] != ele[11][17];
    ele[11][2] != ele[11][18];
    ele[11][2] != ele[11][19];
    ele[11][2] != ele[11][20];
    ele[11][2] != ele[11][21];
    ele[11][2] != ele[11][22];
    ele[11][2] != ele[11][23];
    ele[11][2] != ele[11][24];
    ele[11][2] != ele[11][3];
    ele[11][2] != ele[11][4];
    ele[11][2] != ele[11][5];
    ele[11][2] != ele[11][6];
    ele[11][2] != ele[11][7];
    ele[11][2] != ele[11][8];
    ele[11][2] != ele[11][9];
    ele[11][2] != ele[12][0];
    ele[11][2] != ele[12][1];
    ele[11][2] != ele[12][2];
    ele[11][2] != ele[12][3];
    ele[11][2] != ele[12][4];
    ele[11][2] != ele[13][0];
    ele[11][2] != ele[13][1];
    ele[11][2] != ele[13][2];
    ele[11][2] != ele[13][3];
    ele[11][2] != ele[13][4];
    ele[11][2] != ele[14][0];
    ele[11][2] != ele[14][1];
    ele[11][2] != ele[14][2];
    ele[11][2] != ele[14][3];
    ele[11][2] != ele[14][4];
    ele[11][2] != ele[15][2];
    ele[11][2] != ele[16][2];
    ele[11][2] != ele[17][2];
    ele[11][2] != ele[18][2];
    ele[11][2] != ele[19][2];
    ele[11][2] != ele[20][2];
    ele[11][2] != ele[21][2];
    ele[11][2] != ele[22][2];
    ele[11][2] != ele[23][2];
    ele[11][2] != ele[24][2];
    ele[11][20] != ele[11][21];
    ele[11][20] != ele[11][22];
    ele[11][20] != ele[11][23];
    ele[11][20] != ele[11][24];
    ele[11][20] != ele[12][20];
    ele[11][20] != ele[12][21];
    ele[11][20] != ele[12][22];
    ele[11][20] != ele[12][23];
    ele[11][20] != ele[12][24];
    ele[11][20] != ele[13][20];
    ele[11][20] != ele[13][21];
    ele[11][20] != ele[13][22];
    ele[11][20] != ele[13][23];
    ele[11][20] != ele[13][24];
    ele[11][20] != ele[14][20];
    ele[11][20] != ele[14][21];
    ele[11][20] != ele[14][22];
    ele[11][20] != ele[14][23];
    ele[11][20] != ele[14][24];
    ele[11][20] != ele[15][20];
    ele[11][20] != ele[16][20];
    ele[11][20] != ele[17][20];
    ele[11][20] != ele[18][20];
    ele[11][20] != ele[19][20];
    ele[11][20] != ele[20][20];
    ele[11][20] != ele[21][20];
    ele[11][20] != ele[22][20];
    ele[11][20] != ele[23][20];
    ele[11][20] != ele[24][20];
    ele[11][21] != ele[11][22];
    ele[11][21] != ele[11][23];
    ele[11][21] != ele[11][24];
    ele[11][21] != ele[12][20];
    ele[11][21] != ele[12][21];
    ele[11][21] != ele[12][22];
    ele[11][21] != ele[12][23];
    ele[11][21] != ele[12][24];
    ele[11][21] != ele[13][20];
    ele[11][21] != ele[13][21];
    ele[11][21] != ele[13][22];
    ele[11][21] != ele[13][23];
    ele[11][21] != ele[13][24];
    ele[11][21] != ele[14][20];
    ele[11][21] != ele[14][21];
    ele[11][21] != ele[14][22];
    ele[11][21] != ele[14][23];
    ele[11][21] != ele[14][24];
    ele[11][21] != ele[15][21];
    ele[11][21] != ele[16][21];
    ele[11][21] != ele[17][21];
    ele[11][21] != ele[18][21];
    ele[11][21] != ele[19][21];
    ele[11][21] != ele[20][21];
    ele[11][21] != ele[21][21];
    ele[11][21] != ele[22][21];
    ele[11][21] != ele[23][21];
    ele[11][21] != ele[24][21];
    ele[11][22] != ele[11][23];
    ele[11][22] != ele[11][24];
    ele[11][22] != ele[12][20];
    ele[11][22] != ele[12][21];
    ele[11][22] != ele[12][22];
    ele[11][22] != ele[12][23];
    ele[11][22] != ele[12][24];
    ele[11][22] != ele[13][20];
    ele[11][22] != ele[13][21];
    ele[11][22] != ele[13][22];
    ele[11][22] != ele[13][23];
    ele[11][22] != ele[13][24];
    ele[11][22] != ele[14][20];
    ele[11][22] != ele[14][21];
    ele[11][22] != ele[14][22];
    ele[11][22] != ele[14][23];
    ele[11][22] != ele[14][24];
    ele[11][22] != ele[15][22];
    ele[11][22] != ele[16][22];
    ele[11][22] != ele[17][22];
    ele[11][22] != ele[18][22];
    ele[11][22] != ele[19][22];
    ele[11][22] != ele[20][22];
    ele[11][22] != ele[21][22];
    ele[11][22] != ele[22][22];
    ele[11][22] != ele[23][22];
    ele[11][22] != ele[24][22];
    ele[11][23] != ele[11][24];
    ele[11][23] != ele[12][20];
    ele[11][23] != ele[12][21];
    ele[11][23] != ele[12][22];
    ele[11][23] != ele[12][23];
    ele[11][23] != ele[12][24];
    ele[11][23] != ele[13][20];
    ele[11][23] != ele[13][21];
    ele[11][23] != ele[13][22];
    ele[11][23] != ele[13][23];
    ele[11][23] != ele[13][24];
    ele[11][23] != ele[14][20];
    ele[11][23] != ele[14][21];
    ele[11][23] != ele[14][22];
    ele[11][23] != ele[14][23];
    ele[11][23] != ele[14][24];
    ele[11][23] != ele[15][23];
    ele[11][23] != ele[16][23];
    ele[11][23] != ele[17][23];
    ele[11][23] != ele[18][23];
    ele[11][23] != ele[19][23];
    ele[11][23] != ele[20][23];
    ele[11][23] != ele[21][23];
    ele[11][23] != ele[22][23];
    ele[11][23] != ele[23][23];
    ele[11][23] != ele[24][23];
    ele[11][24] != ele[12][20];
    ele[11][24] != ele[12][21];
    ele[11][24] != ele[12][22];
    ele[11][24] != ele[12][23];
    ele[11][24] != ele[12][24];
    ele[11][24] != ele[13][20];
    ele[11][24] != ele[13][21];
    ele[11][24] != ele[13][22];
    ele[11][24] != ele[13][23];
    ele[11][24] != ele[13][24];
    ele[11][24] != ele[14][20];
    ele[11][24] != ele[14][21];
    ele[11][24] != ele[14][22];
    ele[11][24] != ele[14][23];
    ele[11][24] != ele[14][24];
    ele[11][24] != ele[15][24];
    ele[11][24] != ele[16][24];
    ele[11][24] != ele[17][24];
    ele[11][24] != ele[18][24];
    ele[11][24] != ele[19][24];
    ele[11][24] != ele[20][24];
    ele[11][24] != ele[21][24];
    ele[11][24] != ele[22][24];
    ele[11][24] != ele[23][24];
    ele[11][24] != ele[24][24];
    ele[11][3] != ele[11][10];
    ele[11][3] != ele[11][11];
    ele[11][3] != ele[11][12];
    ele[11][3] != ele[11][13];
    ele[11][3] != ele[11][14];
    ele[11][3] != ele[11][15];
    ele[11][3] != ele[11][16];
    ele[11][3] != ele[11][17];
    ele[11][3] != ele[11][18];
    ele[11][3] != ele[11][19];
    ele[11][3] != ele[11][20];
    ele[11][3] != ele[11][21];
    ele[11][3] != ele[11][22];
    ele[11][3] != ele[11][23];
    ele[11][3] != ele[11][24];
    ele[11][3] != ele[11][4];
    ele[11][3] != ele[11][5];
    ele[11][3] != ele[11][6];
    ele[11][3] != ele[11][7];
    ele[11][3] != ele[11][8];
    ele[11][3] != ele[11][9];
    ele[11][3] != ele[12][0];
    ele[11][3] != ele[12][1];
    ele[11][3] != ele[12][2];
    ele[11][3] != ele[12][3];
    ele[11][3] != ele[12][4];
    ele[11][3] != ele[13][0];
    ele[11][3] != ele[13][1];
    ele[11][3] != ele[13][2];
    ele[11][3] != ele[13][3];
    ele[11][3] != ele[13][4];
    ele[11][3] != ele[14][0];
    ele[11][3] != ele[14][1];
    ele[11][3] != ele[14][2];
    ele[11][3] != ele[14][3];
    ele[11][3] != ele[14][4];
    ele[11][3] != ele[15][3];
    ele[11][3] != ele[16][3];
    ele[11][3] != ele[17][3];
    ele[11][3] != ele[18][3];
    ele[11][3] != ele[19][3];
    ele[11][3] != ele[20][3];
    ele[11][3] != ele[21][3];
    ele[11][3] != ele[22][3];
    ele[11][3] != ele[23][3];
    ele[11][3] != ele[24][3];
    ele[11][4] != ele[11][10];
    ele[11][4] != ele[11][11];
    ele[11][4] != ele[11][12];
    ele[11][4] != ele[11][13];
    ele[11][4] != ele[11][14];
    ele[11][4] != ele[11][15];
    ele[11][4] != ele[11][16];
    ele[11][4] != ele[11][17];
    ele[11][4] != ele[11][18];
    ele[11][4] != ele[11][19];
    ele[11][4] != ele[11][20];
    ele[11][4] != ele[11][21];
    ele[11][4] != ele[11][22];
    ele[11][4] != ele[11][23];
    ele[11][4] != ele[11][24];
    ele[11][4] != ele[11][5];
    ele[11][4] != ele[11][6];
    ele[11][4] != ele[11][7];
    ele[11][4] != ele[11][8];
    ele[11][4] != ele[11][9];
    ele[11][4] != ele[12][0];
    ele[11][4] != ele[12][1];
    ele[11][4] != ele[12][2];
    ele[11][4] != ele[12][3];
    ele[11][4] != ele[12][4];
    ele[11][4] != ele[13][0];
    ele[11][4] != ele[13][1];
    ele[11][4] != ele[13][2];
    ele[11][4] != ele[13][3];
    ele[11][4] != ele[13][4];
    ele[11][4] != ele[14][0];
    ele[11][4] != ele[14][1];
    ele[11][4] != ele[14][2];
    ele[11][4] != ele[14][3];
    ele[11][4] != ele[14][4];
    ele[11][4] != ele[15][4];
    ele[11][4] != ele[16][4];
    ele[11][4] != ele[17][4];
    ele[11][4] != ele[18][4];
    ele[11][4] != ele[19][4];
    ele[11][4] != ele[20][4];
    ele[11][4] != ele[21][4];
    ele[11][4] != ele[22][4];
    ele[11][4] != ele[23][4];
    ele[11][4] != ele[24][4];
    ele[11][5] != ele[11][10];
    ele[11][5] != ele[11][11];
    ele[11][5] != ele[11][12];
    ele[11][5] != ele[11][13];
    ele[11][5] != ele[11][14];
    ele[11][5] != ele[11][15];
    ele[11][5] != ele[11][16];
    ele[11][5] != ele[11][17];
    ele[11][5] != ele[11][18];
    ele[11][5] != ele[11][19];
    ele[11][5] != ele[11][20];
    ele[11][5] != ele[11][21];
    ele[11][5] != ele[11][22];
    ele[11][5] != ele[11][23];
    ele[11][5] != ele[11][24];
    ele[11][5] != ele[11][6];
    ele[11][5] != ele[11][7];
    ele[11][5] != ele[11][8];
    ele[11][5] != ele[11][9];
    ele[11][5] != ele[12][5];
    ele[11][5] != ele[12][6];
    ele[11][5] != ele[12][7];
    ele[11][5] != ele[12][8];
    ele[11][5] != ele[12][9];
    ele[11][5] != ele[13][5];
    ele[11][5] != ele[13][6];
    ele[11][5] != ele[13][7];
    ele[11][5] != ele[13][8];
    ele[11][5] != ele[13][9];
    ele[11][5] != ele[14][5];
    ele[11][5] != ele[14][6];
    ele[11][5] != ele[14][7];
    ele[11][5] != ele[14][8];
    ele[11][5] != ele[14][9];
    ele[11][5] != ele[15][5];
    ele[11][5] != ele[16][5];
    ele[11][5] != ele[17][5];
    ele[11][5] != ele[18][5];
    ele[11][5] != ele[19][5];
    ele[11][5] != ele[20][5];
    ele[11][5] != ele[21][5];
    ele[11][5] != ele[22][5];
    ele[11][5] != ele[23][5];
    ele[11][5] != ele[24][5];
    ele[11][6] != ele[11][10];
    ele[11][6] != ele[11][11];
    ele[11][6] != ele[11][12];
    ele[11][6] != ele[11][13];
    ele[11][6] != ele[11][14];
    ele[11][6] != ele[11][15];
    ele[11][6] != ele[11][16];
    ele[11][6] != ele[11][17];
    ele[11][6] != ele[11][18];
    ele[11][6] != ele[11][19];
    ele[11][6] != ele[11][20];
    ele[11][6] != ele[11][21];
    ele[11][6] != ele[11][22];
    ele[11][6] != ele[11][23];
    ele[11][6] != ele[11][24];
    ele[11][6] != ele[11][7];
    ele[11][6] != ele[11][8];
    ele[11][6] != ele[11][9];
    ele[11][6] != ele[12][5];
    ele[11][6] != ele[12][6];
    ele[11][6] != ele[12][7];
    ele[11][6] != ele[12][8];
    ele[11][6] != ele[12][9];
    ele[11][6] != ele[13][5];
    ele[11][6] != ele[13][6];
    ele[11][6] != ele[13][7];
    ele[11][6] != ele[13][8];
    ele[11][6] != ele[13][9];
    ele[11][6] != ele[14][5];
    ele[11][6] != ele[14][6];
    ele[11][6] != ele[14][7];
    ele[11][6] != ele[14][8];
    ele[11][6] != ele[14][9];
    ele[11][6] != ele[15][6];
    ele[11][6] != ele[16][6];
    ele[11][6] != ele[17][6];
    ele[11][6] != ele[18][6];
    ele[11][6] != ele[19][6];
    ele[11][6] != ele[20][6];
    ele[11][6] != ele[21][6];
    ele[11][6] != ele[22][6];
    ele[11][6] != ele[23][6];
    ele[11][6] != ele[24][6];
    ele[11][7] != ele[11][10];
    ele[11][7] != ele[11][11];
    ele[11][7] != ele[11][12];
    ele[11][7] != ele[11][13];
    ele[11][7] != ele[11][14];
    ele[11][7] != ele[11][15];
    ele[11][7] != ele[11][16];
    ele[11][7] != ele[11][17];
    ele[11][7] != ele[11][18];
    ele[11][7] != ele[11][19];
    ele[11][7] != ele[11][20];
    ele[11][7] != ele[11][21];
    ele[11][7] != ele[11][22];
    ele[11][7] != ele[11][23];
    ele[11][7] != ele[11][24];
    ele[11][7] != ele[11][8];
    ele[11][7] != ele[11][9];
    ele[11][7] != ele[12][5];
    ele[11][7] != ele[12][6];
    ele[11][7] != ele[12][7];
    ele[11][7] != ele[12][8];
    ele[11][7] != ele[12][9];
    ele[11][7] != ele[13][5];
    ele[11][7] != ele[13][6];
    ele[11][7] != ele[13][7];
    ele[11][7] != ele[13][8];
    ele[11][7] != ele[13][9];
    ele[11][7] != ele[14][5];
    ele[11][7] != ele[14][6];
    ele[11][7] != ele[14][7];
    ele[11][7] != ele[14][8];
    ele[11][7] != ele[14][9];
    ele[11][7] != ele[15][7];
    ele[11][7] != ele[16][7];
    ele[11][7] != ele[17][7];
    ele[11][7] != ele[18][7];
    ele[11][7] != ele[19][7];
    ele[11][7] != ele[20][7];
    ele[11][7] != ele[21][7];
    ele[11][7] != ele[22][7];
    ele[11][7] != ele[23][7];
    ele[11][7] != ele[24][7];
    ele[11][8] != ele[11][10];
    ele[11][8] != ele[11][11];
    ele[11][8] != ele[11][12];
    ele[11][8] != ele[11][13];
    ele[11][8] != ele[11][14];
    ele[11][8] != ele[11][15];
    ele[11][8] != ele[11][16];
    ele[11][8] != ele[11][17];
    ele[11][8] != ele[11][18];
    ele[11][8] != ele[11][19];
    ele[11][8] != ele[11][20];
    ele[11][8] != ele[11][21];
    ele[11][8] != ele[11][22];
    ele[11][8] != ele[11][23];
    ele[11][8] != ele[11][24];
    ele[11][8] != ele[11][9];
    ele[11][8] != ele[12][5];
    ele[11][8] != ele[12][6];
    ele[11][8] != ele[12][7];
    ele[11][8] != ele[12][8];
    ele[11][8] != ele[12][9];
    ele[11][8] != ele[13][5];
    ele[11][8] != ele[13][6];
    ele[11][8] != ele[13][7];
    ele[11][8] != ele[13][8];
    ele[11][8] != ele[13][9];
    ele[11][8] != ele[14][5];
    ele[11][8] != ele[14][6];
    ele[11][8] != ele[14][7];
    ele[11][8] != ele[14][8];
    ele[11][8] != ele[14][9];
    ele[11][8] != ele[15][8];
    ele[11][8] != ele[16][8];
    ele[11][8] != ele[17][8];
    ele[11][8] != ele[18][8];
    ele[11][8] != ele[19][8];
    ele[11][8] != ele[20][8];
    ele[11][8] != ele[21][8];
    ele[11][8] != ele[22][8];
    ele[11][8] != ele[23][8];
    ele[11][8] != ele[24][8];
    ele[11][9] != ele[11][10];
    ele[11][9] != ele[11][11];
    ele[11][9] != ele[11][12];
    ele[11][9] != ele[11][13];
    ele[11][9] != ele[11][14];
    ele[11][9] != ele[11][15];
    ele[11][9] != ele[11][16];
    ele[11][9] != ele[11][17];
    ele[11][9] != ele[11][18];
    ele[11][9] != ele[11][19];
    ele[11][9] != ele[11][20];
    ele[11][9] != ele[11][21];
    ele[11][9] != ele[11][22];
    ele[11][9] != ele[11][23];
    ele[11][9] != ele[11][24];
    ele[11][9] != ele[12][5];
    ele[11][9] != ele[12][6];
    ele[11][9] != ele[12][7];
    ele[11][9] != ele[12][8];
    ele[11][9] != ele[12][9];
    ele[11][9] != ele[13][5];
    ele[11][9] != ele[13][6];
    ele[11][9] != ele[13][7];
    ele[11][9] != ele[13][8];
    ele[11][9] != ele[13][9];
    ele[11][9] != ele[14][5];
    ele[11][9] != ele[14][6];
    ele[11][9] != ele[14][7];
    ele[11][9] != ele[14][8];
    ele[11][9] != ele[14][9];
    ele[11][9] != ele[15][9];
    ele[11][9] != ele[16][9];
    ele[11][9] != ele[17][9];
    ele[11][9] != ele[18][9];
    ele[11][9] != ele[19][9];
    ele[11][9] != ele[20][9];
    ele[11][9] != ele[21][9];
    ele[11][9] != ele[22][9];
    ele[11][9] != ele[23][9];
    ele[11][9] != ele[24][9];
    ele[12][0] != ele[12][1];
    ele[12][0] != ele[12][10];
    ele[12][0] != ele[12][11];
    ele[12][0] != ele[12][12];
    ele[12][0] != ele[12][13];
    ele[12][0] != ele[12][14];
    ele[12][0] != ele[12][15];
    ele[12][0] != ele[12][16];
    ele[12][0] != ele[12][17];
    ele[12][0] != ele[12][18];
    ele[12][0] != ele[12][19];
    ele[12][0] != ele[12][2];
    ele[12][0] != ele[12][20];
    ele[12][0] != ele[12][21];
    ele[12][0] != ele[12][22];
    ele[12][0] != ele[12][23];
    ele[12][0] != ele[12][24];
    ele[12][0] != ele[12][3];
    ele[12][0] != ele[12][4];
    ele[12][0] != ele[12][5];
    ele[12][0] != ele[12][6];
    ele[12][0] != ele[12][7];
    ele[12][0] != ele[12][8];
    ele[12][0] != ele[12][9];
    ele[12][0] != ele[13][0];
    ele[12][0] != ele[13][1];
    ele[12][0] != ele[13][2];
    ele[12][0] != ele[13][3];
    ele[12][0] != ele[13][4];
    ele[12][0] != ele[14][0];
    ele[12][0] != ele[14][1];
    ele[12][0] != ele[14][2];
    ele[12][0] != ele[14][3];
    ele[12][0] != ele[14][4];
    ele[12][0] != ele[15][0];
    ele[12][0] != ele[16][0];
    ele[12][0] != ele[17][0];
    ele[12][0] != ele[18][0];
    ele[12][0] != ele[19][0];
    ele[12][0] != ele[20][0];
    ele[12][0] != ele[21][0];
    ele[12][0] != ele[22][0];
    ele[12][0] != ele[23][0];
    ele[12][0] != ele[24][0];
    ele[12][1] != ele[12][10];
    ele[12][1] != ele[12][11];
    ele[12][1] != ele[12][12];
    ele[12][1] != ele[12][13];
    ele[12][1] != ele[12][14];
    ele[12][1] != ele[12][15];
    ele[12][1] != ele[12][16];
    ele[12][1] != ele[12][17];
    ele[12][1] != ele[12][18];
    ele[12][1] != ele[12][19];
    ele[12][1] != ele[12][2];
    ele[12][1] != ele[12][20];
    ele[12][1] != ele[12][21];
    ele[12][1] != ele[12][22];
    ele[12][1] != ele[12][23];
    ele[12][1] != ele[12][24];
    ele[12][1] != ele[12][3];
    ele[12][1] != ele[12][4];
    ele[12][1] != ele[12][5];
    ele[12][1] != ele[12][6];
    ele[12][1] != ele[12][7];
    ele[12][1] != ele[12][8];
    ele[12][1] != ele[12][9];
    ele[12][1] != ele[13][0];
    ele[12][1] != ele[13][1];
    ele[12][1] != ele[13][2];
    ele[12][1] != ele[13][3];
    ele[12][1] != ele[13][4];
    ele[12][1] != ele[14][0];
    ele[12][1] != ele[14][1];
    ele[12][1] != ele[14][2];
    ele[12][1] != ele[14][3];
    ele[12][1] != ele[14][4];
    ele[12][1] != ele[15][1];
    ele[12][1] != ele[16][1];
    ele[12][1] != ele[17][1];
    ele[12][1] != ele[18][1];
    ele[12][1] != ele[19][1];
    ele[12][1] != ele[20][1];
    ele[12][1] != ele[21][1];
    ele[12][1] != ele[22][1];
    ele[12][1] != ele[23][1];
    ele[12][1] != ele[24][1];
    ele[12][10] != ele[12][11];
    ele[12][10] != ele[12][12];
    ele[12][10] != ele[12][13];
    ele[12][10] != ele[12][14];
    ele[12][10] != ele[12][15];
    ele[12][10] != ele[12][16];
    ele[12][10] != ele[12][17];
    ele[12][10] != ele[12][18];
    ele[12][10] != ele[12][19];
    ele[12][10] != ele[12][20];
    ele[12][10] != ele[12][21];
    ele[12][10] != ele[12][22];
    ele[12][10] != ele[12][23];
    ele[12][10] != ele[12][24];
    ele[12][10] != ele[13][10];
    ele[12][10] != ele[13][11];
    ele[12][10] != ele[13][12];
    ele[12][10] != ele[13][13];
    ele[12][10] != ele[13][14];
    ele[12][10] != ele[14][10];
    ele[12][10] != ele[14][11];
    ele[12][10] != ele[14][12];
    ele[12][10] != ele[14][13];
    ele[12][10] != ele[14][14];
    ele[12][10] != ele[15][10];
    ele[12][10] != ele[16][10];
    ele[12][10] != ele[17][10];
    ele[12][10] != ele[18][10];
    ele[12][10] != ele[19][10];
    ele[12][10] != ele[20][10];
    ele[12][10] != ele[21][10];
    ele[12][10] != ele[22][10];
    ele[12][10] != ele[23][10];
    ele[12][10] != ele[24][10];
    ele[12][11] != ele[12][12];
    ele[12][11] != ele[12][13];
    ele[12][11] != ele[12][14];
    ele[12][11] != ele[12][15];
    ele[12][11] != ele[12][16];
    ele[12][11] != ele[12][17];
    ele[12][11] != ele[12][18];
    ele[12][11] != ele[12][19];
    ele[12][11] != ele[12][20];
    ele[12][11] != ele[12][21];
    ele[12][11] != ele[12][22];
    ele[12][11] != ele[12][23];
    ele[12][11] != ele[12][24];
    ele[12][11] != ele[13][10];
    ele[12][11] != ele[13][11];
    ele[12][11] != ele[13][12];
    ele[12][11] != ele[13][13];
    ele[12][11] != ele[13][14];
    ele[12][11] != ele[14][10];
    ele[12][11] != ele[14][11];
    ele[12][11] != ele[14][12];
    ele[12][11] != ele[14][13];
    ele[12][11] != ele[14][14];
    ele[12][11] != ele[15][11];
    ele[12][11] != ele[16][11];
    ele[12][11] != ele[17][11];
    ele[12][11] != ele[18][11];
    ele[12][11] != ele[19][11];
    ele[12][11] != ele[20][11];
    ele[12][11] != ele[21][11];
    ele[12][11] != ele[22][11];
    ele[12][11] != ele[23][11];
    ele[12][11] != ele[24][11];
    ele[12][12] != ele[12][13];
    ele[12][12] != ele[12][14];
    ele[12][12] != ele[12][15];
    ele[12][12] != ele[12][16];
    ele[12][12] != ele[12][17];
    ele[12][12] != ele[12][18];
    ele[12][12] != ele[12][19];
    ele[12][12] != ele[12][20];
    ele[12][12] != ele[12][21];
    ele[12][12] != ele[12][22];
    ele[12][12] != ele[12][23];
    ele[12][12] != ele[12][24];
    ele[12][12] != ele[13][10];
    ele[12][12] != ele[13][11];
    ele[12][12] != ele[13][12];
    ele[12][12] != ele[13][13];
    ele[12][12] != ele[13][14];
    ele[12][12] != ele[14][10];
    ele[12][12] != ele[14][11];
    ele[12][12] != ele[14][12];
    ele[12][12] != ele[14][13];
    ele[12][12] != ele[14][14];
    ele[12][12] != ele[15][12];
    ele[12][12] != ele[16][12];
    ele[12][12] != ele[17][12];
    ele[12][12] != ele[18][12];
    ele[12][12] != ele[19][12];
    ele[12][12] != ele[20][12];
    ele[12][12] != ele[21][12];
    ele[12][12] != ele[22][12];
    ele[12][12] != ele[23][12];
    ele[12][12] != ele[24][12];
    ele[12][13] != ele[12][14];
    ele[12][13] != ele[12][15];
    ele[12][13] != ele[12][16];
    ele[12][13] != ele[12][17];
    ele[12][13] != ele[12][18];
    ele[12][13] != ele[12][19];
    ele[12][13] != ele[12][20];
    ele[12][13] != ele[12][21];
    ele[12][13] != ele[12][22];
    ele[12][13] != ele[12][23];
    ele[12][13] != ele[12][24];
    ele[12][13] != ele[13][10];
    ele[12][13] != ele[13][11];
    ele[12][13] != ele[13][12];
    ele[12][13] != ele[13][13];
    ele[12][13] != ele[13][14];
    ele[12][13] != ele[14][10];
    ele[12][13] != ele[14][11];
    ele[12][13] != ele[14][12];
    ele[12][13] != ele[14][13];
    ele[12][13] != ele[14][14];
    ele[12][13] != ele[15][13];
    ele[12][13] != ele[16][13];
    ele[12][13] != ele[17][13];
    ele[12][13] != ele[18][13];
    ele[12][13] != ele[19][13];
    ele[12][13] != ele[20][13];
    ele[12][13] != ele[21][13];
    ele[12][13] != ele[22][13];
    ele[12][13] != ele[23][13];
    ele[12][13] != ele[24][13];
    ele[12][14] != ele[12][15];
    ele[12][14] != ele[12][16];
    ele[12][14] != ele[12][17];
    ele[12][14] != ele[12][18];
    ele[12][14] != ele[12][19];
    ele[12][14] != ele[12][20];
    ele[12][14] != ele[12][21];
    ele[12][14] != ele[12][22];
    ele[12][14] != ele[12][23];
    ele[12][14] != ele[12][24];
    ele[12][14] != ele[13][10];
    ele[12][14] != ele[13][11];
    ele[12][14] != ele[13][12];
    ele[12][14] != ele[13][13];
    ele[12][14] != ele[13][14];
    ele[12][14] != ele[14][10];
    ele[12][14] != ele[14][11];
    ele[12][14] != ele[14][12];
    ele[12][14] != ele[14][13];
    ele[12][14] != ele[14][14];
    ele[12][14] != ele[15][14];
    ele[12][14] != ele[16][14];
    ele[12][14] != ele[17][14];
    ele[12][14] != ele[18][14];
    ele[12][14] != ele[19][14];
    ele[12][14] != ele[20][14];
    ele[12][14] != ele[21][14];
    ele[12][14] != ele[22][14];
    ele[12][14] != ele[23][14];
    ele[12][14] != ele[24][14];
    ele[12][15] != ele[12][16];
    ele[12][15] != ele[12][17];
    ele[12][15] != ele[12][18];
    ele[12][15] != ele[12][19];
    ele[12][15] != ele[12][20];
    ele[12][15] != ele[12][21];
    ele[12][15] != ele[12][22];
    ele[12][15] != ele[12][23];
    ele[12][15] != ele[12][24];
    ele[12][15] != ele[13][15];
    ele[12][15] != ele[13][16];
    ele[12][15] != ele[13][17];
    ele[12][15] != ele[13][18];
    ele[12][15] != ele[13][19];
    ele[12][15] != ele[14][15];
    ele[12][15] != ele[14][16];
    ele[12][15] != ele[14][17];
    ele[12][15] != ele[14][18];
    ele[12][15] != ele[14][19];
    ele[12][15] != ele[15][15];
    ele[12][15] != ele[16][15];
    ele[12][15] != ele[17][15];
    ele[12][15] != ele[18][15];
    ele[12][15] != ele[19][15];
    ele[12][15] != ele[20][15];
    ele[12][15] != ele[21][15];
    ele[12][15] != ele[22][15];
    ele[12][15] != ele[23][15];
    ele[12][15] != ele[24][15];
    ele[12][16] != ele[12][17];
    ele[12][16] != ele[12][18];
    ele[12][16] != ele[12][19];
    ele[12][16] != ele[12][20];
    ele[12][16] != ele[12][21];
    ele[12][16] != ele[12][22];
    ele[12][16] != ele[12][23];
    ele[12][16] != ele[12][24];
    ele[12][16] != ele[13][15];
    ele[12][16] != ele[13][16];
    ele[12][16] != ele[13][17];
    ele[12][16] != ele[13][18];
    ele[12][16] != ele[13][19];
    ele[12][16] != ele[14][15];
    ele[12][16] != ele[14][16];
    ele[12][16] != ele[14][17];
    ele[12][16] != ele[14][18];
    ele[12][16] != ele[14][19];
    ele[12][16] != ele[15][16];
    ele[12][16] != ele[16][16];
    ele[12][16] != ele[17][16];
    ele[12][16] != ele[18][16];
    ele[12][16] != ele[19][16];
    ele[12][16] != ele[20][16];
    ele[12][16] != ele[21][16];
    ele[12][16] != ele[22][16];
    ele[12][16] != ele[23][16];
    ele[12][16] != ele[24][16];
    ele[12][17] != ele[12][18];
    ele[12][17] != ele[12][19];
    ele[12][17] != ele[12][20];
    ele[12][17] != ele[12][21];
    ele[12][17] != ele[12][22];
    ele[12][17] != ele[12][23];
    ele[12][17] != ele[12][24];
    ele[12][17] != ele[13][15];
    ele[12][17] != ele[13][16];
    ele[12][17] != ele[13][17];
    ele[12][17] != ele[13][18];
    ele[12][17] != ele[13][19];
    ele[12][17] != ele[14][15];
    ele[12][17] != ele[14][16];
    ele[12][17] != ele[14][17];
    ele[12][17] != ele[14][18];
    ele[12][17] != ele[14][19];
    ele[12][17] != ele[15][17];
    ele[12][17] != ele[16][17];
    ele[12][17] != ele[17][17];
    ele[12][17] != ele[18][17];
    ele[12][17] != ele[19][17];
    ele[12][17] != ele[20][17];
    ele[12][17] != ele[21][17];
    ele[12][17] != ele[22][17];
    ele[12][17] != ele[23][17];
    ele[12][17] != ele[24][17];
    ele[12][18] != ele[12][19];
    ele[12][18] != ele[12][20];
    ele[12][18] != ele[12][21];
    ele[12][18] != ele[12][22];
    ele[12][18] != ele[12][23];
    ele[12][18] != ele[12][24];
    ele[12][18] != ele[13][15];
    ele[12][18] != ele[13][16];
    ele[12][18] != ele[13][17];
    ele[12][18] != ele[13][18];
    ele[12][18] != ele[13][19];
    ele[12][18] != ele[14][15];
    ele[12][18] != ele[14][16];
    ele[12][18] != ele[14][17];
    ele[12][18] != ele[14][18];
    ele[12][18] != ele[14][19];
    ele[12][18] != ele[15][18];
    ele[12][18] != ele[16][18];
    ele[12][18] != ele[17][18];
    ele[12][18] != ele[18][18];
    ele[12][18] != ele[19][18];
    ele[12][18] != ele[20][18];
    ele[12][18] != ele[21][18];
    ele[12][18] != ele[22][18];
    ele[12][18] != ele[23][18];
    ele[12][18] != ele[24][18];
    ele[12][19] != ele[12][20];
    ele[12][19] != ele[12][21];
    ele[12][19] != ele[12][22];
    ele[12][19] != ele[12][23];
    ele[12][19] != ele[12][24];
    ele[12][19] != ele[13][15];
    ele[12][19] != ele[13][16];
    ele[12][19] != ele[13][17];
    ele[12][19] != ele[13][18];
    ele[12][19] != ele[13][19];
    ele[12][19] != ele[14][15];
    ele[12][19] != ele[14][16];
    ele[12][19] != ele[14][17];
    ele[12][19] != ele[14][18];
    ele[12][19] != ele[14][19];
    ele[12][19] != ele[15][19];
    ele[12][19] != ele[16][19];
    ele[12][19] != ele[17][19];
    ele[12][19] != ele[18][19];
    ele[12][19] != ele[19][19];
    ele[12][19] != ele[20][19];
    ele[12][19] != ele[21][19];
    ele[12][19] != ele[22][19];
    ele[12][19] != ele[23][19];
    ele[12][19] != ele[24][19];
    ele[12][2] != ele[12][10];
    ele[12][2] != ele[12][11];
    ele[12][2] != ele[12][12];
    ele[12][2] != ele[12][13];
    ele[12][2] != ele[12][14];
    ele[12][2] != ele[12][15];
    ele[12][2] != ele[12][16];
    ele[12][2] != ele[12][17];
    ele[12][2] != ele[12][18];
    ele[12][2] != ele[12][19];
    ele[12][2] != ele[12][20];
    ele[12][2] != ele[12][21];
    ele[12][2] != ele[12][22];
    ele[12][2] != ele[12][23];
    ele[12][2] != ele[12][24];
    ele[12][2] != ele[12][3];
    ele[12][2] != ele[12][4];
    ele[12][2] != ele[12][5];
    ele[12][2] != ele[12][6];
    ele[12][2] != ele[12][7];
    ele[12][2] != ele[12][8];
    ele[12][2] != ele[12][9];
    ele[12][2] != ele[13][0];
    ele[12][2] != ele[13][1];
    ele[12][2] != ele[13][2];
    ele[12][2] != ele[13][3];
    ele[12][2] != ele[13][4];
    ele[12][2] != ele[14][0];
    ele[12][2] != ele[14][1];
    ele[12][2] != ele[14][2];
    ele[12][2] != ele[14][3];
    ele[12][2] != ele[14][4];
    ele[12][2] != ele[15][2];
    ele[12][2] != ele[16][2];
    ele[12][2] != ele[17][2];
    ele[12][2] != ele[18][2];
    ele[12][2] != ele[19][2];
    ele[12][2] != ele[20][2];
    ele[12][2] != ele[21][2];
    ele[12][2] != ele[22][2];
    ele[12][2] != ele[23][2];
    ele[12][2] != ele[24][2];
    ele[12][20] != ele[12][21];
    ele[12][20] != ele[12][22];
    ele[12][20] != ele[12][23];
    ele[12][20] != ele[12][24];
    ele[12][20] != ele[13][20];
    ele[12][20] != ele[13][21];
    ele[12][20] != ele[13][22];
    ele[12][20] != ele[13][23];
    ele[12][20] != ele[13][24];
    ele[12][20] != ele[14][20];
    ele[12][20] != ele[14][21];
    ele[12][20] != ele[14][22];
    ele[12][20] != ele[14][23];
    ele[12][20] != ele[14][24];
    ele[12][20] != ele[15][20];
    ele[12][20] != ele[16][20];
    ele[12][20] != ele[17][20];
    ele[12][20] != ele[18][20];
    ele[12][20] != ele[19][20];
    ele[12][20] != ele[20][20];
    ele[12][20] != ele[21][20];
    ele[12][20] != ele[22][20];
    ele[12][20] != ele[23][20];
    ele[12][20] != ele[24][20];
    ele[12][21] != ele[12][22];
    ele[12][21] != ele[12][23];
    ele[12][21] != ele[12][24];
    ele[12][21] != ele[13][20];
    ele[12][21] != ele[13][21];
    ele[12][21] != ele[13][22];
    ele[12][21] != ele[13][23];
    ele[12][21] != ele[13][24];
    ele[12][21] != ele[14][20];
    ele[12][21] != ele[14][21];
    ele[12][21] != ele[14][22];
    ele[12][21] != ele[14][23];
    ele[12][21] != ele[14][24];
    ele[12][21] != ele[15][21];
    ele[12][21] != ele[16][21];
    ele[12][21] != ele[17][21];
    ele[12][21] != ele[18][21];
    ele[12][21] != ele[19][21];
    ele[12][21] != ele[20][21];
    ele[12][21] != ele[21][21];
    ele[12][21] != ele[22][21];
    ele[12][21] != ele[23][21];
    ele[12][21] != ele[24][21];
    ele[12][22] != ele[12][23];
    ele[12][22] != ele[12][24];
    ele[12][22] != ele[13][20];
    ele[12][22] != ele[13][21];
    ele[12][22] != ele[13][22];
    ele[12][22] != ele[13][23];
    ele[12][22] != ele[13][24];
    ele[12][22] != ele[14][20];
    ele[12][22] != ele[14][21];
    ele[12][22] != ele[14][22];
    ele[12][22] != ele[14][23];
    ele[12][22] != ele[14][24];
    ele[12][22] != ele[15][22];
    ele[12][22] != ele[16][22];
    ele[12][22] != ele[17][22];
    ele[12][22] != ele[18][22];
    ele[12][22] != ele[19][22];
    ele[12][22] != ele[20][22];
    ele[12][22] != ele[21][22];
    ele[12][22] != ele[22][22];
    ele[12][22] != ele[23][22];
    ele[12][22] != ele[24][22];
    ele[12][23] != ele[12][24];
    ele[12][23] != ele[13][20];
    ele[12][23] != ele[13][21];
    ele[12][23] != ele[13][22];
    ele[12][23] != ele[13][23];
    ele[12][23] != ele[13][24];
    ele[12][23] != ele[14][20];
    ele[12][23] != ele[14][21];
    ele[12][23] != ele[14][22];
    ele[12][23] != ele[14][23];
    ele[12][23] != ele[14][24];
    ele[12][23] != ele[15][23];
    ele[12][23] != ele[16][23];
    ele[12][23] != ele[17][23];
    ele[12][23] != ele[18][23];
    ele[12][23] != ele[19][23];
    ele[12][23] != ele[20][23];
    ele[12][23] != ele[21][23];
    ele[12][23] != ele[22][23];
    ele[12][23] != ele[23][23];
    ele[12][23] != ele[24][23];
    ele[12][24] != ele[13][20];
    ele[12][24] != ele[13][21];
    ele[12][24] != ele[13][22];
    ele[12][24] != ele[13][23];
    ele[12][24] != ele[13][24];
    ele[12][24] != ele[14][20];
    ele[12][24] != ele[14][21];
    ele[12][24] != ele[14][22];
    ele[12][24] != ele[14][23];
    ele[12][24] != ele[14][24];
    ele[12][24] != ele[15][24];
    ele[12][24] != ele[16][24];
    ele[12][24] != ele[17][24];
    ele[12][24] != ele[18][24];
    ele[12][24] != ele[19][24];
    ele[12][24] != ele[20][24];
    ele[12][24] != ele[21][24];
    ele[12][24] != ele[22][24];
    ele[12][24] != ele[23][24];
    ele[12][24] != ele[24][24];
    ele[12][3] != ele[12][10];
    ele[12][3] != ele[12][11];
    ele[12][3] != ele[12][12];
    ele[12][3] != ele[12][13];
    ele[12][3] != ele[12][14];
    ele[12][3] != ele[12][15];
    ele[12][3] != ele[12][16];
    ele[12][3] != ele[12][17];
    ele[12][3] != ele[12][18];
    ele[12][3] != ele[12][19];
    ele[12][3] != ele[12][20];
    ele[12][3] != ele[12][21];
    ele[12][3] != ele[12][22];
    ele[12][3] != ele[12][23];
    ele[12][3] != ele[12][24];
    ele[12][3] != ele[12][4];
    ele[12][3] != ele[12][5];
    ele[12][3] != ele[12][6];
    ele[12][3] != ele[12][7];
    ele[12][3] != ele[12][8];
    ele[12][3] != ele[12][9];
    ele[12][3] != ele[13][0];
    ele[12][3] != ele[13][1];
    ele[12][3] != ele[13][2];
    ele[12][3] != ele[13][3];
    ele[12][3] != ele[13][4];
    ele[12][3] != ele[14][0];
    ele[12][3] != ele[14][1];
    ele[12][3] != ele[14][2];
    ele[12][3] != ele[14][3];
    ele[12][3] != ele[14][4];
    ele[12][3] != ele[15][3];
    ele[12][3] != ele[16][3];
    ele[12][3] != ele[17][3];
    ele[12][3] != ele[18][3];
    ele[12][3] != ele[19][3];
    ele[12][3] != ele[20][3];
    ele[12][3] != ele[21][3];
    ele[12][3] != ele[22][3];
    ele[12][3] != ele[23][3];
    ele[12][3] != ele[24][3];
    ele[12][4] != ele[12][10];
    ele[12][4] != ele[12][11];
    ele[12][4] != ele[12][12];
    ele[12][4] != ele[12][13];
    ele[12][4] != ele[12][14];
    ele[12][4] != ele[12][15];
    ele[12][4] != ele[12][16];
    ele[12][4] != ele[12][17];
    ele[12][4] != ele[12][18];
    ele[12][4] != ele[12][19];
    ele[12][4] != ele[12][20];
    ele[12][4] != ele[12][21];
    ele[12][4] != ele[12][22];
    ele[12][4] != ele[12][23];
    ele[12][4] != ele[12][24];
    ele[12][4] != ele[12][5];
    ele[12][4] != ele[12][6];
    ele[12][4] != ele[12][7];
    ele[12][4] != ele[12][8];
    ele[12][4] != ele[12][9];
    ele[12][4] != ele[13][0];
    ele[12][4] != ele[13][1];
    ele[12][4] != ele[13][2];
    ele[12][4] != ele[13][3];
    ele[12][4] != ele[13][4];
    ele[12][4] != ele[14][0];
    ele[12][4] != ele[14][1];
    ele[12][4] != ele[14][2];
    ele[12][4] != ele[14][3];
    ele[12][4] != ele[14][4];
    ele[12][4] != ele[15][4];
    ele[12][4] != ele[16][4];
    ele[12][4] != ele[17][4];
    ele[12][4] != ele[18][4];
    ele[12][4] != ele[19][4];
    ele[12][4] != ele[20][4];
    ele[12][4] != ele[21][4];
    ele[12][4] != ele[22][4];
    ele[12][4] != ele[23][4];
    ele[12][4] != ele[24][4];
    ele[12][5] != ele[12][10];
    ele[12][5] != ele[12][11];
    ele[12][5] != ele[12][12];
    ele[12][5] != ele[12][13];
    ele[12][5] != ele[12][14];
    ele[12][5] != ele[12][15];
    ele[12][5] != ele[12][16];
    ele[12][5] != ele[12][17];
    ele[12][5] != ele[12][18];
    ele[12][5] != ele[12][19];
    ele[12][5] != ele[12][20];
    ele[12][5] != ele[12][21];
    ele[12][5] != ele[12][22];
    ele[12][5] != ele[12][23];
    ele[12][5] != ele[12][24];
    ele[12][5] != ele[12][6];
    ele[12][5] != ele[12][7];
    ele[12][5] != ele[12][8];
    ele[12][5] != ele[12][9];
    ele[12][5] != ele[13][5];
    ele[12][5] != ele[13][6];
    ele[12][5] != ele[13][7];
    ele[12][5] != ele[13][8];
    ele[12][5] != ele[13][9];
    ele[12][5] != ele[14][5];
    ele[12][5] != ele[14][6];
    ele[12][5] != ele[14][7];
    ele[12][5] != ele[14][8];
    ele[12][5] != ele[14][9];
    ele[12][5] != ele[15][5];
    ele[12][5] != ele[16][5];
    ele[12][5] != ele[17][5];
    ele[12][5] != ele[18][5];
    ele[12][5] != ele[19][5];
    ele[12][5] != ele[20][5];
    ele[12][5] != ele[21][5];
    ele[12][5] != ele[22][5];
    ele[12][5] != ele[23][5];
    ele[12][5] != ele[24][5];
    ele[12][6] != ele[12][10];
    ele[12][6] != ele[12][11];
    ele[12][6] != ele[12][12];
    ele[12][6] != ele[12][13];
    ele[12][6] != ele[12][14];
    ele[12][6] != ele[12][15];
    ele[12][6] != ele[12][16];
    ele[12][6] != ele[12][17];
    ele[12][6] != ele[12][18];
    ele[12][6] != ele[12][19];
    ele[12][6] != ele[12][20];
    ele[12][6] != ele[12][21];
    ele[12][6] != ele[12][22];
    ele[12][6] != ele[12][23];
    ele[12][6] != ele[12][24];
    ele[12][6] != ele[12][7];
    ele[12][6] != ele[12][8];
    ele[12][6] != ele[12][9];
    ele[12][6] != ele[13][5];
    ele[12][6] != ele[13][6];
    ele[12][6] != ele[13][7];
    ele[12][6] != ele[13][8];
    ele[12][6] != ele[13][9];
    ele[12][6] != ele[14][5];
    ele[12][6] != ele[14][6];
    ele[12][6] != ele[14][7];
    ele[12][6] != ele[14][8];
    ele[12][6] != ele[14][9];
    ele[12][6] != ele[15][6];
    ele[12][6] != ele[16][6];
    ele[12][6] != ele[17][6];
    ele[12][6] != ele[18][6];
    ele[12][6] != ele[19][6];
    ele[12][6] != ele[20][6];
    ele[12][6] != ele[21][6];
    ele[12][6] != ele[22][6];
    ele[12][6] != ele[23][6];
    ele[12][6] != ele[24][6];
    ele[12][7] != ele[12][10];
    ele[12][7] != ele[12][11];
    ele[12][7] != ele[12][12];
    ele[12][7] != ele[12][13];
    ele[12][7] != ele[12][14];
    ele[12][7] != ele[12][15];
    ele[12][7] != ele[12][16];
    ele[12][7] != ele[12][17];
    ele[12][7] != ele[12][18];
    ele[12][7] != ele[12][19];
    ele[12][7] != ele[12][20];
    ele[12][7] != ele[12][21];
    ele[12][7] != ele[12][22];
    ele[12][7] != ele[12][23];
    ele[12][7] != ele[12][24];
    ele[12][7] != ele[12][8];
    ele[12][7] != ele[12][9];
    ele[12][7] != ele[13][5];
    ele[12][7] != ele[13][6];
    ele[12][7] != ele[13][7];
    ele[12][7] != ele[13][8];
    ele[12][7] != ele[13][9];
    ele[12][7] != ele[14][5];
    ele[12][7] != ele[14][6];
    ele[12][7] != ele[14][7];
    ele[12][7] != ele[14][8];
    ele[12][7] != ele[14][9];
    ele[12][7] != ele[15][7];
    ele[12][7] != ele[16][7];
    ele[12][7] != ele[17][7];
    ele[12][7] != ele[18][7];
    ele[12][7] != ele[19][7];
    ele[12][7] != ele[20][7];
    ele[12][7] != ele[21][7];
    ele[12][7] != ele[22][7];
    ele[12][7] != ele[23][7];
    ele[12][7] != ele[24][7];
    ele[12][8] != ele[12][10];
    ele[12][8] != ele[12][11];
    ele[12][8] != ele[12][12];
    ele[12][8] != ele[12][13];
    ele[12][8] != ele[12][14];
    ele[12][8] != ele[12][15];
    ele[12][8] != ele[12][16];
    ele[12][8] != ele[12][17];
    ele[12][8] != ele[12][18];
    ele[12][8] != ele[12][19];
    ele[12][8] != ele[12][20];
    ele[12][8] != ele[12][21];
    ele[12][8] != ele[12][22];
    ele[12][8] != ele[12][23];
    ele[12][8] != ele[12][24];
    ele[12][8] != ele[12][9];
    ele[12][8] != ele[13][5];
    ele[12][8] != ele[13][6];
    ele[12][8] != ele[13][7];
    ele[12][8] != ele[13][8];
    ele[12][8] != ele[13][9];
    ele[12][8] != ele[14][5];
    ele[12][8] != ele[14][6];
    ele[12][8] != ele[14][7];
    ele[12][8] != ele[14][8];
    ele[12][8] != ele[14][9];
    ele[12][8] != ele[15][8];
    ele[12][8] != ele[16][8];
    ele[12][8] != ele[17][8];
    ele[12][8] != ele[18][8];
    ele[12][8] != ele[19][8];
    ele[12][8] != ele[20][8];
    ele[12][8] != ele[21][8];
    ele[12][8] != ele[22][8];
    ele[12][8] != ele[23][8];
    ele[12][8] != ele[24][8];
    ele[12][9] != ele[12][10];
    ele[12][9] != ele[12][11];
    ele[12][9] != ele[12][12];
    ele[12][9] != ele[12][13];
    ele[12][9] != ele[12][14];
    ele[12][9] != ele[12][15];
    ele[12][9] != ele[12][16];
    ele[12][9] != ele[12][17];
    ele[12][9] != ele[12][18];
    ele[12][9] != ele[12][19];
    ele[12][9] != ele[12][20];
    ele[12][9] != ele[12][21];
    ele[12][9] != ele[12][22];
    ele[12][9] != ele[12][23];
    ele[12][9] != ele[12][24];
    ele[12][9] != ele[13][5];
    ele[12][9] != ele[13][6];
    ele[12][9] != ele[13][7];
    ele[12][9] != ele[13][8];
    ele[12][9] != ele[13][9];
    ele[12][9] != ele[14][5];
    ele[12][9] != ele[14][6];
    ele[12][9] != ele[14][7];
    ele[12][9] != ele[14][8];
    ele[12][9] != ele[14][9];
    ele[12][9] != ele[15][9];
    ele[12][9] != ele[16][9];
    ele[12][9] != ele[17][9];
    ele[12][9] != ele[18][9];
    ele[12][9] != ele[19][9];
    ele[12][9] != ele[20][9];
    ele[12][9] != ele[21][9];
    ele[12][9] != ele[22][9];
    ele[12][9] != ele[23][9];
    ele[12][9] != ele[24][9];
    ele[13][0] != ele[13][1];
    ele[13][0] != ele[13][10];
    ele[13][0] != ele[13][11];
    ele[13][0] != ele[13][12];
    ele[13][0] != ele[13][13];
    ele[13][0] != ele[13][14];
    ele[13][0] != ele[13][15];
    ele[13][0] != ele[13][16];
    ele[13][0] != ele[13][17];
    ele[13][0] != ele[13][18];
    ele[13][0] != ele[13][19];
    ele[13][0] != ele[13][2];
    ele[13][0] != ele[13][20];
    ele[13][0] != ele[13][21];
    ele[13][0] != ele[13][22];
    ele[13][0] != ele[13][23];
    ele[13][0] != ele[13][24];
    ele[13][0] != ele[13][3];
    ele[13][0] != ele[13][4];
    ele[13][0] != ele[13][5];
    ele[13][0] != ele[13][6];
    ele[13][0] != ele[13][7];
    ele[13][0] != ele[13][8];
    ele[13][0] != ele[13][9];
    ele[13][0] != ele[14][0];
    ele[13][0] != ele[14][1];
    ele[13][0] != ele[14][2];
    ele[13][0] != ele[14][3];
    ele[13][0] != ele[14][4];
    ele[13][0] != ele[15][0];
    ele[13][0] != ele[16][0];
    ele[13][0] != ele[17][0];
    ele[13][0] != ele[18][0];
    ele[13][0] != ele[19][0];
    ele[13][0] != ele[20][0];
    ele[13][0] != ele[21][0];
    ele[13][0] != ele[22][0];
    ele[13][0] != ele[23][0];
    ele[13][0] != ele[24][0];
    ele[13][1] != ele[13][10];
    ele[13][1] != ele[13][11];
    ele[13][1] != ele[13][12];
    ele[13][1] != ele[13][13];
    ele[13][1] != ele[13][14];
    ele[13][1] != ele[13][15];
    ele[13][1] != ele[13][16];
    ele[13][1] != ele[13][17];
    ele[13][1] != ele[13][18];
    ele[13][1] != ele[13][19];
    ele[13][1] != ele[13][2];
    ele[13][1] != ele[13][20];
    ele[13][1] != ele[13][21];
    ele[13][1] != ele[13][22];
    ele[13][1] != ele[13][23];
    ele[13][1] != ele[13][24];
    ele[13][1] != ele[13][3];
    ele[13][1] != ele[13][4];
    ele[13][1] != ele[13][5];
    ele[13][1] != ele[13][6];
    ele[13][1] != ele[13][7];
    ele[13][1] != ele[13][8];
    ele[13][1] != ele[13][9];
    ele[13][1] != ele[14][0];
    ele[13][1] != ele[14][1];
    ele[13][1] != ele[14][2];
    ele[13][1] != ele[14][3];
    ele[13][1] != ele[14][4];
    ele[13][1] != ele[15][1];
    ele[13][1] != ele[16][1];
    ele[13][1] != ele[17][1];
    ele[13][1] != ele[18][1];
    ele[13][1] != ele[19][1];
    ele[13][1] != ele[20][1];
    ele[13][1] != ele[21][1];
    ele[13][1] != ele[22][1];
    ele[13][1] != ele[23][1];
    ele[13][1] != ele[24][1];
    ele[13][10] != ele[13][11];
    ele[13][10] != ele[13][12];
    ele[13][10] != ele[13][13];
    ele[13][10] != ele[13][14];
    ele[13][10] != ele[13][15];
    ele[13][10] != ele[13][16];
    ele[13][10] != ele[13][17];
    ele[13][10] != ele[13][18];
    ele[13][10] != ele[13][19];
    ele[13][10] != ele[13][20];
    ele[13][10] != ele[13][21];
    ele[13][10] != ele[13][22];
    ele[13][10] != ele[13][23];
    ele[13][10] != ele[13][24];
    ele[13][10] != ele[14][10];
    ele[13][10] != ele[14][11];
    ele[13][10] != ele[14][12];
    ele[13][10] != ele[14][13];
    ele[13][10] != ele[14][14];
    ele[13][10] != ele[15][10];
    ele[13][10] != ele[16][10];
    ele[13][10] != ele[17][10];
    ele[13][10] != ele[18][10];
    ele[13][10] != ele[19][10];
    ele[13][10] != ele[20][10];
    ele[13][10] != ele[21][10];
    ele[13][10] != ele[22][10];
    ele[13][10] != ele[23][10];
    ele[13][10] != ele[24][10];
    ele[13][11] != ele[13][12];
    ele[13][11] != ele[13][13];
    ele[13][11] != ele[13][14];
    ele[13][11] != ele[13][15];
    ele[13][11] != ele[13][16];
    ele[13][11] != ele[13][17];
    ele[13][11] != ele[13][18];
    ele[13][11] != ele[13][19];
    ele[13][11] != ele[13][20];
    ele[13][11] != ele[13][21];
    ele[13][11] != ele[13][22];
    ele[13][11] != ele[13][23];
    ele[13][11] != ele[13][24];
    ele[13][11] != ele[14][10];
    ele[13][11] != ele[14][11];
    ele[13][11] != ele[14][12];
    ele[13][11] != ele[14][13];
    ele[13][11] != ele[14][14];
    ele[13][11] != ele[15][11];
    ele[13][11] != ele[16][11];
    ele[13][11] != ele[17][11];
    ele[13][11] != ele[18][11];
    ele[13][11] != ele[19][11];
    ele[13][11] != ele[20][11];
    ele[13][11] != ele[21][11];
    ele[13][11] != ele[22][11];
    ele[13][11] != ele[23][11];
    ele[13][11] != ele[24][11];
    ele[13][12] != ele[13][13];
    ele[13][12] != ele[13][14];
    ele[13][12] != ele[13][15];
    ele[13][12] != ele[13][16];
    ele[13][12] != ele[13][17];
    ele[13][12] != ele[13][18];
    ele[13][12] != ele[13][19];
    ele[13][12] != ele[13][20];
    ele[13][12] != ele[13][21];
    ele[13][12] != ele[13][22];
    ele[13][12] != ele[13][23];
    ele[13][12] != ele[13][24];
    ele[13][12] != ele[14][10];
    ele[13][12] != ele[14][11];
    ele[13][12] != ele[14][12];
    ele[13][12] != ele[14][13];
    ele[13][12] != ele[14][14];
    ele[13][12] != ele[15][12];
    ele[13][12] != ele[16][12];
    ele[13][12] != ele[17][12];
    ele[13][12] != ele[18][12];
    ele[13][12] != ele[19][12];
    ele[13][12] != ele[20][12];
    ele[13][12] != ele[21][12];
    ele[13][12] != ele[22][12];
    ele[13][12] != ele[23][12];
    ele[13][12] != ele[24][12];
    ele[13][13] != ele[13][14];
    ele[13][13] != ele[13][15];
    ele[13][13] != ele[13][16];
    ele[13][13] != ele[13][17];
    ele[13][13] != ele[13][18];
    ele[13][13] != ele[13][19];
    ele[13][13] != ele[13][20];
    ele[13][13] != ele[13][21];
    ele[13][13] != ele[13][22];
    ele[13][13] != ele[13][23];
    ele[13][13] != ele[13][24];
    ele[13][13] != ele[14][10];
    ele[13][13] != ele[14][11];
    ele[13][13] != ele[14][12];
    ele[13][13] != ele[14][13];
    ele[13][13] != ele[14][14];
    ele[13][13] != ele[15][13];
    ele[13][13] != ele[16][13];
    ele[13][13] != ele[17][13];
    ele[13][13] != ele[18][13];
    ele[13][13] != ele[19][13];
    ele[13][13] != ele[20][13];
    ele[13][13] != ele[21][13];
    ele[13][13] != ele[22][13];
    ele[13][13] != ele[23][13];
    ele[13][13] != ele[24][13];
    ele[13][14] != ele[13][15];
    ele[13][14] != ele[13][16];
    ele[13][14] != ele[13][17];
    ele[13][14] != ele[13][18];
    ele[13][14] != ele[13][19];
    ele[13][14] != ele[13][20];
    ele[13][14] != ele[13][21];
    ele[13][14] != ele[13][22];
    ele[13][14] != ele[13][23];
    ele[13][14] != ele[13][24];
    ele[13][14] != ele[14][10];
    ele[13][14] != ele[14][11];
    ele[13][14] != ele[14][12];
    ele[13][14] != ele[14][13];
    ele[13][14] != ele[14][14];
    ele[13][14] != ele[15][14];
    ele[13][14] != ele[16][14];
    ele[13][14] != ele[17][14];
    ele[13][14] != ele[18][14];
    ele[13][14] != ele[19][14];
    ele[13][14] != ele[20][14];
    ele[13][14] != ele[21][14];
    ele[13][14] != ele[22][14];
    ele[13][14] != ele[23][14];
    ele[13][14] != ele[24][14];
    ele[13][15] != ele[13][16];
    ele[13][15] != ele[13][17];
    ele[13][15] != ele[13][18];
    ele[13][15] != ele[13][19];
    ele[13][15] != ele[13][20];
    ele[13][15] != ele[13][21];
    ele[13][15] != ele[13][22];
    ele[13][15] != ele[13][23];
    ele[13][15] != ele[13][24];
    ele[13][15] != ele[14][15];
    ele[13][15] != ele[14][16];
    ele[13][15] != ele[14][17];
    ele[13][15] != ele[14][18];
    ele[13][15] != ele[14][19];
    ele[13][15] != ele[15][15];
    ele[13][15] != ele[16][15];
    ele[13][15] != ele[17][15];
    ele[13][15] != ele[18][15];
    ele[13][15] != ele[19][15];
    ele[13][15] != ele[20][15];
    ele[13][15] != ele[21][15];
    ele[13][15] != ele[22][15];
    ele[13][15] != ele[23][15];
    ele[13][15] != ele[24][15];
    ele[13][16] != ele[13][17];
    ele[13][16] != ele[13][18];
    ele[13][16] != ele[13][19];
    ele[13][16] != ele[13][20];
    ele[13][16] != ele[13][21];
    ele[13][16] != ele[13][22];
    ele[13][16] != ele[13][23];
    ele[13][16] != ele[13][24];
    ele[13][16] != ele[14][15];
    ele[13][16] != ele[14][16];
    ele[13][16] != ele[14][17];
    ele[13][16] != ele[14][18];
    ele[13][16] != ele[14][19];
    ele[13][16] != ele[15][16];
    ele[13][16] != ele[16][16];
    ele[13][16] != ele[17][16];
    ele[13][16] != ele[18][16];
    ele[13][16] != ele[19][16];
    ele[13][16] != ele[20][16];
    ele[13][16] != ele[21][16];
    ele[13][16] != ele[22][16];
    ele[13][16] != ele[23][16];
    ele[13][16] != ele[24][16];
    ele[13][17] != ele[13][18];
    ele[13][17] != ele[13][19];
    ele[13][17] != ele[13][20];
    ele[13][17] != ele[13][21];
    ele[13][17] != ele[13][22];
    ele[13][17] != ele[13][23];
    ele[13][17] != ele[13][24];
    ele[13][17] != ele[14][15];
    ele[13][17] != ele[14][16];
    ele[13][17] != ele[14][17];
    ele[13][17] != ele[14][18];
    ele[13][17] != ele[14][19];
    ele[13][17] != ele[15][17];
    ele[13][17] != ele[16][17];
    ele[13][17] != ele[17][17];
    ele[13][17] != ele[18][17];
    ele[13][17] != ele[19][17];
    ele[13][17] != ele[20][17];
    ele[13][17] != ele[21][17];
    ele[13][17] != ele[22][17];
    ele[13][17] != ele[23][17];
    ele[13][17] != ele[24][17];
    ele[13][18] != ele[13][19];
    ele[13][18] != ele[13][20];
    ele[13][18] != ele[13][21];
    ele[13][18] != ele[13][22];
    ele[13][18] != ele[13][23];
    ele[13][18] != ele[13][24];
    ele[13][18] != ele[14][15];
    ele[13][18] != ele[14][16];
    ele[13][18] != ele[14][17];
    ele[13][18] != ele[14][18];
    ele[13][18] != ele[14][19];
    ele[13][18] != ele[15][18];
    ele[13][18] != ele[16][18];
    ele[13][18] != ele[17][18];
    ele[13][18] != ele[18][18];
    ele[13][18] != ele[19][18];
    ele[13][18] != ele[20][18];
    ele[13][18] != ele[21][18];
    ele[13][18] != ele[22][18];
    ele[13][18] != ele[23][18];
    ele[13][18] != ele[24][18];
    ele[13][19] != ele[13][20];
    ele[13][19] != ele[13][21];
    ele[13][19] != ele[13][22];
    ele[13][19] != ele[13][23];
    ele[13][19] != ele[13][24];
    ele[13][19] != ele[14][15];
    ele[13][19] != ele[14][16];
    ele[13][19] != ele[14][17];
    ele[13][19] != ele[14][18];
    ele[13][19] != ele[14][19];
    ele[13][19] != ele[15][19];
    ele[13][19] != ele[16][19];
    ele[13][19] != ele[17][19];
    ele[13][19] != ele[18][19];
    ele[13][19] != ele[19][19];
    ele[13][19] != ele[20][19];
    ele[13][19] != ele[21][19];
    ele[13][19] != ele[22][19];
    ele[13][19] != ele[23][19];
    ele[13][19] != ele[24][19];
    ele[13][2] != ele[13][10];
    ele[13][2] != ele[13][11];
    ele[13][2] != ele[13][12];
    ele[13][2] != ele[13][13];
    ele[13][2] != ele[13][14];
    ele[13][2] != ele[13][15];
    ele[13][2] != ele[13][16];
    ele[13][2] != ele[13][17];
    ele[13][2] != ele[13][18];
    ele[13][2] != ele[13][19];
    ele[13][2] != ele[13][20];
    ele[13][2] != ele[13][21];
    ele[13][2] != ele[13][22];
    ele[13][2] != ele[13][23];
    ele[13][2] != ele[13][24];
    ele[13][2] != ele[13][3];
    ele[13][2] != ele[13][4];
    ele[13][2] != ele[13][5];
    ele[13][2] != ele[13][6];
    ele[13][2] != ele[13][7];
    ele[13][2] != ele[13][8];
    ele[13][2] != ele[13][9];
    ele[13][2] != ele[14][0];
    ele[13][2] != ele[14][1];
    ele[13][2] != ele[14][2];
    ele[13][2] != ele[14][3];
    ele[13][2] != ele[14][4];
    ele[13][2] != ele[15][2];
    ele[13][2] != ele[16][2];
    ele[13][2] != ele[17][2];
    ele[13][2] != ele[18][2];
    ele[13][2] != ele[19][2];
    ele[13][2] != ele[20][2];
    ele[13][2] != ele[21][2];
    ele[13][2] != ele[22][2];
    ele[13][2] != ele[23][2];
    ele[13][2] != ele[24][2];
    ele[13][20] != ele[13][21];
    ele[13][20] != ele[13][22];
    ele[13][20] != ele[13][23];
    ele[13][20] != ele[13][24];
    ele[13][20] != ele[14][20];
    ele[13][20] != ele[14][21];
    ele[13][20] != ele[14][22];
    ele[13][20] != ele[14][23];
    ele[13][20] != ele[14][24];
    ele[13][20] != ele[15][20];
    ele[13][20] != ele[16][20];
    ele[13][20] != ele[17][20];
    ele[13][20] != ele[18][20];
    ele[13][20] != ele[19][20];
    ele[13][20] != ele[20][20];
    ele[13][20] != ele[21][20];
    ele[13][20] != ele[22][20];
    ele[13][20] != ele[23][20];
    ele[13][20] != ele[24][20];
    ele[13][21] != ele[13][22];
    ele[13][21] != ele[13][23];
    ele[13][21] != ele[13][24];
    ele[13][21] != ele[14][20];
    ele[13][21] != ele[14][21];
    ele[13][21] != ele[14][22];
    ele[13][21] != ele[14][23];
    ele[13][21] != ele[14][24];
    ele[13][21] != ele[15][21];
    ele[13][21] != ele[16][21];
    ele[13][21] != ele[17][21];
    ele[13][21] != ele[18][21];
    ele[13][21] != ele[19][21];
    ele[13][21] != ele[20][21];
    ele[13][21] != ele[21][21];
    ele[13][21] != ele[22][21];
    ele[13][21] != ele[23][21];
    ele[13][21] != ele[24][21];
    ele[13][22] != ele[13][23];
    ele[13][22] != ele[13][24];
    ele[13][22] != ele[14][20];
    ele[13][22] != ele[14][21];
    ele[13][22] != ele[14][22];
    ele[13][22] != ele[14][23];
    ele[13][22] != ele[14][24];
    ele[13][22] != ele[15][22];
    ele[13][22] != ele[16][22];
    ele[13][22] != ele[17][22];
    ele[13][22] != ele[18][22];
    ele[13][22] != ele[19][22];
    ele[13][22] != ele[20][22];
    ele[13][22] != ele[21][22];
    ele[13][22] != ele[22][22];
    ele[13][22] != ele[23][22];
    ele[13][22] != ele[24][22];
    ele[13][23] != ele[13][24];
    ele[13][23] != ele[14][20];
    ele[13][23] != ele[14][21];
    ele[13][23] != ele[14][22];
    ele[13][23] != ele[14][23];
    ele[13][23] != ele[14][24];
    ele[13][23] != ele[15][23];
    ele[13][23] != ele[16][23];
    ele[13][23] != ele[17][23];
    ele[13][23] != ele[18][23];
    ele[13][23] != ele[19][23];
    ele[13][23] != ele[20][23];
    ele[13][23] != ele[21][23];
    ele[13][23] != ele[22][23];
    ele[13][23] != ele[23][23];
    ele[13][23] != ele[24][23];
    ele[13][24] != ele[14][20];
    ele[13][24] != ele[14][21];
    ele[13][24] != ele[14][22];
    ele[13][24] != ele[14][23];
    ele[13][24] != ele[14][24];
    ele[13][24] != ele[15][24];
    ele[13][24] != ele[16][24];
    ele[13][24] != ele[17][24];
    ele[13][24] != ele[18][24];
    ele[13][24] != ele[19][24];
    ele[13][24] != ele[20][24];
    ele[13][24] != ele[21][24];
    ele[13][24] != ele[22][24];
    ele[13][24] != ele[23][24];
    ele[13][24] != ele[24][24];
    ele[13][3] != ele[13][10];
    ele[13][3] != ele[13][11];
    ele[13][3] != ele[13][12];
    ele[13][3] != ele[13][13];
    ele[13][3] != ele[13][14];
    ele[13][3] != ele[13][15];
    ele[13][3] != ele[13][16];
    ele[13][3] != ele[13][17];
    ele[13][3] != ele[13][18];
    ele[13][3] != ele[13][19];
    ele[13][3] != ele[13][20];
    ele[13][3] != ele[13][21];
    ele[13][3] != ele[13][22];
    ele[13][3] != ele[13][23];
    ele[13][3] != ele[13][24];
    ele[13][3] != ele[13][4];
    ele[13][3] != ele[13][5];
    ele[13][3] != ele[13][6];
    ele[13][3] != ele[13][7];
    ele[13][3] != ele[13][8];
    ele[13][3] != ele[13][9];
    ele[13][3] != ele[14][0];
    ele[13][3] != ele[14][1];
    ele[13][3] != ele[14][2];
    ele[13][3] != ele[14][3];
    ele[13][3] != ele[14][4];
    ele[13][3] != ele[15][3];
    ele[13][3] != ele[16][3];
    ele[13][3] != ele[17][3];
    ele[13][3] != ele[18][3];
    ele[13][3] != ele[19][3];
    ele[13][3] != ele[20][3];
    ele[13][3] != ele[21][3];
    ele[13][3] != ele[22][3];
    ele[13][3] != ele[23][3];
    ele[13][3] != ele[24][3];
    ele[13][4] != ele[13][10];
    ele[13][4] != ele[13][11];
    ele[13][4] != ele[13][12];
    ele[13][4] != ele[13][13];
    ele[13][4] != ele[13][14];
    ele[13][4] != ele[13][15];
    ele[13][4] != ele[13][16];
    ele[13][4] != ele[13][17];
    ele[13][4] != ele[13][18];
    ele[13][4] != ele[13][19];
    ele[13][4] != ele[13][20];
    ele[13][4] != ele[13][21];
    ele[13][4] != ele[13][22];
    ele[13][4] != ele[13][23];
    ele[13][4] != ele[13][24];
    ele[13][4] != ele[13][5];
    ele[13][4] != ele[13][6];
    ele[13][4] != ele[13][7];
    ele[13][4] != ele[13][8];
    ele[13][4] != ele[13][9];
    ele[13][4] != ele[14][0];
    ele[13][4] != ele[14][1];
    ele[13][4] != ele[14][2];
    ele[13][4] != ele[14][3];
    ele[13][4] != ele[14][4];
    ele[13][4] != ele[15][4];
    ele[13][4] != ele[16][4];
    ele[13][4] != ele[17][4];
    ele[13][4] != ele[18][4];
    ele[13][4] != ele[19][4];
    ele[13][4] != ele[20][4];
    ele[13][4] != ele[21][4];
    ele[13][4] != ele[22][4];
    ele[13][4] != ele[23][4];
    ele[13][4] != ele[24][4];
    ele[13][5] != ele[13][10];
    ele[13][5] != ele[13][11];
    ele[13][5] != ele[13][12];
    ele[13][5] != ele[13][13];
    ele[13][5] != ele[13][14];
    ele[13][5] != ele[13][15];
    ele[13][5] != ele[13][16];
    ele[13][5] != ele[13][17];
    ele[13][5] != ele[13][18];
    ele[13][5] != ele[13][19];
    ele[13][5] != ele[13][20];
    ele[13][5] != ele[13][21];
    ele[13][5] != ele[13][22];
    ele[13][5] != ele[13][23];
    ele[13][5] != ele[13][24];
    ele[13][5] != ele[13][6];
    ele[13][5] != ele[13][7];
    ele[13][5] != ele[13][8];
    ele[13][5] != ele[13][9];
    ele[13][5] != ele[14][5];
    ele[13][5] != ele[14][6];
    ele[13][5] != ele[14][7];
    ele[13][5] != ele[14][8];
    ele[13][5] != ele[14][9];
    ele[13][5] != ele[15][5];
    ele[13][5] != ele[16][5];
    ele[13][5] != ele[17][5];
    ele[13][5] != ele[18][5];
    ele[13][5] != ele[19][5];
    ele[13][5] != ele[20][5];
    ele[13][5] != ele[21][5];
    ele[13][5] != ele[22][5];
    ele[13][5] != ele[23][5];
    ele[13][5] != ele[24][5];
    ele[13][6] != ele[13][10];
    ele[13][6] != ele[13][11];
    ele[13][6] != ele[13][12];
    ele[13][6] != ele[13][13];
    ele[13][6] != ele[13][14];
    ele[13][6] != ele[13][15];
    ele[13][6] != ele[13][16];
    ele[13][6] != ele[13][17];
    ele[13][6] != ele[13][18];
    ele[13][6] != ele[13][19];
    ele[13][6] != ele[13][20];
    ele[13][6] != ele[13][21];
    ele[13][6] != ele[13][22];
    ele[13][6] != ele[13][23];
    ele[13][6] != ele[13][24];
    ele[13][6] != ele[13][7];
    ele[13][6] != ele[13][8];
    ele[13][6] != ele[13][9];
    ele[13][6] != ele[14][5];
    ele[13][6] != ele[14][6];
    ele[13][6] != ele[14][7];
    ele[13][6] != ele[14][8];
    ele[13][6] != ele[14][9];
    ele[13][6] != ele[15][6];
    ele[13][6] != ele[16][6];
    ele[13][6] != ele[17][6];
    ele[13][6] != ele[18][6];
    ele[13][6] != ele[19][6];
    ele[13][6] != ele[20][6];
    ele[13][6] != ele[21][6];
    ele[13][6] != ele[22][6];
    ele[13][6] != ele[23][6];
    ele[13][6] != ele[24][6];
    ele[13][7] != ele[13][10];
    ele[13][7] != ele[13][11];
    ele[13][7] != ele[13][12];
    ele[13][7] != ele[13][13];
    ele[13][7] != ele[13][14];
    ele[13][7] != ele[13][15];
    ele[13][7] != ele[13][16];
    ele[13][7] != ele[13][17];
    ele[13][7] != ele[13][18];
    ele[13][7] != ele[13][19];
    ele[13][7] != ele[13][20];
    ele[13][7] != ele[13][21];
    ele[13][7] != ele[13][22];
    ele[13][7] != ele[13][23];
    ele[13][7] != ele[13][24];
    ele[13][7] != ele[13][8];
    ele[13][7] != ele[13][9];
    ele[13][7] != ele[14][5];
    ele[13][7] != ele[14][6];
    ele[13][7] != ele[14][7];
    ele[13][7] != ele[14][8];
    ele[13][7] != ele[14][9];
    ele[13][7] != ele[15][7];
    ele[13][7] != ele[16][7];
    ele[13][7] != ele[17][7];
    ele[13][7] != ele[18][7];
    ele[13][7] != ele[19][7];
    ele[13][7] != ele[20][7];
    ele[13][7] != ele[21][7];
    ele[13][7] != ele[22][7];
    ele[13][7] != ele[23][7];
    ele[13][7] != ele[24][7];
    ele[13][8] != ele[13][10];
    ele[13][8] != ele[13][11];
    ele[13][8] != ele[13][12];
    ele[13][8] != ele[13][13];
    ele[13][8] != ele[13][14];
    ele[13][8] != ele[13][15];
    ele[13][8] != ele[13][16];
    ele[13][8] != ele[13][17];
    ele[13][8] != ele[13][18];
    ele[13][8] != ele[13][19];
    ele[13][8] != ele[13][20];
    ele[13][8] != ele[13][21];
    ele[13][8] != ele[13][22];
    ele[13][8] != ele[13][23];
    ele[13][8] != ele[13][24];
    ele[13][8] != ele[13][9];
    ele[13][8] != ele[14][5];
    ele[13][8] != ele[14][6];
    ele[13][8] != ele[14][7];
    ele[13][8] != ele[14][8];
    ele[13][8] != ele[14][9];
    ele[13][8] != ele[15][8];
    ele[13][8] != ele[16][8];
    ele[13][8] != ele[17][8];
    ele[13][8] != ele[18][8];
    ele[13][8] != ele[19][8];
    ele[13][8] != ele[20][8];
    ele[13][8] != ele[21][8];
    ele[13][8] != ele[22][8];
    ele[13][8] != ele[23][8];
    ele[13][8] != ele[24][8];
    ele[13][9] != ele[13][10];
    ele[13][9] != ele[13][11];
    ele[13][9] != ele[13][12];
    ele[13][9] != ele[13][13];
    ele[13][9] != ele[13][14];
    ele[13][9] != ele[13][15];
    ele[13][9] != ele[13][16];
    ele[13][9] != ele[13][17];
    ele[13][9] != ele[13][18];
    ele[13][9] != ele[13][19];
    ele[13][9] != ele[13][20];
    ele[13][9] != ele[13][21];
    ele[13][9] != ele[13][22];
    ele[13][9] != ele[13][23];
    ele[13][9] != ele[13][24];
    ele[13][9] != ele[14][5];
    ele[13][9] != ele[14][6];
    ele[13][9] != ele[14][7];
    ele[13][9] != ele[14][8];
    ele[13][9] != ele[14][9];
    ele[13][9] != ele[15][9];
    ele[13][9] != ele[16][9];
    ele[13][9] != ele[17][9];
    ele[13][9] != ele[18][9];
    ele[13][9] != ele[19][9];
    ele[13][9] != ele[20][9];
    ele[13][9] != ele[21][9];
    ele[13][9] != ele[22][9];
    ele[13][9] != ele[23][9];
    ele[13][9] != ele[24][9];
    ele[14][0] != ele[14][1];
    ele[14][0] != ele[14][10];
    ele[14][0] != ele[14][11];
    ele[14][0] != ele[14][12];
    ele[14][0] != ele[14][13];
    ele[14][0] != ele[14][14];
    ele[14][0] != ele[14][15];
    ele[14][0] != ele[14][16];
    ele[14][0] != ele[14][17];
    ele[14][0] != ele[14][18];
    ele[14][0] != ele[14][19];
    ele[14][0] != ele[14][2];
    ele[14][0] != ele[14][20];
    ele[14][0] != ele[14][21];
    ele[14][0] != ele[14][22];
    ele[14][0] != ele[14][23];
    ele[14][0] != ele[14][24];
    ele[14][0] != ele[14][3];
    ele[14][0] != ele[14][4];
    ele[14][0] != ele[14][5];
    ele[14][0] != ele[14][6];
    ele[14][0] != ele[14][7];
    ele[14][0] != ele[14][8];
    ele[14][0] != ele[14][9];
    ele[14][0] != ele[15][0];
    ele[14][0] != ele[16][0];
    ele[14][0] != ele[17][0];
    ele[14][0] != ele[18][0];
    ele[14][0] != ele[19][0];
    ele[14][0] != ele[20][0];
    ele[14][0] != ele[21][0];
    ele[14][0] != ele[22][0];
    ele[14][0] != ele[23][0];
    ele[14][0] != ele[24][0];
    ele[14][1] != ele[14][10];
    ele[14][1] != ele[14][11];
    ele[14][1] != ele[14][12];
    ele[14][1] != ele[14][13];
    ele[14][1] != ele[14][14];
    ele[14][1] != ele[14][15];
    ele[14][1] != ele[14][16];
    ele[14][1] != ele[14][17];
    ele[14][1] != ele[14][18];
    ele[14][1] != ele[14][19];
    ele[14][1] != ele[14][2];
    ele[14][1] != ele[14][20];
    ele[14][1] != ele[14][21];
    ele[14][1] != ele[14][22];
    ele[14][1] != ele[14][23];
    ele[14][1] != ele[14][24];
    ele[14][1] != ele[14][3];
    ele[14][1] != ele[14][4];
    ele[14][1] != ele[14][5];
    ele[14][1] != ele[14][6];
    ele[14][1] != ele[14][7];
    ele[14][1] != ele[14][8];
    ele[14][1] != ele[14][9];
    ele[14][1] != ele[15][1];
    ele[14][1] != ele[16][1];
    ele[14][1] != ele[17][1];
    ele[14][1] != ele[18][1];
    ele[14][1] != ele[19][1];
    ele[14][1] != ele[20][1];
    ele[14][1] != ele[21][1];
    ele[14][1] != ele[22][1];
    ele[14][1] != ele[23][1];
    ele[14][1] != ele[24][1];
    ele[14][10] != ele[14][11];
    ele[14][10] != ele[14][12];
    ele[14][10] != ele[14][13];
    ele[14][10] != ele[14][14];
    ele[14][10] != ele[14][15];
    ele[14][10] != ele[14][16];
    ele[14][10] != ele[14][17];
    ele[14][10] != ele[14][18];
    ele[14][10] != ele[14][19];
    ele[14][10] != ele[14][20];
    ele[14][10] != ele[14][21];
    ele[14][10] != ele[14][22];
    ele[14][10] != ele[14][23];
    ele[14][10] != ele[14][24];
    ele[14][10] != ele[15][10];
    ele[14][10] != ele[16][10];
    ele[14][10] != ele[17][10];
    ele[14][10] != ele[18][10];
    ele[14][10] != ele[19][10];
    ele[14][10] != ele[20][10];
    ele[14][10] != ele[21][10];
    ele[14][10] != ele[22][10];
    ele[14][10] != ele[23][10];
    ele[14][10] != ele[24][10];
    ele[14][11] != ele[14][12];
    ele[14][11] != ele[14][13];
    ele[14][11] != ele[14][14];
    ele[14][11] != ele[14][15];
    ele[14][11] != ele[14][16];
    ele[14][11] != ele[14][17];
    ele[14][11] != ele[14][18];
    ele[14][11] != ele[14][19];
    ele[14][11] != ele[14][20];
    ele[14][11] != ele[14][21];
    ele[14][11] != ele[14][22];
    ele[14][11] != ele[14][23];
    ele[14][11] != ele[14][24];
    ele[14][11] != ele[15][11];
    ele[14][11] != ele[16][11];
    ele[14][11] != ele[17][11];
    ele[14][11] != ele[18][11];
    ele[14][11] != ele[19][11];
    ele[14][11] != ele[20][11];
    ele[14][11] != ele[21][11];
    ele[14][11] != ele[22][11];
    ele[14][11] != ele[23][11];
    ele[14][11] != ele[24][11];
    ele[14][12] != ele[14][13];
    ele[14][12] != ele[14][14];
    ele[14][12] != ele[14][15];
    ele[14][12] != ele[14][16];
    ele[14][12] != ele[14][17];
    ele[14][12] != ele[14][18];
    ele[14][12] != ele[14][19];
    ele[14][12] != ele[14][20];
    ele[14][12] != ele[14][21];
    ele[14][12] != ele[14][22];
    ele[14][12] != ele[14][23];
    ele[14][12] != ele[14][24];
    ele[14][12] != ele[15][12];
    ele[14][12] != ele[16][12];
    ele[14][12] != ele[17][12];
    ele[14][12] != ele[18][12];
    ele[14][12] != ele[19][12];
    ele[14][12] != ele[20][12];
    ele[14][12] != ele[21][12];
    ele[14][12] != ele[22][12];
    ele[14][12] != ele[23][12];
    ele[14][12] != ele[24][12];
    ele[14][13] != ele[14][14];
    ele[14][13] != ele[14][15];
    ele[14][13] != ele[14][16];
    ele[14][13] != ele[14][17];
    ele[14][13] != ele[14][18];
    ele[14][13] != ele[14][19];
    ele[14][13] != ele[14][20];
    ele[14][13] != ele[14][21];
    ele[14][13] != ele[14][22];
    ele[14][13] != ele[14][23];
    ele[14][13] != ele[14][24];
    ele[14][13] != ele[15][13];
    ele[14][13] != ele[16][13];
    ele[14][13] != ele[17][13];
    ele[14][13] != ele[18][13];
    ele[14][13] != ele[19][13];
    ele[14][13] != ele[20][13];
    ele[14][13] != ele[21][13];
    ele[14][13] != ele[22][13];
    ele[14][13] != ele[23][13];
    ele[14][13] != ele[24][13];
    ele[14][14] != ele[14][15];
    ele[14][14] != ele[14][16];
    ele[14][14] != ele[14][17];
    ele[14][14] != ele[14][18];
    ele[14][14] != ele[14][19];
    ele[14][14] != ele[14][20];
    ele[14][14] != ele[14][21];
    ele[14][14] != ele[14][22];
    ele[14][14] != ele[14][23];
    ele[14][14] != ele[14][24];
    ele[14][14] != ele[15][14];
    ele[14][14] != ele[16][14];
    ele[14][14] != ele[17][14];
    ele[14][14] != ele[18][14];
    ele[14][14] != ele[19][14];
    ele[14][14] != ele[20][14];
    ele[14][14] != ele[21][14];
    ele[14][14] != ele[22][14];
    ele[14][14] != ele[23][14];
    ele[14][14] != ele[24][14];
    ele[14][15] != ele[14][16];
    ele[14][15] != ele[14][17];
    ele[14][15] != ele[14][18];
    ele[14][15] != ele[14][19];
    ele[14][15] != ele[14][20];
    ele[14][15] != ele[14][21];
    ele[14][15] != ele[14][22];
    ele[14][15] != ele[14][23];
    ele[14][15] != ele[14][24];
    ele[14][15] != ele[15][15];
    ele[14][15] != ele[16][15];
    ele[14][15] != ele[17][15];
    ele[14][15] != ele[18][15];
    ele[14][15] != ele[19][15];
    ele[14][15] != ele[20][15];
    ele[14][15] != ele[21][15];
    ele[14][15] != ele[22][15];
    ele[14][15] != ele[23][15];
    ele[14][15] != ele[24][15];
    ele[14][16] != ele[14][17];
    ele[14][16] != ele[14][18];
    ele[14][16] != ele[14][19];
    ele[14][16] != ele[14][20];
    ele[14][16] != ele[14][21];
    ele[14][16] != ele[14][22];
    ele[14][16] != ele[14][23];
    ele[14][16] != ele[14][24];
    ele[14][16] != ele[15][16];
    ele[14][16] != ele[16][16];
    ele[14][16] != ele[17][16];
    ele[14][16] != ele[18][16];
    ele[14][16] != ele[19][16];
    ele[14][16] != ele[20][16];
    ele[14][16] != ele[21][16];
    ele[14][16] != ele[22][16];
    ele[14][16] != ele[23][16];
    ele[14][16] != ele[24][16];
    ele[14][17] != ele[14][18];
    ele[14][17] != ele[14][19];
    ele[14][17] != ele[14][20];
    ele[14][17] != ele[14][21];
    ele[14][17] != ele[14][22];
    ele[14][17] != ele[14][23];
    ele[14][17] != ele[14][24];
    ele[14][17] != ele[15][17];
    ele[14][17] != ele[16][17];
    ele[14][17] != ele[17][17];
    ele[14][17] != ele[18][17];
    ele[14][17] != ele[19][17];
    ele[14][17] != ele[20][17];
    ele[14][17] != ele[21][17];
    ele[14][17] != ele[22][17];
    ele[14][17] != ele[23][17];
    ele[14][17] != ele[24][17];
    ele[14][18] != ele[14][19];
    ele[14][18] != ele[14][20];
    ele[14][18] != ele[14][21];
    ele[14][18] != ele[14][22];
    ele[14][18] != ele[14][23];
    ele[14][18] != ele[14][24];
    ele[14][18] != ele[15][18];
    ele[14][18] != ele[16][18];
    ele[14][18] != ele[17][18];
    ele[14][18] != ele[18][18];
    ele[14][18] != ele[19][18];
    ele[14][18] != ele[20][18];
    ele[14][18] != ele[21][18];
    ele[14][18] != ele[22][18];
    ele[14][18] != ele[23][18];
    ele[14][18] != ele[24][18];
    ele[14][19] != ele[14][20];
    ele[14][19] != ele[14][21];
    ele[14][19] != ele[14][22];
    ele[14][19] != ele[14][23];
    ele[14][19] != ele[14][24];
    ele[14][19] != ele[15][19];
    ele[14][19] != ele[16][19];
    ele[14][19] != ele[17][19];
    ele[14][19] != ele[18][19];
    ele[14][19] != ele[19][19];
    ele[14][19] != ele[20][19];
    ele[14][19] != ele[21][19];
    ele[14][19] != ele[22][19];
    ele[14][19] != ele[23][19];
    ele[14][19] != ele[24][19];
    ele[14][2] != ele[14][10];
    ele[14][2] != ele[14][11];
    ele[14][2] != ele[14][12];
    ele[14][2] != ele[14][13];
    ele[14][2] != ele[14][14];
    ele[14][2] != ele[14][15];
    ele[14][2] != ele[14][16];
    ele[14][2] != ele[14][17];
    ele[14][2] != ele[14][18];
    ele[14][2] != ele[14][19];
    ele[14][2] != ele[14][20];
    ele[14][2] != ele[14][21];
    ele[14][2] != ele[14][22];
    ele[14][2] != ele[14][23];
    ele[14][2] != ele[14][24];
    ele[14][2] != ele[14][3];
    ele[14][2] != ele[14][4];
    ele[14][2] != ele[14][5];
    ele[14][2] != ele[14][6];
    ele[14][2] != ele[14][7];
    ele[14][2] != ele[14][8];
    ele[14][2] != ele[14][9];
    ele[14][2] != ele[15][2];
    ele[14][2] != ele[16][2];
    ele[14][2] != ele[17][2];
    ele[14][2] != ele[18][2];
    ele[14][2] != ele[19][2];
    ele[14][2] != ele[20][2];
    ele[14][2] != ele[21][2];
    ele[14][2] != ele[22][2];
    ele[14][2] != ele[23][2];
    ele[14][2] != ele[24][2];
    ele[14][20] != ele[14][21];
    ele[14][20] != ele[14][22];
    ele[14][20] != ele[14][23];
    ele[14][20] != ele[14][24];
    ele[14][20] != ele[15][20];
    ele[14][20] != ele[16][20];
    ele[14][20] != ele[17][20];
    ele[14][20] != ele[18][20];
    ele[14][20] != ele[19][20];
    ele[14][20] != ele[20][20];
    ele[14][20] != ele[21][20];
    ele[14][20] != ele[22][20];
    ele[14][20] != ele[23][20];
    ele[14][20] != ele[24][20];
    ele[14][21] != ele[14][22];
    ele[14][21] != ele[14][23];
    ele[14][21] != ele[14][24];
    ele[14][21] != ele[15][21];
    ele[14][21] != ele[16][21];
    ele[14][21] != ele[17][21];
    ele[14][21] != ele[18][21];
    ele[14][21] != ele[19][21];
    ele[14][21] != ele[20][21];
    ele[14][21] != ele[21][21];
    ele[14][21] != ele[22][21];
    ele[14][21] != ele[23][21];
    ele[14][21] != ele[24][21];
    ele[14][22] != ele[14][23];
    ele[14][22] != ele[14][24];
    ele[14][22] != ele[15][22];
    ele[14][22] != ele[16][22];
    ele[14][22] != ele[17][22];
    ele[14][22] != ele[18][22];
    ele[14][22] != ele[19][22];
    ele[14][22] != ele[20][22];
    ele[14][22] != ele[21][22];
    ele[14][22] != ele[22][22];
    ele[14][22] != ele[23][22];
    ele[14][22] != ele[24][22];
    ele[14][23] != ele[14][24];
    ele[14][23] != ele[15][23];
    ele[14][23] != ele[16][23];
    ele[14][23] != ele[17][23];
    ele[14][23] != ele[18][23];
    ele[14][23] != ele[19][23];
    ele[14][23] != ele[20][23];
    ele[14][23] != ele[21][23];
    ele[14][23] != ele[22][23];
    ele[14][23] != ele[23][23];
    ele[14][23] != ele[24][23];
    ele[14][24] != ele[15][24];
    ele[14][24] != ele[16][24];
    ele[14][24] != ele[17][24];
    ele[14][24] != ele[18][24];
    ele[14][24] != ele[19][24];
    ele[14][24] != ele[20][24];
    ele[14][24] != ele[21][24];
    ele[14][24] != ele[22][24];
    ele[14][24] != ele[23][24];
    ele[14][24] != ele[24][24];
    ele[14][3] != ele[14][10];
    ele[14][3] != ele[14][11];
    ele[14][3] != ele[14][12];
    ele[14][3] != ele[14][13];
    ele[14][3] != ele[14][14];
    ele[14][3] != ele[14][15];
    ele[14][3] != ele[14][16];
    ele[14][3] != ele[14][17];
    ele[14][3] != ele[14][18];
    ele[14][3] != ele[14][19];
    ele[14][3] != ele[14][20];
    ele[14][3] != ele[14][21];
    ele[14][3] != ele[14][22];
    ele[14][3] != ele[14][23];
    ele[14][3] != ele[14][24];
    ele[14][3] != ele[14][4];
    ele[14][3] != ele[14][5];
    ele[14][3] != ele[14][6];
    ele[14][3] != ele[14][7];
    ele[14][3] != ele[14][8];
    ele[14][3] != ele[14][9];
    ele[14][3] != ele[15][3];
    ele[14][3] != ele[16][3];
    ele[14][3] != ele[17][3];
    ele[14][3] != ele[18][3];
    ele[14][3] != ele[19][3];
    ele[14][3] != ele[20][3];
    ele[14][3] != ele[21][3];
    ele[14][3] != ele[22][3];
    ele[14][3] != ele[23][3];
    ele[14][3] != ele[24][3];
    ele[14][4] != ele[14][10];
    ele[14][4] != ele[14][11];
    ele[14][4] != ele[14][12];
    ele[14][4] != ele[14][13];
    ele[14][4] != ele[14][14];
    ele[14][4] != ele[14][15];
    ele[14][4] != ele[14][16];
    ele[14][4] != ele[14][17];
    ele[14][4] != ele[14][18];
    ele[14][4] != ele[14][19];
    ele[14][4] != ele[14][20];
    ele[14][4] != ele[14][21];
    ele[14][4] != ele[14][22];
    ele[14][4] != ele[14][23];
    ele[14][4] != ele[14][24];
    ele[14][4] != ele[14][5];
    ele[14][4] != ele[14][6];
    ele[14][4] != ele[14][7];
    ele[14][4] != ele[14][8];
    ele[14][4] != ele[14][9];
    ele[14][4] != ele[15][4];
    ele[14][4] != ele[16][4];
    ele[14][4] != ele[17][4];
    ele[14][4] != ele[18][4];
    ele[14][4] != ele[19][4];
    ele[14][4] != ele[20][4];
    ele[14][4] != ele[21][4];
    ele[14][4] != ele[22][4];
    ele[14][4] != ele[23][4];
    ele[14][4] != ele[24][4];
    ele[14][5] != ele[14][10];
    ele[14][5] != ele[14][11];
    ele[14][5] != ele[14][12];
    ele[14][5] != ele[14][13];
    ele[14][5] != ele[14][14];
    ele[14][5] != ele[14][15];
    ele[14][5] != ele[14][16];
    ele[14][5] != ele[14][17];
    ele[14][5] != ele[14][18];
    ele[14][5] != ele[14][19];
    ele[14][5] != ele[14][20];
    ele[14][5] != ele[14][21];
    ele[14][5] != ele[14][22];
    ele[14][5] != ele[14][23];
    ele[14][5] != ele[14][24];
    ele[14][5] != ele[14][6];
    ele[14][5] != ele[14][7];
    ele[14][5] != ele[14][8];
    ele[14][5] != ele[14][9];
    ele[14][5] != ele[15][5];
    ele[14][5] != ele[16][5];
    ele[14][5] != ele[17][5];
    ele[14][5] != ele[18][5];
    ele[14][5] != ele[19][5];
    ele[14][5] != ele[20][5];
    ele[14][5] != ele[21][5];
    ele[14][5] != ele[22][5];
    ele[14][5] != ele[23][5];
    ele[14][5] != ele[24][5];
    ele[14][6] != ele[14][10];
    ele[14][6] != ele[14][11];
    ele[14][6] != ele[14][12];
    ele[14][6] != ele[14][13];
    ele[14][6] != ele[14][14];
    ele[14][6] != ele[14][15];
    ele[14][6] != ele[14][16];
    ele[14][6] != ele[14][17];
    ele[14][6] != ele[14][18];
    ele[14][6] != ele[14][19];
    ele[14][6] != ele[14][20];
    ele[14][6] != ele[14][21];
    ele[14][6] != ele[14][22];
    ele[14][6] != ele[14][23];
    ele[14][6] != ele[14][24];
    ele[14][6] != ele[14][7];
    ele[14][6] != ele[14][8];
    ele[14][6] != ele[14][9];
    ele[14][6] != ele[15][6];
    ele[14][6] != ele[16][6];
    ele[14][6] != ele[17][6];
    ele[14][6] != ele[18][6];
    ele[14][6] != ele[19][6];
    ele[14][6] != ele[20][6];
    ele[14][6] != ele[21][6];
    ele[14][6] != ele[22][6];
    ele[14][6] != ele[23][6];
    ele[14][6] != ele[24][6];
    ele[14][7] != ele[14][10];
    ele[14][7] != ele[14][11];
    ele[14][7] != ele[14][12];
    ele[14][7] != ele[14][13];
    ele[14][7] != ele[14][14];
    ele[14][7] != ele[14][15];
    ele[14][7] != ele[14][16];
    ele[14][7] != ele[14][17];
    ele[14][7] != ele[14][18];
    ele[14][7] != ele[14][19];
    ele[14][7] != ele[14][20];
    ele[14][7] != ele[14][21];
    ele[14][7] != ele[14][22];
    ele[14][7] != ele[14][23];
    ele[14][7] != ele[14][24];
    ele[14][7] != ele[14][8];
    ele[14][7] != ele[14][9];
    ele[14][7] != ele[15][7];
    ele[14][7] != ele[16][7];
    ele[14][7] != ele[17][7];
    ele[14][7] != ele[18][7];
    ele[14][7] != ele[19][7];
    ele[14][7] != ele[20][7];
    ele[14][7] != ele[21][7];
    ele[14][7] != ele[22][7];
    ele[14][7] != ele[23][7];
    ele[14][7] != ele[24][7];
    ele[14][8] != ele[14][10];
    ele[14][8] != ele[14][11];
    ele[14][8] != ele[14][12];
    ele[14][8] != ele[14][13];
    ele[14][8] != ele[14][14];
    ele[14][8] != ele[14][15];
    ele[14][8] != ele[14][16];
    ele[14][8] != ele[14][17];
    ele[14][8] != ele[14][18];
    ele[14][8] != ele[14][19];
    ele[14][8] != ele[14][20];
    ele[14][8] != ele[14][21];
    ele[14][8] != ele[14][22];
    ele[14][8] != ele[14][23];
    ele[14][8] != ele[14][24];
    ele[14][8] != ele[14][9];
    ele[14][8] != ele[15][8];
    ele[14][8] != ele[16][8];
    ele[14][8] != ele[17][8];
    ele[14][8] != ele[18][8];
    ele[14][8] != ele[19][8];
    ele[14][8] != ele[20][8];
    ele[14][8] != ele[21][8];
    ele[14][8] != ele[22][8];
    ele[14][8] != ele[23][8];
    ele[14][8] != ele[24][8];
    ele[14][9] != ele[14][10];
    ele[14][9] != ele[14][11];
    ele[14][9] != ele[14][12];
    ele[14][9] != ele[14][13];
    ele[14][9] != ele[14][14];
    ele[14][9] != ele[14][15];
    ele[14][9] != ele[14][16];
    ele[14][9] != ele[14][17];
    ele[14][9] != ele[14][18];
    ele[14][9] != ele[14][19];
    ele[14][9] != ele[14][20];
    ele[14][9] != ele[14][21];
    ele[14][9] != ele[14][22];
    ele[14][9] != ele[14][23];
    ele[14][9] != ele[14][24];
    ele[14][9] != ele[15][9];
    ele[14][9] != ele[16][9];
    ele[14][9] != ele[17][9];
    ele[14][9] != ele[18][9];
    ele[14][9] != ele[19][9];
    ele[14][9] != ele[20][9];
    ele[14][9] != ele[21][9];
    ele[14][9] != ele[22][9];
    ele[14][9] != ele[23][9];
    ele[14][9] != ele[24][9];
    ele[15][0] != ele[15][1];
    ele[15][0] != ele[15][10];
    ele[15][0] != ele[15][11];
    ele[15][0] != ele[15][12];
    ele[15][0] != ele[15][13];
    ele[15][0] != ele[15][14];
    ele[15][0] != ele[15][15];
    ele[15][0] != ele[15][16];
    ele[15][0] != ele[15][17];
    ele[15][0] != ele[15][18];
    ele[15][0] != ele[15][19];
    ele[15][0] != ele[15][2];
    ele[15][0] != ele[15][20];
    ele[15][0] != ele[15][21];
    ele[15][0] != ele[15][22];
    ele[15][0] != ele[15][23];
    ele[15][0] != ele[15][24];
    ele[15][0] != ele[15][3];
    ele[15][0] != ele[15][4];
    ele[15][0] != ele[15][5];
    ele[15][0] != ele[15][6];
    ele[15][0] != ele[15][7];
    ele[15][0] != ele[15][8];
    ele[15][0] != ele[15][9];
    ele[15][0] != ele[16][0];
    ele[15][0] != ele[16][1];
    ele[15][0] != ele[16][2];
    ele[15][0] != ele[16][3];
    ele[15][0] != ele[16][4];
    ele[15][0] != ele[17][0];
    ele[15][0] != ele[17][1];
    ele[15][0] != ele[17][2];
    ele[15][0] != ele[17][3];
    ele[15][0] != ele[17][4];
    ele[15][0] != ele[18][0];
    ele[15][0] != ele[18][1];
    ele[15][0] != ele[18][2];
    ele[15][0] != ele[18][3];
    ele[15][0] != ele[18][4];
    ele[15][0] != ele[19][0];
    ele[15][0] != ele[19][1];
    ele[15][0] != ele[19][2];
    ele[15][0] != ele[19][3];
    ele[15][0] != ele[19][4];
    ele[15][0] != ele[20][0];
    ele[15][0] != ele[21][0];
    ele[15][0] != ele[22][0];
    ele[15][0] != ele[23][0];
    ele[15][0] != ele[24][0];
    ele[15][1] != ele[15][10];
    ele[15][1] != ele[15][11];
    ele[15][1] != ele[15][12];
    ele[15][1] != ele[15][13];
    ele[15][1] != ele[15][14];
    ele[15][1] != ele[15][15];
    ele[15][1] != ele[15][16];
    ele[15][1] != ele[15][17];
    ele[15][1] != ele[15][18];
    ele[15][1] != ele[15][19];
    ele[15][1] != ele[15][2];
    ele[15][1] != ele[15][20];
    ele[15][1] != ele[15][21];
    ele[15][1] != ele[15][22];
    ele[15][1] != ele[15][23];
    ele[15][1] != ele[15][24];
    ele[15][1] != ele[15][3];
    ele[15][1] != ele[15][4];
    ele[15][1] != ele[15][5];
    ele[15][1] != ele[15][6];
    ele[15][1] != ele[15][7];
    ele[15][1] != ele[15][8];
    ele[15][1] != ele[15][9];
    ele[15][1] != ele[16][0];
    ele[15][1] != ele[16][1];
    ele[15][1] != ele[16][2];
    ele[15][1] != ele[16][3];
    ele[15][1] != ele[16][4];
    ele[15][1] != ele[17][0];
    ele[15][1] != ele[17][1];
    ele[15][1] != ele[17][2];
    ele[15][1] != ele[17][3];
    ele[15][1] != ele[17][4];
    ele[15][1] != ele[18][0];
    ele[15][1] != ele[18][1];
    ele[15][1] != ele[18][2];
    ele[15][1] != ele[18][3];
    ele[15][1] != ele[18][4];
    ele[15][1] != ele[19][0];
    ele[15][1] != ele[19][1];
    ele[15][1] != ele[19][2];
    ele[15][1] != ele[19][3];
    ele[15][1] != ele[19][4];
    ele[15][1] != ele[20][1];
    ele[15][1] != ele[21][1];
    ele[15][1] != ele[22][1];
    ele[15][1] != ele[23][1];
    ele[15][1] != ele[24][1];
    ele[15][10] != ele[15][11];
    ele[15][10] != ele[15][12];
    ele[15][10] != ele[15][13];
    ele[15][10] != ele[15][14];
    ele[15][10] != ele[15][15];
    ele[15][10] != ele[15][16];
    ele[15][10] != ele[15][17];
    ele[15][10] != ele[15][18];
    ele[15][10] != ele[15][19];
    ele[15][10] != ele[15][20];
    ele[15][10] != ele[15][21];
    ele[15][10] != ele[15][22];
    ele[15][10] != ele[15][23];
    ele[15][10] != ele[15][24];
    ele[15][10] != ele[16][10];
    ele[15][10] != ele[16][11];
    ele[15][10] != ele[16][12];
    ele[15][10] != ele[16][13];
    ele[15][10] != ele[16][14];
    ele[15][10] != ele[17][10];
    ele[15][10] != ele[17][11];
    ele[15][10] != ele[17][12];
    ele[15][10] != ele[17][13];
    ele[15][10] != ele[17][14];
    ele[15][10] != ele[18][10];
    ele[15][10] != ele[18][11];
    ele[15][10] != ele[18][12];
    ele[15][10] != ele[18][13];
    ele[15][10] != ele[18][14];
    ele[15][10] != ele[19][10];
    ele[15][10] != ele[19][11];
    ele[15][10] != ele[19][12];
    ele[15][10] != ele[19][13];
    ele[15][10] != ele[19][14];
    ele[15][10] != ele[20][10];
    ele[15][10] != ele[21][10];
    ele[15][10] != ele[22][10];
    ele[15][10] != ele[23][10];
    ele[15][10] != ele[24][10];
    ele[15][11] != ele[15][12];
    ele[15][11] != ele[15][13];
    ele[15][11] != ele[15][14];
    ele[15][11] != ele[15][15];
    ele[15][11] != ele[15][16];
    ele[15][11] != ele[15][17];
    ele[15][11] != ele[15][18];
    ele[15][11] != ele[15][19];
    ele[15][11] != ele[15][20];
    ele[15][11] != ele[15][21];
    ele[15][11] != ele[15][22];
    ele[15][11] != ele[15][23];
    ele[15][11] != ele[15][24];
    ele[15][11] != ele[16][10];
    ele[15][11] != ele[16][11];
    ele[15][11] != ele[16][12];
    ele[15][11] != ele[16][13];
    ele[15][11] != ele[16][14];
    ele[15][11] != ele[17][10];
    ele[15][11] != ele[17][11];
    ele[15][11] != ele[17][12];
    ele[15][11] != ele[17][13];
    ele[15][11] != ele[17][14];
    ele[15][11] != ele[18][10];
    ele[15][11] != ele[18][11];
    ele[15][11] != ele[18][12];
    ele[15][11] != ele[18][13];
    ele[15][11] != ele[18][14];
    ele[15][11] != ele[19][10];
    ele[15][11] != ele[19][11];
    ele[15][11] != ele[19][12];
    ele[15][11] != ele[19][13];
    ele[15][11] != ele[19][14];
    ele[15][11] != ele[20][11];
    ele[15][11] != ele[21][11];
    ele[15][11] != ele[22][11];
    ele[15][11] != ele[23][11];
    ele[15][11] != ele[24][11];
    ele[15][12] != ele[15][13];
    ele[15][12] != ele[15][14];
    ele[15][12] != ele[15][15];
    ele[15][12] != ele[15][16];
    ele[15][12] != ele[15][17];
    ele[15][12] != ele[15][18];
    ele[15][12] != ele[15][19];
    ele[15][12] != ele[15][20];
    ele[15][12] != ele[15][21];
    ele[15][12] != ele[15][22];
    ele[15][12] != ele[15][23];
    ele[15][12] != ele[15][24];
    ele[15][12] != ele[16][10];
    ele[15][12] != ele[16][11];
    ele[15][12] != ele[16][12];
    ele[15][12] != ele[16][13];
    ele[15][12] != ele[16][14];
    ele[15][12] != ele[17][10];
    ele[15][12] != ele[17][11];
    ele[15][12] != ele[17][12];
    ele[15][12] != ele[17][13];
    ele[15][12] != ele[17][14];
    ele[15][12] != ele[18][10];
    ele[15][12] != ele[18][11];
    ele[15][12] != ele[18][12];
    ele[15][12] != ele[18][13];
    ele[15][12] != ele[18][14];
    ele[15][12] != ele[19][10];
    ele[15][12] != ele[19][11];
    ele[15][12] != ele[19][12];
    ele[15][12] != ele[19][13];
    ele[15][12] != ele[19][14];
    ele[15][12] != ele[20][12];
    ele[15][12] != ele[21][12];
    ele[15][12] != ele[22][12];
    ele[15][12] != ele[23][12];
    ele[15][12] != ele[24][12];
    ele[15][13] != ele[15][14];
    ele[15][13] != ele[15][15];
    ele[15][13] != ele[15][16];
    ele[15][13] != ele[15][17];
    ele[15][13] != ele[15][18];
    ele[15][13] != ele[15][19];
    ele[15][13] != ele[15][20];
    ele[15][13] != ele[15][21];
    ele[15][13] != ele[15][22];
    ele[15][13] != ele[15][23];
    ele[15][13] != ele[15][24];
    ele[15][13] != ele[16][10];
    ele[15][13] != ele[16][11];
    ele[15][13] != ele[16][12];
    ele[15][13] != ele[16][13];
    ele[15][13] != ele[16][14];
    ele[15][13] != ele[17][10];
    ele[15][13] != ele[17][11];
    ele[15][13] != ele[17][12];
    ele[15][13] != ele[17][13];
    ele[15][13] != ele[17][14];
    ele[15][13] != ele[18][10];
    ele[15][13] != ele[18][11];
    ele[15][13] != ele[18][12];
    ele[15][13] != ele[18][13];
    ele[15][13] != ele[18][14];
    ele[15][13] != ele[19][10];
    ele[15][13] != ele[19][11];
    ele[15][13] != ele[19][12];
    ele[15][13] != ele[19][13];
    ele[15][13] != ele[19][14];
    ele[15][13] != ele[20][13];
    ele[15][13] != ele[21][13];
    ele[15][13] != ele[22][13];
    ele[15][13] != ele[23][13];
    ele[15][13] != ele[24][13];
    ele[15][14] != ele[15][15];
    ele[15][14] != ele[15][16];
    ele[15][14] != ele[15][17];
    ele[15][14] != ele[15][18];
    ele[15][14] != ele[15][19];
    ele[15][14] != ele[15][20];
    ele[15][14] != ele[15][21];
    ele[15][14] != ele[15][22];
    ele[15][14] != ele[15][23];
    ele[15][14] != ele[15][24];
    ele[15][14] != ele[16][10];
    ele[15][14] != ele[16][11];
    ele[15][14] != ele[16][12];
    ele[15][14] != ele[16][13];
    ele[15][14] != ele[16][14];
    ele[15][14] != ele[17][10];
    ele[15][14] != ele[17][11];
    ele[15][14] != ele[17][12];
    ele[15][14] != ele[17][13];
    ele[15][14] != ele[17][14];
    ele[15][14] != ele[18][10];
    ele[15][14] != ele[18][11];
    ele[15][14] != ele[18][12];
    ele[15][14] != ele[18][13];
    ele[15][14] != ele[18][14];
    ele[15][14] != ele[19][10];
    ele[15][14] != ele[19][11];
    ele[15][14] != ele[19][12];
    ele[15][14] != ele[19][13];
    ele[15][14] != ele[19][14];
    ele[15][14] != ele[20][14];
    ele[15][14] != ele[21][14];
    ele[15][14] != ele[22][14];
    ele[15][14] != ele[23][14];
    ele[15][14] != ele[24][14];
    ele[15][15] != ele[15][16];
    ele[15][15] != ele[15][17];
    ele[15][15] != ele[15][18];
    ele[15][15] != ele[15][19];
    ele[15][15] != ele[15][20];
    ele[15][15] != ele[15][21];
    ele[15][15] != ele[15][22];
    ele[15][15] != ele[15][23];
    ele[15][15] != ele[15][24];
    ele[15][15] != ele[16][15];
    ele[15][15] != ele[16][16];
    ele[15][15] != ele[16][17];
    ele[15][15] != ele[16][18];
    ele[15][15] != ele[16][19];
    ele[15][15] != ele[17][15];
    ele[15][15] != ele[17][16];
    ele[15][15] != ele[17][17];
    ele[15][15] != ele[17][18];
    ele[15][15] != ele[17][19];
    ele[15][15] != ele[18][15];
    ele[15][15] != ele[18][16];
    ele[15][15] != ele[18][17];
    ele[15][15] != ele[18][18];
    ele[15][15] != ele[18][19];
    ele[15][15] != ele[19][15];
    ele[15][15] != ele[19][16];
    ele[15][15] != ele[19][17];
    ele[15][15] != ele[19][18];
    ele[15][15] != ele[19][19];
    ele[15][15] != ele[20][15];
    ele[15][15] != ele[21][15];
    ele[15][15] != ele[22][15];
    ele[15][15] != ele[23][15];
    ele[15][15] != ele[24][15];
    ele[15][16] != ele[15][17];
    ele[15][16] != ele[15][18];
    ele[15][16] != ele[15][19];
    ele[15][16] != ele[15][20];
    ele[15][16] != ele[15][21];
    ele[15][16] != ele[15][22];
    ele[15][16] != ele[15][23];
    ele[15][16] != ele[15][24];
    ele[15][16] != ele[16][15];
    ele[15][16] != ele[16][16];
    ele[15][16] != ele[16][17];
    ele[15][16] != ele[16][18];
    ele[15][16] != ele[16][19];
    ele[15][16] != ele[17][15];
    ele[15][16] != ele[17][16];
    ele[15][16] != ele[17][17];
    ele[15][16] != ele[17][18];
    ele[15][16] != ele[17][19];
    ele[15][16] != ele[18][15];
    ele[15][16] != ele[18][16];
    ele[15][16] != ele[18][17];
    ele[15][16] != ele[18][18];
    ele[15][16] != ele[18][19];
    ele[15][16] != ele[19][15];
    ele[15][16] != ele[19][16];
    ele[15][16] != ele[19][17];
    ele[15][16] != ele[19][18];
    ele[15][16] != ele[19][19];
    ele[15][16] != ele[20][16];
    ele[15][16] != ele[21][16];
    ele[15][16] != ele[22][16];
    ele[15][16] != ele[23][16];
    ele[15][16] != ele[24][16];
    ele[15][17] != ele[15][18];
    ele[15][17] != ele[15][19];
    ele[15][17] != ele[15][20];
    ele[15][17] != ele[15][21];
    ele[15][17] != ele[15][22];
    ele[15][17] != ele[15][23];
    ele[15][17] != ele[15][24];
    ele[15][17] != ele[16][15];
    ele[15][17] != ele[16][16];
    ele[15][17] != ele[16][17];
    ele[15][17] != ele[16][18];
    ele[15][17] != ele[16][19];
    ele[15][17] != ele[17][15];
    ele[15][17] != ele[17][16];
    ele[15][17] != ele[17][17];
    ele[15][17] != ele[17][18];
    ele[15][17] != ele[17][19];
    ele[15][17] != ele[18][15];
    ele[15][17] != ele[18][16];
    ele[15][17] != ele[18][17];
    ele[15][17] != ele[18][18];
    ele[15][17] != ele[18][19];
    ele[15][17] != ele[19][15];
    ele[15][17] != ele[19][16];
    ele[15][17] != ele[19][17];
    ele[15][17] != ele[19][18];
    ele[15][17] != ele[19][19];
    ele[15][17] != ele[20][17];
    ele[15][17] != ele[21][17];
    ele[15][17] != ele[22][17];
    ele[15][17] != ele[23][17];
    ele[15][17] != ele[24][17];
    ele[15][18] != ele[15][19];
    ele[15][18] != ele[15][20];
    ele[15][18] != ele[15][21];
    ele[15][18] != ele[15][22];
    ele[15][18] != ele[15][23];
    ele[15][18] != ele[15][24];
    ele[15][18] != ele[16][15];
    ele[15][18] != ele[16][16];
    ele[15][18] != ele[16][17];
    ele[15][18] != ele[16][18];
    ele[15][18] != ele[16][19];
    ele[15][18] != ele[17][15];
    ele[15][18] != ele[17][16];
    ele[15][18] != ele[17][17];
    ele[15][18] != ele[17][18];
    ele[15][18] != ele[17][19];
    ele[15][18] != ele[18][15];
    ele[15][18] != ele[18][16];
    ele[15][18] != ele[18][17];
    ele[15][18] != ele[18][18];
    ele[15][18] != ele[18][19];
    ele[15][18] != ele[19][15];
    ele[15][18] != ele[19][16];
    ele[15][18] != ele[19][17];
    ele[15][18] != ele[19][18];
    ele[15][18] != ele[19][19];
    ele[15][18] != ele[20][18];
    ele[15][18] != ele[21][18];
    ele[15][18] != ele[22][18];
    ele[15][18] != ele[23][18];
    ele[15][18] != ele[24][18];
    ele[15][19] != ele[15][20];
    ele[15][19] != ele[15][21];
    ele[15][19] != ele[15][22];
    ele[15][19] != ele[15][23];
    ele[15][19] != ele[15][24];
    ele[15][19] != ele[16][15];
    ele[15][19] != ele[16][16];
    ele[15][19] != ele[16][17];
    ele[15][19] != ele[16][18];
    ele[15][19] != ele[16][19];
    ele[15][19] != ele[17][15];
    ele[15][19] != ele[17][16];
    ele[15][19] != ele[17][17];
    ele[15][19] != ele[17][18];
    ele[15][19] != ele[17][19];
    ele[15][19] != ele[18][15];
    ele[15][19] != ele[18][16];
    ele[15][19] != ele[18][17];
    ele[15][19] != ele[18][18];
    ele[15][19] != ele[18][19];
    ele[15][19] != ele[19][15];
    ele[15][19] != ele[19][16];
    ele[15][19] != ele[19][17];
    ele[15][19] != ele[19][18];
    ele[15][19] != ele[19][19];
    ele[15][19] != ele[20][19];
    ele[15][19] != ele[21][19];
    ele[15][19] != ele[22][19];
    ele[15][19] != ele[23][19];
    ele[15][19] != ele[24][19];
    ele[15][2] != ele[15][10];
    ele[15][2] != ele[15][11];
    ele[15][2] != ele[15][12];
    ele[15][2] != ele[15][13];
    ele[15][2] != ele[15][14];
    ele[15][2] != ele[15][15];
    ele[15][2] != ele[15][16];
    ele[15][2] != ele[15][17];
    ele[15][2] != ele[15][18];
    ele[15][2] != ele[15][19];
    ele[15][2] != ele[15][20];
    ele[15][2] != ele[15][21];
    ele[15][2] != ele[15][22];
    ele[15][2] != ele[15][23];
    ele[15][2] != ele[15][24];
    ele[15][2] != ele[15][3];
    ele[15][2] != ele[15][4];
    ele[15][2] != ele[15][5];
    ele[15][2] != ele[15][6];
    ele[15][2] != ele[15][7];
    ele[15][2] != ele[15][8];
    ele[15][2] != ele[15][9];
    ele[15][2] != ele[16][0];
    ele[15][2] != ele[16][1];
    ele[15][2] != ele[16][2];
    ele[15][2] != ele[16][3];
    ele[15][2] != ele[16][4];
    ele[15][2] != ele[17][0];
    ele[15][2] != ele[17][1];
    ele[15][2] != ele[17][2];
    ele[15][2] != ele[17][3];
    ele[15][2] != ele[17][4];
    ele[15][2] != ele[18][0];
    ele[15][2] != ele[18][1];
    ele[15][2] != ele[18][2];
    ele[15][2] != ele[18][3];
    ele[15][2] != ele[18][4];
    ele[15][2] != ele[19][0];
    ele[15][2] != ele[19][1];
    ele[15][2] != ele[19][2];
    ele[15][2] != ele[19][3];
    ele[15][2] != ele[19][4];
    ele[15][2] != ele[20][2];
    ele[15][2] != ele[21][2];
    ele[15][2] != ele[22][2];
    ele[15][2] != ele[23][2];
    ele[15][2] != ele[24][2];
    ele[15][20] != ele[15][21];
    ele[15][20] != ele[15][22];
    ele[15][20] != ele[15][23];
    ele[15][20] != ele[15][24];
    ele[15][20] != ele[16][20];
    ele[15][20] != ele[16][21];
    ele[15][20] != ele[16][22];
    ele[15][20] != ele[16][23];
    ele[15][20] != ele[16][24];
    ele[15][20] != ele[17][20];
    ele[15][20] != ele[17][21];
    ele[15][20] != ele[17][22];
    ele[15][20] != ele[17][23];
    ele[15][20] != ele[17][24];
    ele[15][20] != ele[18][20];
    ele[15][20] != ele[18][21];
    ele[15][20] != ele[18][22];
    ele[15][20] != ele[18][23];
    ele[15][20] != ele[18][24];
    ele[15][20] != ele[19][20];
    ele[15][20] != ele[19][21];
    ele[15][20] != ele[19][22];
    ele[15][20] != ele[19][23];
    ele[15][20] != ele[19][24];
    ele[15][20] != ele[20][20];
    ele[15][20] != ele[21][20];
    ele[15][20] != ele[22][20];
    ele[15][20] != ele[23][20];
    ele[15][20] != ele[24][20];
    ele[15][21] != ele[15][22];
    ele[15][21] != ele[15][23];
    ele[15][21] != ele[15][24];
    ele[15][21] != ele[16][20];
    ele[15][21] != ele[16][21];
    ele[15][21] != ele[16][22];
    ele[15][21] != ele[16][23];
    ele[15][21] != ele[16][24];
    ele[15][21] != ele[17][20];
    ele[15][21] != ele[17][21];
    ele[15][21] != ele[17][22];
    ele[15][21] != ele[17][23];
    ele[15][21] != ele[17][24];
    ele[15][21] != ele[18][20];
    ele[15][21] != ele[18][21];
    ele[15][21] != ele[18][22];
    ele[15][21] != ele[18][23];
    ele[15][21] != ele[18][24];
    ele[15][21] != ele[19][20];
    ele[15][21] != ele[19][21];
    ele[15][21] != ele[19][22];
    ele[15][21] != ele[19][23];
    ele[15][21] != ele[19][24];
    ele[15][21] != ele[20][21];
    ele[15][21] != ele[21][21];
    ele[15][21] != ele[22][21];
    ele[15][21] != ele[23][21];
    ele[15][21] != ele[24][21];
    ele[15][22] != ele[15][23];
    ele[15][22] != ele[15][24];
    ele[15][22] != ele[16][20];
    ele[15][22] != ele[16][21];
    ele[15][22] != ele[16][22];
    ele[15][22] != ele[16][23];
    ele[15][22] != ele[16][24];
    ele[15][22] != ele[17][20];
    ele[15][22] != ele[17][21];
    ele[15][22] != ele[17][22];
    ele[15][22] != ele[17][23];
    ele[15][22] != ele[17][24];
    ele[15][22] != ele[18][20];
    ele[15][22] != ele[18][21];
    ele[15][22] != ele[18][22];
    ele[15][22] != ele[18][23];
    ele[15][22] != ele[18][24];
    ele[15][22] != ele[19][20];
    ele[15][22] != ele[19][21];
    ele[15][22] != ele[19][22];
    ele[15][22] != ele[19][23];
    ele[15][22] != ele[19][24];
    ele[15][22] != ele[20][22];
    ele[15][22] != ele[21][22];
    ele[15][22] != ele[22][22];
    ele[15][22] != ele[23][22];
    ele[15][22] != ele[24][22];
    ele[15][23] != ele[15][24];
    ele[15][23] != ele[16][20];
    ele[15][23] != ele[16][21];
    ele[15][23] != ele[16][22];
    ele[15][23] != ele[16][23];
    ele[15][23] != ele[16][24];
    ele[15][23] != ele[17][20];
    ele[15][23] != ele[17][21];
    ele[15][23] != ele[17][22];
    ele[15][23] != ele[17][23];
    ele[15][23] != ele[17][24];
    ele[15][23] != ele[18][20];
    ele[15][23] != ele[18][21];
    ele[15][23] != ele[18][22];
    ele[15][23] != ele[18][23];
    ele[15][23] != ele[18][24];
    ele[15][23] != ele[19][20];
    ele[15][23] != ele[19][21];
    ele[15][23] != ele[19][22];
    ele[15][23] != ele[19][23];
    ele[15][23] != ele[19][24];
    ele[15][23] != ele[20][23];
    ele[15][23] != ele[21][23];
    ele[15][23] != ele[22][23];
    ele[15][23] != ele[23][23];
    ele[15][23] != ele[24][23];
    ele[15][24] != ele[16][20];
    ele[15][24] != ele[16][21];
    ele[15][24] != ele[16][22];
    ele[15][24] != ele[16][23];
    ele[15][24] != ele[16][24];
    ele[15][24] != ele[17][20];
    ele[15][24] != ele[17][21];
    ele[15][24] != ele[17][22];
    ele[15][24] != ele[17][23];
    ele[15][24] != ele[17][24];
    ele[15][24] != ele[18][20];
    ele[15][24] != ele[18][21];
    ele[15][24] != ele[18][22];
    ele[15][24] != ele[18][23];
    ele[15][24] != ele[18][24];
    ele[15][24] != ele[19][20];
    ele[15][24] != ele[19][21];
    ele[15][24] != ele[19][22];
    ele[15][24] != ele[19][23];
    ele[15][24] != ele[19][24];
    ele[15][24] != ele[20][24];
    ele[15][24] != ele[21][24];
    ele[15][24] != ele[22][24];
    ele[15][24] != ele[23][24];
    ele[15][24] != ele[24][24];
    ele[15][3] != ele[15][10];
    ele[15][3] != ele[15][11];
    ele[15][3] != ele[15][12];
    ele[15][3] != ele[15][13];
    ele[15][3] != ele[15][14];
    ele[15][3] != ele[15][15];
    ele[15][3] != ele[15][16];
    ele[15][3] != ele[15][17];
    ele[15][3] != ele[15][18];
    ele[15][3] != ele[15][19];
    ele[15][3] != ele[15][20];
    ele[15][3] != ele[15][21];
    ele[15][3] != ele[15][22];
    ele[15][3] != ele[15][23];
    ele[15][3] != ele[15][24];
    ele[15][3] != ele[15][4];
    ele[15][3] != ele[15][5];
    ele[15][3] != ele[15][6];
    ele[15][3] != ele[15][7];
    ele[15][3] != ele[15][8];
    ele[15][3] != ele[15][9];
    ele[15][3] != ele[16][0];
    ele[15][3] != ele[16][1];
    ele[15][3] != ele[16][2];
    ele[15][3] != ele[16][3];
    ele[15][3] != ele[16][4];
    ele[15][3] != ele[17][0];
    ele[15][3] != ele[17][1];
    ele[15][3] != ele[17][2];
    ele[15][3] != ele[17][3];
    ele[15][3] != ele[17][4];
    ele[15][3] != ele[18][0];
    ele[15][3] != ele[18][1];
    ele[15][3] != ele[18][2];
    ele[15][3] != ele[18][3];
    ele[15][3] != ele[18][4];
    ele[15][3] != ele[19][0];
    ele[15][3] != ele[19][1];
    ele[15][3] != ele[19][2];
    ele[15][3] != ele[19][3];
    ele[15][3] != ele[19][4];
    ele[15][3] != ele[20][3];
    ele[15][3] != ele[21][3];
    ele[15][3] != ele[22][3];
    ele[15][3] != ele[23][3];
    ele[15][3] != ele[24][3];
    ele[15][4] != ele[15][10];
    ele[15][4] != ele[15][11];
    ele[15][4] != ele[15][12];
    ele[15][4] != ele[15][13];
    ele[15][4] != ele[15][14];
    ele[15][4] != ele[15][15];
    ele[15][4] != ele[15][16];
    ele[15][4] != ele[15][17];
    ele[15][4] != ele[15][18];
    ele[15][4] != ele[15][19];
    ele[15][4] != ele[15][20];
    ele[15][4] != ele[15][21];
    ele[15][4] != ele[15][22];
    ele[15][4] != ele[15][23];
    ele[15][4] != ele[15][24];
    ele[15][4] != ele[15][5];
    ele[15][4] != ele[15][6];
    ele[15][4] != ele[15][7];
    ele[15][4] != ele[15][8];
    ele[15][4] != ele[15][9];
    ele[15][4] != ele[16][0];
    ele[15][4] != ele[16][1];
    ele[15][4] != ele[16][2];
    ele[15][4] != ele[16][3];
    ele[15][4] != ele[16][4];
    ele[15][4] != ele[17][0];
    ele[15][4] != ele[17][1];
    ele[15][4] != ele[17][2];
    ele[15][4] != ele[17][3];
    ele[15][4] != ele[17][4];
    ele[15][4] != ele[18][0];
    ele[15][4] != ele[18][1];
    ele[15][4] != ele[18][2];
    ele[15][4] != ele[18][3];
    ele[15][4] != ele[18][4];
    ele[15][4] != ele[19][0];
    ele[15][4] != ele[19][1];
    ele[15][4] != ele[19][2];
    ele[15][4] != ele[19][3];
    ele[15][4] != ele[19][4];
    ele[15][4] != ele[20][4];
    ele[15][4] != ele[21][4];
    ele[15][4] != ele[22][4];
    ele[15][4] != ele[23][4];
    ele[15][4] != ele[24][4];
    ele[15][5] != ele[15][10];
    ele[15][5] != ele[15][11];
    ele[15][5] != ele[15][12];
    ele[15][5] != ele[15][13];
    ele[15][5] != ele[15][14];
    ele[15][5] != ele[15][15];
    ele[15][5] != ele[15][16];
    ele[15][5] != ele[15][17];
    ele[15][5] != ele[15][18];
    ele[15][5] != ele[15][19];
    ele[15][5] != ele[15][20];
    ele[15][5] != ele[15][21];
    ele[15][5] != ele[15][22];
    ele[15][5] != ele[15][23];
    ele[15][5] != ele[15][24];
    ele[15][5] != ele[15][6];
    ele[15][5] != ele[15][7];
    ele[15][5] != ele[15][8];
    ele[15][5] != ele[15][9];
    ele[15][5] != ele[16][5];
    ele[15][5] != ele[16][6];
    ele[15][5] != ele[16][7];
    ele[15][5] != ele[16][8];
    ele[15][5] != ele[16][9];
    ele[15][5] != ele[17][5];
    ele[15][5] != ele[17][6];
    ele[15][5] != ele[17][7];
    ele[15][5] != ele[17][8];
    ele[15][5] != ele[17][9];
    ele[15][5] != ele[18][5];
    ele[15][5] != ele[18][6];
    ele[15][5] != ele[18][7];
    ele[15][5] != ele[18][8];
    ele[15][5] != ele[18][9];
    ele[15][5] != ele[19][5];
    ele[15][5] != ele[19][6];
    ele[15][5] != ele[19][7];
    ele[15][5] != ele[19][8];
    ele[15][5] != ele[19][9];
    ele[15][5] != ele[20][5];
    ele[15][5] != ele[21][5];
    ele[15][5] != ele[22][5];
    ele[15][5] != ele[23][5];
    ele[15][5] != ele[24][5];
    ele[15][6] != ele[15][10];
    ele[15][6] != ele[15][11];
    ele[15][6] != ele[15][12];
    ele[15][6] != ele[15][13];
    ele[15][6] != ele[15][14];
    ele[15][6] != ele[15][15];
    ele[15][6] != ele[15][16];
    ele[15][6] != ele[15][17];
    ele[15][6] != ele[15][18];
    ele[15][6] != ele[15][19];
    ele[15][6] != ele[15][20];
    ele[15][6] != ele[15][21];
    ele[15][6] != ele[15][22];
    ele[15][6] != ele[15][23];
    ele[15][6] != ele[15][24];
    ele[15][6] != ele[15][7];
    ele[15][6] != ele[15][8];
    ele[15][6] != ele[15][9];
    ele[15][6] != ele[16][5];
    ele[15][6] != ele[16][6];
    ele[15][6] != ele[16][7];
    ele[15][6] != ele[16][8];
    ele[15][6] != ele[16][9];
    ele[15][6] != ele[17][5];
    ele[15][6] != ele[17][6];
    ele[15][6] != ele[17][7];
    ele[15][6] != ele[17][8];
    ele[15][6] != ele[17][9];
    ele[15][6] != ele[18][5];
    ele[15][6] != ele[18][6];
    ele[15][6] != ele[18][7];
    ele[15][6] != ele[18][8];
    ele[15][6] != ele[18][9];
    ele[15][6] != ele[19][5];
    ele[15][6] != ele[19][6];
    ele[15][6] != ele[19][7];
    ele[15][6] != ele[19][8];
    ele[15][6] != ele[19][9];
    ele[15][6] != ele[20][6];
    ele[15][6] != ele[21][6];
    ele[15][6] != ele[22][6];
    ele[15][6] != ele[23][6];
    ele[15][6] != ele[24][6];
    ele[15][7] != ele[15][10];
    ele[15][7] != ele[15][11];
    ele[15][7] != ele[15][12];
    ele[15][7] != ele[15][13];
    ele[15][7] != ele[15][14];
    ele[15][7] != ele[15][15];
    ele[15][7] != ele[15][16];
    ele[15][7] != ele[15][17];
    ele[15][7] != ele[15][18];
    ele[15][7] != ele[15][19];
    ele[15][7] != ele[15][20];
    ele[15][7] != ele[15][21];
    ele[15][7] != ele[15][22];
    ele[15][7] != ele[15][23];
    ele[15][7] != ele[15][24];
    ele[15][7] != ele[15][8];
    ele[15][7] != ele[15][9];
    ele[15][7] != ele[16][5];
    ele[15][7] != ele[16][6];
    ele[15][7] != ele[16][7];
    ele[15][7] != ele[16][8];
    ele[15][7] != ele[16][9];
    ele[15][7] != ele[17][5];
    ele[15][7] != ele[17][6];
    ele[15][7] != ele[17][7];
    ele[15][7] != ele[17][8];
    ele[15][7] != ele[17][9];
    ele[15][7] != ele[18][5];
    ele[15][7] != ele[18][6];
    ele[15][7] != ele[18][7];
    ele[15][7] != ele[18][8];
    ele[15][7] != ele[18][9];
    ele[15][7] != ele[19][5];
    ele[15][7] != ele[19][6];
    ele[15][7] != ele[19][7];
    ele[15][7] != ele[19][8];
    ele[15][7] != ele[19][9];
    ele[15][7] != ele[20][7];
    ele[15][7] != ele[21][7];
    ele[15][7] != ele[22][7];
    ele[15][7] != ele[23][7];
    ele[15][7] != ele[24][7];
    ele[15][8] != ele[15][10];
    ele[15][8] != ele[15][11];
    ele[15][8] != ele[15][12];
    ele[15][8] != ele[15][13];
    ele[15][8] != ele[15][14];
    ele[15][8] != ele[15][15];
    ele[15][8] != ele[15][16];
    ele[15][8] != ele[15][17];
    ele[15][8] != ele[15][18];
    ele[15][8] != ele[15][19];
    ele[15][8] != ele[15][20];
    ele[15][8] != ele[15][21];
    ele[15][8] != ele[15][22];
    ele[15][8] != ele[15][23];
    ele[15][8] != ele[15][24];
    ele[15][8] != ele[15][9];
    ele[15][8] != ele[16][5];
    ele[15][8] != ele[16][6];
    ele[15][8] != ele[16][7];
    ele[15][8] != ele[16][8];
    ele[15][8] != ele[16][9];
    ele[15][8] != ele[17][5];
    ele[15][8] != ele[17][6];
    ele[15][8] != ele[17][7];
    ele[15][8] != ele[17][8];
    ele[15][8] != ele[17][9];
    ele[15][8] != ele[18][5];
    ele[15][8] != ele[18][6];
    ele[15][8] != ele[18][7];
    ele[15][8] != ele[18][8];
    ele[15][8] != ele[18][9];
    ele[15][8] != ele[19][5];
    ele[15][8] != ele[19][6];
    ele[15][8] != ele[19][7];
    ele[15][8] != ele[19][8];
    ele[15][8] != ele[19][9];
    ele[15][8] != ele[20][8];
    ele[15][8] != ele[21][8];
    ele[15][8] != ele[22][8];
    ele[15][8] != ele[23][8];
    ele[15][8] != ele[24][8];
    ele[15][9] != ele[15][10];
    ele[15][9] != ele[15][11];
    ele[15][9] != ele[15][12];
    ele[15][9] != ele[15][13];
    ele[15][9] != ele[15][14];
    ele[15][9] != ele[15][15];
    ele[15][9] != ele[15][16];
    ele[15][9] != ele[15][17];
    ele[15][9] != ele[15][18];
    ele[15][9] != ele[15][19];
    ele[15][9] != ele[15][20];
    ele[15][9] != ele[15][21];
    ele[15][9] != ele[15][22];
    ele[15][9] != ele[15][23];
    ele[15][9] != ele[15][24];
    ele[15][9] != ele[16][5];
    ele[15][9] != ele[16][6];
    ele[15][9] != ele[16][7];
    ele[15][9] != ele[16][8];
    ele[15][9] != ele[16][9];
    ele[15][9] != ele[17][5];
    ele[15][9] != ele[17][6];
    ele[15][9] != ele[17][7];
    ele[15][9] != ele[17][8];
    ele[15][9] != ele[17][9];
    ele[15][9] != ele[18][5];
    ele[15][9] != ele[18][6];
    ele[15][9] != ele[18][7];
    ele[15][9] != ele[18][8];
    ele[15][9] != ele[18][9];
    ele[15][9] != ele[19][5];
    ele[15][9] != ele[19][6];
    ele[15][9] != ele[19][7];
    ele[15][9] != ele[19][8];
    ele[15][9] != ele[19][9];
    ele[15][9] != ele[20][9];
    ele[15][9] != ele[21][9];
    ele[15][9] != ele[22][9];
    ele[15][9] != ele[23][9];
    ele[15][9] != ele[24][9];
    ele[16][0] != ele[16][1];
    ele[16][0] != ele[16][10];
    ele[16][0] != ele[16][11];
    ele[16][0] != ele[16][12];
    ele[16][0] != ele[16][13];
    ele[16][0] != ele[16][14];
    ele[16][0] != ele[16][15];
    ele[16][0] != ele[16][16];
    ele[16][0] != ele[16][17];
    ele[16][0] != ele[16][18];
    ele[16][0] != ele[16][19];
    ele[16][0] != ele[16][2];
    ele[16][0] != ele[16][20];
    ele[16][0] != ele[16][21];
    ele[16][0] != ele[16][22];
    ele[16][0] != ele[16][23];
    ele[16][0] != ele[16][24];
    ele[16][0] != ele[16][3];
    ele[16][0] != ele[16][4];
    ele[16][0] != ele[16][5];
    ele[16][0] != ele[16][6];
    ele[16][0] != ele[16][7];
    ele[16][0] != ele[16][8];
    ele[16][0] != ele[16][9];
    ele[16][0] != ele[17][0];
    ele[16][0] != ele[17][1];
    ele[16][0] != ele[17][2];
    ele[16][0] != ele[17][3];
    ele[16][0] != ele[17][4];
    ele[16][0] != ele[18][0];
    ele[16][0] != ele[18][1];
    ele[16][0] != ele[18][2];
    ele[16][0] != ele[18][3];
    ele[16][0] != ele[18][4];
    ele[16][0] != ele[19][0];
    ele[16][0] != ele[19][1];
    ele[16][0] != ele[19][2];
    ele[16][0] != ele[19][3];
    ele[16][0] != ele[19][4];
    ele[16][0] != ele[20][0];
    ele[16][0] != ele[21][0];
    ele[16][0] != ele[22][0];
    ele[16][0] != ele[23][0];
    ele[16][0] != ele[24][0];
    ele[16][1] != ele[16][10];
    ele[16][1] != ele[16][11];
    ele[16][1] != ele[16][12];
    ele[16][1] != ele[16][13];
    ele[16][1] != ele[16][14];
    ele[16][1] != ele[16][15];
    ele[16][1] != ele[16][16];
    ele[16][1] != ele[16][17];
    ele[16][1] != ele[16][18];
    ele[16][1] != ele[16][19];
    ele[16][1] != ele[16][2];
    ele[16][1] != ele[16][20];
    ele[16][1] != ele[16][21];
    ele[16][1] != ele[16][22];
    ele[16][1] != ele[16][23];
    ele[16][1] != ele[16][24];
    ele[16][1] != ele[16][3];
    ele[16][1] != ele[16][4];
    ele[16][1] != ele[16][5];
    ele[16][1] != ele[16][6];
    ele[16][1] != ele[16][7];
    ele[16][1] != ele[16][8];
    ele[16][1] != ele[16][9];
    ele[16][1] != ele[17][0];
    ele[16][1] != ele[17][1];
    ele[16][1] != ele[17][2];
    ele[16][1] != ele[17][3];
    ele[16][1] != ele[17][4];
    ele[16][1] != ele[18][0];
    ele[16][1] != ele[18][1];
    ele[16][1] != ele[18][2];
    ele[16][1] != ele[18][3];
    ele[16][1] != ele[18][4];
    ele[16][1] != ele[19][0];
    ele[16][1] != ele[19][1];
    ele[16][1] != ele[19][2];
    ele[16][1] != ele[19][3];
    ele[16][1] != ele[19][4];
    ele[16][1] != ele[20][1];
    ele[16][1] != ele[21][1];
    ele[16][1] != ele[22][1];
    ele[16][1] != ele[23][1];
    ele[16][1] != ele[24][1];
    ele[16][10] != ele[16][11];
    ele[16][10] != ele[16][12];
    ele[16][10] != ele[16][13];
    ele[16][10] != ele[16][14];
    ele[16][10] != ele[16][15];
    ele[16][10] != ele[16][16];
    ele[16][10] != ele[16][17];
    ele[16][10] != ele[16][18];
    ele[16][10] != ele[16][19];
    ele[16][10] != ele[16][20];
    ele[16][10] != ele[16][21];
    ele[16][10] != ele[16][22];
    ele[16][10] != ele[16][23];
    ele[16][10] != ele[16][24];
    ele[16][10] != ele[17][10];
    ele[16][10] != ele[17][11];
    ele[16][10] != ele[17][12];
    ele[16][10] != ele[17][13];
    ele[16][10] != ele[17][14];
    ele[16][10] != ele[18][10];
    ele[16][10] != ele[18][11];
    ele[16][10] != ele[18][12];
    ele[16][10] != ele[18][13];
    ele[16][10] != ele[18][14];
    ele[16][10] != ele[19][10];
    ele[16][10] != ele[19][11];
    ele[16][10] != ele[19][12];
    ele[16][10] != ele[19][13];
    ele[16][10] != ele[19][14];
    ele[16][10] != ele[20][10];
    ele[16][10] != ele[21][10];
    ele[16][10] != ele[22][10];
    ele[16][10] != ele[23][10];
    ele[16][10] != ele[24][10];
    ele[16][11] != ele[16][12];
    ele[16][11] != ele[16][13];
    ele[16][11] != ele[16][14];
    ele[16][11] != ele[16][15];
    ele[16][11] != ele[16][16];
    ele[16][11] != ele[16][17];
    ele[16][11] != ele[16][18];
    ele[16][11] != ele[16][19];
    ele[16][11] != ele[16][20];
    ele[16][11] != ele[16][21];
    ele[16][11] != ele[16][22];
    ele[16][11] != ele[16][23];
    ele[16][11] != ele[16][24];
    ele[16][11] != ele[17][10];
    ele[16][11] != ele[17][11];
    ele[16][11] != ele[17][12];
    ele[16][11] != ele[17][13];
    ele[16][11] != ele[17][14];
    ele[16][11] != ele[18][10];
    ele[16][11] != ele[18][11];
    ele[16][11] != ele[18][12];
    ele[16][11] != ele[18][13];
    ele[16][11] != ele[18][14];
    ele[16][11] != ele[19][10];
    ele[16][11] != ele[19][11];
    ele[16][11] != ele[19][12];
    ele[16][11] != ele[19][13];
    ele[16][11] != ele[19][14];
    ele[16][11] != ele[20][11];
    ele[16][11] != ele[21][11];
    ele[16][11] != ele[22][11];
    ele[16][11] != ele[23][11];
    ele[16][11] != ele[24][11];
    ele[16][12] != ele[16][13];
    ele[16][12] != ele[16][14];
    ele[16][12] != ele[16][15];
    ele[16][12] != ele[16][16];
    ele[16][12] != ele[16][17];
    ele[16][12] != ele[16][18];
    ele[16][12] != ele[16][19];
    ele[16][12] != ele[16][20];
    ele[16][12] != ele[16][21];
    ele[16][12] != ele[16][22];
    ele[16][12] != ele[16][23];
    ele[16][12] != ele[16][24];
    ele[16][12] != ele[17][10];
    ele[16][12] != ele[17][11];
    ele[16][12] != ele[17][12];
    ele[16][12] != ele[17][13];
    ele[16][12] != ele[17][14];
    ele[16][12] != ele[18][10];
    ele[16][12] != ele[18][11];
    ele[16][12] != ele[18][12];
    ele[16][12] != ele[18][13];
    ele[16][12] != ele[18][14];
    ele[16][12] != ele[19][10];
    ele[16][12] != ele[19][11];
    ele[16][12] != ele[19][12];
    ele[16][12] != ele[19][13];
    ele[16][12] != ele[19][14];
    ele[16][12] != ele[20][12];
    ele[16][12] != ele[21][12];
    ele[16][12] != ele[22][12];
    ele[16][12] != ele[23][12];
    ele[16][12] != ele[24][12];
    ele[16][13] != ele[16][14];
    ele[16][13] != ele[16][15];
    ele[16][13] != ele[16][16];
    ele[16][13] != ele[16][17];
    ele[16][13] != ele[16][18];
    ele[16][13] != ele[16][19];
    ele[16][13] != ele[16][20];
    ele[16][13] != ele[16][21];
    ele[16][13] != ele[16][22];
    ele[16][13] != ele[16][23];
    ele[16][13] != ele[16][24];
    ele[16][13] != ele[17][10];
    ele[16][13] != ele[17][11];
    ele[16][13] != ele[17][12];
    ele[16][13] != ele[17][13];
    ele[16][13] != ele[17][14];
    ele[16][13] != ele[18][10];
    ele[16][13] != ele[18][11];
    ele[16][13] != ele[18][12];
    ele[16][13] != ele[18][13];
    ele[16][13] != ele[18][14];
    ele[16][13] != ele[19][10];
    ele[16][13] != ele[19][11];
    ele[16][13] != ele[19][12];
    ele[16][13] != ele[19][13];
    ele[16][13] != ele[19][14];
    ele[16][13] != ele[20][13];
    ele[16][13] != ele[21][13];
    ele[16][13] != ele[22][13];
    ele[16][13] != ele[23][13];
    ele[16][13] != ele[24][13];
    ele[16][14] != ele[16][15];
    ele[16][14] != ele[16][16];
    ele[16][14] != ele[16][17];
    ele[16][14] != ele[16][18];
    ele[16][14] != ele[16][19];
    ele[16][14] != ele[16][20];
    ele[16][14] != ele[16][21];
    ele[16][14] != ele[16][22];
    ele[16][14] != ele[16][23];
    ele[16][14] != ele[16][24];
    ele[16][14] != ele[17][10];
    ele[16][14] != ele[17][11];
    ele[16][14] != ele[17][12];
    ele[16][14] != ele[17][13];
    ele[16][14] != ele[17][14];
    ele[16][14] != ele[18][10];
    ele[16][14] != ele[18][11];
    ele[16][14] != ele[18][12];
    ele[16][14] != ele[18][13];
    ele[16][14] != ele[18][14];
    ele[16][14] != ele[19][10];
    ele[16][14] != ele[19][11];
    ele[16][14] != ele[19][12];
    ele[16][14] != ele[19][13];
    ele[16][14] != ele[19][14];
    ele[16][14] != ele[20][14];
    ele[16][14] != ele[21][14];
    ele[16][14] != ele[22][14];
    ele[16][14] != ele[23][14];
    ele[16][14] != ele[24][14];
    ele[16][15] != ele[16][16];
    ele[16][15] != ele[16][17];
    ele[16][15] != ele[16][18];
    ele[16][15] != ele[16][19];
    ele[16][15] != ele[16][20];
    ele[16][15] != ele[16][21];
    ele[16][15] != ele[16][22];
    ele[16][15] != ele[16][23];
    ele[16][15] != ele[16][24];
    ele[16][15] != ele[17][15];
    ele[16][15] != ele[17][16];
    ele[16][15] != ele[17][17];
    ele[16][15] != ele[17][18];
    ele[16][15] != ele[17][19];
    ele[16][15] != ele[18][15];
    ele[16][15] != ele[18][16];
    ele[16][15] != ele[18][17];
    ele[16][15] != ele[18][18];
    ele[16][15] != ele[18][19];
    ele[16][15] != ele[19][15];
    ele[16][15] != ele[19][16];
    ele[16][15] != ele[19][17];
    ele[16][15] != ele[19][18];
    ele[16][15] != ele[19][19];
    ele[16][15] != ele[20][15];
    ele[16][15] != ele[21][15];
    ele[16][15] != ele[22][15];
    ele[16][15] != ele[23][15];
    ele[16][15] != ele[24][15];
    ele[16][16] != ele[16][17];
    ele[16][16] != ele[16][18];
    ele[16][16] != ele[16][19];
    ele[16][16] != ele[16][20];
    ele[16][16] != ele[16][21];
    ele[16][16] != ele[16][22];
    ele[16][16] != ele[16][23];
    ele[16][16] != ele[16][24];
    ele[16][16] != ele[17][15];
    ele[16][16] != ele[17][16];
    ele[16][16] != ele[17][17];
    ele[16][16] != ele[17][18];
    ele[16][16] != ele[17][19];
    ele[16][16] != ele[18][15];
    ele[16][16] != ele[18][16];
    ele[16][16] != ele[18][17];
    ele[16][16] != ele[18][18];
    ele[16][16] != ele[18][19];
    ele[16][16] != ele[19][15];
    ele[16][16] != ele[19][16];
    ele[16][16] != ele[19][17];
    ele[16][16] != ele[19][18];
    ele[16][16] != ele[19][19];
    ele[16][16] != ele[20][16];
    ele[16][16] != ele[21][16];
    ele[16][16] != ele[22][16];
    ele[16][16] != ele[23][16];
    ele[16][16] != ele[24][16];
    ele[16][17] != ele[16][18];
    ele[16][17] != ele[16][19];
    ele[16][17] != ele[16][20];
    ele[16][17] != ele[16][21];
    ele[16][17] != ele[16][22];
    ele[16][17] != ele[16][23];
    ele[16][17] != ele[16][24];
    ele[16][17] != ele[17][15];
    ele[16][17] != ele[17][16];
    ele[16][17] != ele[17][17];
    ele[16][17] != ele[17][18];
    ele[16][17] != ele[17][19];
    ele[16][17] != ele[18][15];
    ele[16][17] != ele[18][16];
    ele[16][17] != ele[18][17];
    ele[16][17] != ele[18][18];
    ele[16][17] != ele[18][19];
    ele[16][17] != ele[19][15];
    ele[16][17] != ele[19][16];
    ele[16][17] != ele[19][17];
    ele[16][17] != ele[19][18];
    ele[16][17] != ele[19][19];
    ele[16][17] != ele[20][17];
    ele[16][17] != ele[21][17];
    ele[16][17] != ele[22][17];
    ele[16][17] != ele[23][17];
    ele[16][17] != ele[24][17];
    ele[16][18] != ele[16][19];
    ele[16][18] != ele[16][20];
    ele[16][18] != ele[16][21];
    ele[16][18] != ele[16][22];
    ele[16][18] != ele[16][23];
    ele[16][18] != ele[16][24];
    ele[16][18] != ele[17][15];
    ele[16][18] != ele[17][16];
    ele[16][18] != ele[17][17];
    ele[16][18] != ele[17][18];
    ele[16][18] != ele[17][19];
    ele[16][18] != ele[18][15];
    ele[16][18] != ele[18][16];
    ele[16][18] != ele[18][17];
    ele[16][18] != ele[18][18];
    ele[16][18] != ele[18][19];
    ele[16][18] != ele[19][15];
    ele[16][18] != ele[19][16];
    ele[16][18] != ele[19][17];
    ele[16][18] != ele[19][18];
    ele[16][18] != ele[19][19];
    ele[16][18] != ele[20][18];
    ele[16][18] != ele[21][18];
    ele[16][18] != ele[22][18];
    ele[16][18] != ele[23][18];
    ele[16][18] != ele[24][18];
    ele[16][19] != ele[16][20];
    ele[16][19] != ele[16][21];
    ele[16][19] != ele[16][22];
    ele[16][19] != ele[16][23];
    ele[16][19] != ele[16][24];
    ele[16][19] != ele[17][15];
    ele[16][19] != ele[17][16];
    ele[16][19] != ele[17][17];
    ele[16][19] != ele[17][18];
    ele[16][19] != ele[17][19];
    ele[16][19] != ele[18][15];
    ele[16][19] != ele[18][16];
    ele[16][19] != ele[18][17];
    ele[16][19] != ele[18][18];
    ele[16][19] != ele[18][19];
    ele[16][19] != ele[19][15];
    ele[16][19] != ele[19][16];
    ele[16][19] != ele[19][17];
    ele[16][19] != ele[19][18];
    ele[16][19] != ele[19][19];
    ele[16][19] != ele[20][19];
    ele[16][19] != ele[21][19];
    ele[16][19] != ele[22][19];
    ele[16][19] != ele[23][19];
    ele[16][19] != ele[24][19];
    ele[16][2] != ele[16][10];
    ele[16][2] != ele[16][11];
    ele[16][2] != ele[16][12];
    ele[16][2] != ele[16][13];
    ele[16][2] != ele[16][14];
    ele[16][2] != ele[16][15];
    ele[16][2] != ele[16][16];
    ele[16][2] != ele[16][17];
    ele[16][2] != ele[16][18];
    ele[16][2] != ele[16][19];
    ele[16][2] != ele[16][20];
    ele[16][2] != ele[16][21];
    ele[16][2] != ele[16][22];
    ele[16][2] != ele[16][23];
    ele[16][2] != ele[16][24];
    ele[16][2] != ele[16][3];
    ele[16][2] != ele[16][4];
    ele[16][2] != ele[16][5];
    ele[16][2] != ele[16][6];
    ele[16][2] != ele[16][7];
    ele[16][2] != ele[16][8];
    ele[16][2] != ele[16][9];
    ele[16][2] != ele[17][0];
    ele[16][2] != ele[17][1];
    ele[16][2] != ele[17][2];
    ele[16][2] != ele[17][3];
    ele[16][2] != ele[17][4];
    ele[16][2] != ele[18][0];
    ele[16][2] != ele[18][1];
    ele[16][2] != ele[18][2];
    ele[16][2] != ele[18][3];
    ele[16][2] != ele[18][4];
    ele[16][2] != ele[19][0];
    ele[16][2] != ele[19][1];
    ele[16][2] != ele[19][2];
    ele[16][2] != ele[19][3];
    ele[16][2] != ele[19][4];
    ele[16][2] != ele[20][2];
    ele[16][2] != ele[21][2];
    ele[16][2] != ele[22][2];
    ele[16][2] != ele[23][2];
    ele[16][2] != ele[24][2];
    ele[16][20] != ele[16][21];
    ele[16][20] != ele[16][22];
    ele[16][20] != ele[16][23];
    ele[16][20] != ele[16][24];
    ele[16][20] != ele[17][20];
    ele[16][20] != ele[17][21];
    ele[16][20] != ele[17][22];
    ele[16][20] != ele[17][23];
    ele[16][20] != ele[17][24];
    ele[16][20] != ele[18][20];
    ele[16][20] != ele[18][21];
    ele[16][20] != ele[18][22];
    ele[16][20] != ele[18][23];
    ele[16][20] != ele[18][24];
    ele[16][20] != ele[19][20];
    ele[16][20] != ele[19][21];
    ele[16][20] != ele[19][22];
    ele[16][20] != ele[19][23];
    ele[16][20] != ele[19][24];
    ele[16][20] != ele[20][20];
    ele[16][20] != ele[21][20];
    ele[16][20] != ele[22][20];
    ele[16][20] != ele[23][20];
    ele[16][20] != ele[24][20];
    ele[16][21] != ele[16][22];
    ele[16][21] != ele[16][23];
    ele[16][21] != ele[16][24];
    ele[16][21] != ele[17][20];
    ele[16][21] != ele[17][21];
    ele[16][21] != ele[17][22];
    ele[16][21] != ele[17][23];
    ele[16][21] != ele[17][24];
    ele[16][21] != ele[18][20];
    ele[16][21] != ele[18][21];
    ele[16][21] != ele[18][22];
    ele[16][21] != ele[18][23];
    ele[16][21] != ele[18][24];
    ele[16][21] != ele[19][20];
    ele[16][21] != ele[19][21];
    ele[16][21] != ele[19][22];
    ele[16][21] != ele[19][23];
    ele[16][21] != ele[19][24];
    ele[16][21] != ele[20][21];
    ele[16][21] != ele[21][21];
    ele[16][21] != ele[22][21];
    ele[16][21] != ele[23][21];
    ele[16][21] != ele[24][21];
    ele[16][22] != ele[16][23];
    ele[16][22] != ele[16][24];
    ele[16][22] != ele[17][20];
    ele[16][22] != ele[17][21];
    ele[16][22] != ele[17][22];
    ele[16][22] != ele[17][23];
    ele[16][22] != ele[17][24];
    ele[16][22] != ele[18][20];
    ele[16][22] != ele[18][21];
    ele[16][22] != ele[18][22];
    ele[16][22] != ele[18][23];
    ele[16][22] != ele[18][24];
    ele[16][22] != ele[19][20];
    ele[16][22] != ele[19][21];
    ele[16][22] != ele[19][22];
    ele[16][22] != ele[19][23];
    ele[16][22] != ele[19][24];
    ele[16][22] != ele[20][22];
    ele[16][22] != ele[21][22];
    ele[16][22] != ele[22][22];
    ele[16][22] != ele[23][22];
    ele[16][22] != ele[24][22];
    ele[16][23] != ele[16][24];
    ele[16][23] != ele[17][20];
    ele[16][23] != ele[17][21];
    ele[16][23] != ele[17][22];
    ele[16][23] != ele[17][23];
    ele[16][23] != ele[17][24];
    ele[16][23] != ele[18][20];
    ele[16][23] != ele[18][21];
    ele[16][23] != ele[18][22];
    ele[16][23] != ele[18][23];
    ele[16][23] != ele[18][24];
    ele[16][23] != ele[19][20];
    ele[16][23] != ele[19][21];
    ele[16][23] != ele[19][22];
    ele[16][23] != ele[19][23];
    ele[16][23] != ele[19][24];
    ele[16][23] != ele[20][23];
    ele[16][23] != ele[21][23];
    ele[16][23] != ele[22][23];
    ele[16][23] != ele[23][23];
    ele[16][23] != ele[24][23];
    ele[16][24] != ele[17][20];
    ele[16][24] != ele[17][21];
    ele[16][24] != ele[17][22];
    ele[16][24] != ele[17][23];
    ele[16][24] != ele[17][24];
    ele[16][24] != ele[18][20];
    ele[16][24] != ele[18][21];
    ele[16][24] != ele[18][22];
    ele[16][24] != ele[18][23];
    ele[16][24] != ele[18][24];
    ele[16][24] != ele[19][20];
    ele[16][24] != ele[19][21];
    ele[16][24] != ele[19][22];
    ele[16][24] != ele[19][23];
    ele[16][24] != ele[19][24];
    ele[16][24] != ele[20][24];
    ele[16][24] != ele[21][24];
    ele[16][24] != ele[22][24];
    ele[16][24] != ele[23][24];
    ele[16][24] != ele[24][24];
    ele[16][3] != ele[16][10];
    ele[16][3] != ele[16][11];
    ele[16][3] != ele[16][12];
    ele[16][3] != ele[16][13];
    ele[16][3] != ele[16][14];
    ele[16][3] != ele[16][15];
    ele[16][3] != ele[16][16];
    ele[16][3] != ele[16][17];
    ele[16][3] != ele[16][18];
    ele[16][3] != ele[16][19];
    ele[16][3] != ele[16][20];
    ele[16][3] != ele[16][21];
    ele[16][3] != ele[16][22];
    ele[16][3] != ele[16][23];
    ele[16][3] != ele[16][24];
    ele[16][3] != ele[16][4];
    ele[16][3] != ele[16][5];
    ele[16][3] != ele[16][6];
    ele[16][3] != ele[16][7];
    ele[16][3] != ele[16][8];
    ele[16][3] != ele[16][9];
    ele[16][3] != ele[17][0];
    ele[16][3] != ele[17][1];
    ele[16][3] != ele[17][2];
    ele[16][3] != ele[17][3];
    ele[16][3] != ele[17][4];
    ele[16][3] != ele[18][0];
    ele[16][3] != ele[18][1];
    ele[16][3] != ele[18][2];
    ele[16][3] != ele[18][3];
    ele[16][3] != ele[18][4];
    ele[16][3] != ele[19][0];
    ele[16][3] != ele[19][1];
    ele[16][3] != ele[19][2];
    ele[16][3] != ele[19][3];
    ele[16][3] != ele[19][4];
    ele[16][3] != ele[20][3];
    ele[16][3] != ele[21][3];
    ele[16][3] != ele[22][3];
    ele[16][3] != ele[23][3];
    ele[16][3] != ele[24][3];
    ele[16][4] != ele[16][10];
    ele[16][4] != ele[16][11];
    ele[16][4] != ele[16][12];
    ele[16][4] != ele[16][13];
    ele[16][4] != ele[16][14];
    ele[16][4] != ele[16][15];
    ele[16][4] != ele[16][16];
    ele[16][4] != ele[16][17];
    ele[16][4] != ele[16][18];
    ele[16][4] != ele[16][19];
    ele[16][4] != ele[16][20];
    ele[16][4] != ele[16][21];
    ele[16][4] != ele[16][22];
    ele[16][4] != ele[16][23];
    ele[16][4] != ele[16][24];
    ele[16][4] != ele[16][5];
    ele[16][4] != ele[16][6];
    ele[16][4] != ele[16][7];
    ele[16][4] != ele[16][8];
    ele[16][4] != ele[16][9];
    ele[16][4] != ele[17][0];
    ele[16][4] != ele[17][1];
    ele[16][4] != ele[17][2];
    ele[16][4] != ele[17][3];
    ele[16][4] != ele[17][4];
    ele[16][4] != ele[18][0];
    ele[16][4] != ele[18][1];
    ele[16][4] != ele[18][2];
    ele[16][4] != ele[18][3];
    ele[16][4] != ele[18][4];
    ele[16][4] != ele[19][0];
    ele[16][4] != ele[19][1];
    ele[16][4] != ele[19][2];
    ele[16][4] != ele[19][3];
    ele[16][4] != ele[19][4];
    ele[16][4] != ele[20][4];
    ele[16][4] != ele[21][4];
    ele[16][4] != ele[22][4];
    ele[16][4] != ele[23][4];
    ele[16][4] != ele[24][4];
    ele[16][5] != ele[16][10];
    ele[16][5] != ele[16][11];
    ele[16][5] != ele[16][12];
    ele[16][5] != ele[16][13];
    ele[16][5] != ele[16][14];
    ele[16][5] != ele[16][15];
    ele[16][5] != ele[16][16];
    ele[16][5] != ele[16][17];
    ele[16][5] != ele[16][18];
    ele[16][5] != ele[16][19];
    ele[16][5] != ele[16][20];
    ele[16][5] != ele[16][21];
    ele[16][5] != ele[16][22];
    ele[16][5] != ele[16][23];
    ele[16][5] != ele[16][24];
    ele[16][5] != ele[16][6];
    ele[16][5] != ele[16][7];
    ele[16][5] != ele[16][8];
    ele[16][5] != ele[16][9];
    ele[16][5] != ele[17][5];
    ele[16][5] != ele[17][6];
    ele[16][5] != ele[17][7];
    ele[16][5] != ele[17][8];
    ele[16][5] != ele[17][9];
    ele[16][5] != ele[18][5];
    ele[16][5] != ele[18][6];
    ele[16][5] != ele[18][7];
    ele[16][5] != ele[18][8];
    ele[16][5] != ele[18][9];
    ele[16][5] != ele[19][5];
    ele[16][5] != ele[19][6];
    ele[16][5] != ele[19][7];
    ele[16][5] != ele[19][8];
    ele[16][5] != ele[19][9];
    ele[16][5] != ele[20][5];
    ele[16][5] != ele[21][5];
    ele[16][5] != ele[22][5];
    ele[16][5] != ele[23][5];
    ele[16][5] != ele[24][5];
    ele[16][6] != ele[16][10];
    ele[16][6] != ele[16][11];
    ele[16][6] != ele[16][12];
    ele[16][6] != ele[16][13];
    ele[16][6] != ele[16][14];
    ele[16][6] != ele[16][15];
    ele[16][6] != ele[16][16];
    ele[16][6] != ele[16][17];
    ele[16][6] != ele[16][18];
    ele[16][6] != ele[16][19];
    ele[16][6] != ele[16][20];
    ele[16][6] != ele[16][21];
    ele[16][6] != ele[16][22];
    ele[16][6] != ele[16][23];
    ele[16][6] != ele[16][24];
    ele[16][6] != ele[16][7];
    ele[16][6] != ele[16][8];
    ele[16][6] != ele[16][9];
    ele[16][6] != ele[17][5];
    ele[16][6] != ele[17][6];
    ele[16][6] != ele[17][7];
    ele[16][6] != ele[17][8];
    ele[16][6] != ele[17][9];
    ele[16][6] != ele[18][5];
    ele[16][6] != ele[18][6];
    ele[16][6] != ele[18][7];
    ele[16][6] != ele[18][8];
    ele[16][6] != ele[18][9];
    ele[16][6] != ele[19][5];
    ele[16][6] != ele[19][6];
    ele[16][6] != ele[19][7];
    ele[16][6] != ele[19][8];
    ele[16][6] != ele[19][9];
    ele[16][6] != ele[20][6];
    ele[16][6] != ele[21][6];
    ele[16][6] != ele[22][6];
    ele[16][6] != ele[23][6];
    ele[16][6] != ele[24][6];
    ele[16][7] != ele[16][10];
    ele[16][7] != ele[16][11];
    ele[16][7] != ele[16][12];
    ele[16][7] != ele[16][13];
    ele[16][7] != ele[16][14];
    ele[16][7] != ele[16][15];
    ele[16][7] != ele[16][16];
    ele[16][7] != ele[16][17];
    ele[16][7] != ele[16][18];
    ele[16][7] != ele[16][19];
    ele[16][7] != ele[16][20];
    ele[16][7] != ele[16][21];
    ele[16][7] != ele[16][22];
    ele[16][7] != ele[16][23];
    ele[16][7] != ele[16][24];
    ele[16][7] != ele[16][8];
    ele[16][7] != ele[16][9];
    ele[16][7] != ele[17][5];
    ele[16][7] != ele[17][6];
    ele[16][7] != ele[17][7];
    ele[16][7] != ele[17][8];
    ele[16][7] != ele[17][9];
    ele[16][7] != ele[18][5];
    ele[16][7] != ele[18][6];
    ele[16][7] != ele[18][7];
    ele[16][7] != ele[18][8];
    ele[16][7] != ele[18][9];
    ele[16][7] != ele[19][5];
    ele[16][7] != ele[19][6];
    ele[16][7] != ele[19][7];
    ele[16][7] != ele[19][8];
    ele[16][7] != ele[19][9];
    ele[16][7] != ele[20][7];
    ele[16][7] != ele[21][7];
    ele[16][7] != ele[22][7];
    ele[16][7] != ele[23][7];
    ele[16][7] != ele[24][7];
    ele[16][8] != ele[16][10];
    ele[16][8] != ele[16][11];
    ele[16][8] != ele[16][12];
    ele[16][8] != ele[16][13];
    ele[16][8] != ele[16][14];
    ele[16][8] != ele[16][15];
    ele[16][8] != ele[16][16];
    ele[16][8] != ele[16][17];
    ele[16][8] != ele[16][18];
    ele[16][8] != ele[16][19];
    ele[16][8] != ele[16][20];
    ele[16][8] != ele[16][21];
    ele[16][8] != ele[16][22];
    ele[16][8] != ele[16][23];
    ele[16][8] != ele[16][24];
    ele[16][8] != ele[16][9];
    ele[16][8] != ele[17][5];
    ele[16][8] != ele[17][6];
    ele[16][8] != ele[17][7];
    ele[16][8] != ele[17][8];
    ele[16][8] != ele[17][9];
    ele[16][8] != ele[18][5];
    ele[16][8] != ele[18][6];
    ele[16][8] != ele[18][7];
    ele[16][8] != ele[18][8];
    ele[16][8] != ele[18][9];
    ele[16][8] != ele[19][5];
    ele[16][8] != ele[19][6];
    ele[16][8] != ele[19][7];
    ele[16][8] != ele[19][8];
    ele[16][8] != ele[19][9];
    ele[16][8] != ele[20][8];
    ele[16][8] != ele[21][8];
    ele[16][8] != ele[22][8];
    ele[16][8] != ele[23][8];
    ele[16][8] != ele[24][8];
    ele[16][9] != ele[16][10];
    ele[16][9] != ele[16][11];
    ele[16][9] != ele[16][12];
    ele[16][9] != ele[16][13];
    ele[16][9] != ele[16][14];
    ele[16][9] != ele[16][15];
    ele[16][9] != ele[16][16];
    ele[16][9] != ele[16][17];
    ele[16][9] != ele[16][18];
    ele[16][9] != ele[16][19];
    ele[16][9] != ele[16][20];
    ele[16][9] != ele[16][21];
    ele[16][9] != ele[16][22];
    ele[16][9] != ele[16][23];
    ele[16][9] != ele[16][24];
    ele[16][9] != ele[17][5];
    ele[16][9] != ele[17][6];
    ele[16][9] != ele[17][7];
    ele[16][9] != ele[17][8];
    ele[16][9] != ele[17][9];
    ele[16][9] != ele[18][5];
    ele[16][9] != ele[18][6];
    ele[16][9] != ele[18][7];
    ele[16][9] != ele[18][8];
    ele[16][9] != ele[18][9];
    ele[16][9] != ele[19][5];
    ele[16][9] != ele[19][6];
    ele[16][9] != ele[19][7];
    ele[16][9] != ele[19][8];
    ele[16][9] != ele[19][9];
    ele[16][9] != ele[20][9];
    ele[16][9] != ele[21][9];
    ele[16][9] != ele[22][9];
    ele[16][9] != ele[23][9];
    ele[16][9] != ele[24][9];
    ele[17][0] != ele[17][1];
    ele[17][0] != ele[17][10];
    ele[17][0] != ele[17][11];
    ele[17][0] != ele[17][12];
    ele[17][0] != ele[17][13];
    ele[17][0] != ele[17][14];
    ele[17][0] != ele[17][15];
    ele[17][0] != ele[17][16];
    ele[17][0] != ele[17][17];
    ele[17][0] != ele[17][18];
    ele[17][0] != ele[17][19];
    ele[17][0] != ele[17][2];
    ele[17][0] != ele[17][20];
    ele[17][0] != ele[17][21];
    ele[17][0] != ele[17][22];
    ele[17][0] != ele[17][23];
    ele[17][0] != ele[17][24];
    ele[17][0] != ele[17][3];
    ele[17][0] != ele[17][4];
    ele[17][0] != ele[17][5];
    ele[17][0] != ele[17][6];
    ele[17][0] != ele[17][7];
    ele[17][0] != ele[17][8];
    ele[17][0] != ele[17][9];
    ele[17][0] != ele[18][0];
    ele[17][0] != ele[18][1];
    ele[17][0] != ele[18][2];
    ele[17][0] != ele[18][3];
    ele[17][0] != ele[18][4];
    ele[17][0] != ele[19][0];
    ele[17][0] != ele[19][1];
    ele[17][0] != ele[19][2];
    ele[17][0] != ele[19][3];
    ele[17][0] != ele[19][4];
    ele[17][0] != ele[20][0];
    ele[17][0] != ele[21][0];
    ele[17][0] != ele[22][0];
    ele[17][0] != ele[23][0];
    ele[17][0] != ele[24][0];
    ele[17][1] != ele[17][10];
    ele[17][1] != ele[17][11];
    ele[17][1] != ele[17][12];
    ele[17][1] != ele[17][13];
    ele[17][1] != ele[17][14];
    ele[17][1] != ele[17][15];
    ele[17][1] != ele[17][16];
    ele[17][1] != ele[17][17];
    ele[17][1] != ele[17][18];
    ele[17][1] != ele[17][19];
    ele[17][1] != ele[17][2];
    ele[17][1] != ele[17][20];
    ele[17][1] != ele[17][21];
    ele[17][1] != ele[17][22];
    ele[17][1] != ele[17][23];
    ele[17][1] != ele[17][24];
    ele[17][1] != ele[17][3];
    ele[17][1] != ele[17][4];
    ele[17][1] != ele[17][5];
    ele[17][1] != ele[17][6];
    ele[17][1] != ele[17][7];
    ele[17][1] != ele[17][8];
    ele[17][1] != ele[17][9];
    ele[17][1] != ele[18][0];
    ele[17][1] != ele[18][1];
    ele[17][1] != ele[18][2];
    ele[17][1] != ele[18][3];
    ele[17][1] != ele[18][4];
    ele[17][1] != ele[19][0];
    ele[17][1] != ele[19][1];
    ele[17][1] != ele[19][2];
    ele[17][1] != ele[19][3];
    ele[17][1] != ele[19][4];
    ele[17][1] != ele[20][1];
    ele[17][1] != ele[21][1];
    ele[17][1] != ele[22][1];
    ele[17][1] != ele[23][1];
    ele[17][1] != ele[24][1];
    ele[17][10] != ele[17][11];
    ele[17][10] != ele[17][12];
    ele[17][10] != ele[17][13];
    ele[17][10] != ele[17][14];
    ele[17][10] != ele[17][15];
    ele[17][10] != ele[17][16];
    ele[17][10] != ele[17][17];
    ele[17][10] != ele[17][18];
    ele[17][10] != ele[17][19];
    ele[17][10] != ele[17][20];
    ele[17][10] != ele[17][21];
    ele[17][10] != ele[17][22];
    ele[17][10] != ele[17][23];
    ele[17][10] != ele[17][24];
    ele[17][10] != ele[18][10];
    ele[17][10] != ele[18][11];
    ele[17][10] != ele[18][12];
    ele[17][10] != ele[18][13];
    ele[17][10] != ele[18][14];
    ele[17][10] != ele[19][10];
    ele[17][10] != ele[19][11];
    ele[17][10] != ele[19][12];
    ele[17][10] != ele[19][13];
    ele[17][10] != ele[19][14];
    ele[17][10] != ele[20][10];
    ele[17][10] != ele[21][10];
    ele[17][10] != ele[22][10];
    ele[17][10] != ele[23][10];
    ele[17][10] != ele[24][10];
    ele[17][11] != ele[17][12];
    ele[17][11] != ele[17][13];
    ele[17][11] != ele[17][14];
    ele[17][11] != ele[17][15];
    ele[17][11] != ele[17][16];
    ele[17][11] != ele[17][17];
    ele[17][11] != ele[17][18];
    ele[17][11] != ele[17][19];
    ele[17][11] != ele[17][20];
    ele[17][11] != ele[17][21];
    ele[17][11] != ele[17][22];
    ele[17][11] != ele[17][23];
    ele[17][11] != ele[17][24];
    ele[17][11] != ele[18][10];
    ele[17][11] != ele[18][11];
    ele[17][11] != ele[18][12];
    ele[17][11] != ele[18][13];
    ele[17][11] != ele[18][14];
    ele[17][11] != ele[19][10];
    ele[17][11] != ele[19][11];
    ele[17][11] != ele[19][12];
    ele[17][11] != ele[19][13];
    ele[17][11] != ele[19][14];
    ele[17][11] != ele[20][11];
    ele[17][11] != ele[21][11];
    ele[17][11] != ele[22][11];
    ele[17][11] != ele[23][11];
    ele[17][11] != ele[24][11];
    ele[17][12] != ele[17][13];
    ele[17][12] != ele[17][14];
    ele[17][12] != ele[17][15];
    ele[17][12] != ele[17][16];
    ele[17][12] != ele[17][17];
    ele[17][12] != ele[17][18];
    ele[17][12] != ele[17][19];
    ele[17][12] != ele[17][20];
    ele[17][12] != ele[17][21];
    ele[17][12] != ele[17][22];
    ele[17][12] != ele[17][23];
    ele[17][12] != ele[17][24];
    ele[17][12] != ele[18][10];
    ele[17][12] != ele[18][11];
    ele[17][12] != ele[18][12];
    ele[17][12] != ele[18][13];
    ele[17][12] != ele[18][14];
    ele[17][12] != ele[19][10];
    ele[17][12] != ele[19][11];
    ele[17][12] != ele[19][12];
    ele[17][12] != ele[19][13];
    ele[17][12] != ele[19][14];
    ele[17][12] != ele[20][12];
    ele[17][12] != ele[21][12];
    ele[17][12] != ele[22][12];
    ele[17][12] != ele[23][12];
    ele[17][12] != ele[24][12];
    ele[17][13] != ele[17][14];
    ele[17][13] != ele[17][15];
    ele[17][13] != ele[17][16];
    ele[17][13] != ele[17][17];
    ele[17][13] != ele[17][18];
    ele[17][13] != ele[17][19];
    ele[17][13] != ele[17][20];
    ele[17][13] != ele[17][21];
    ele[17][13] != ele[17][22];
    ele[17][13] != ele[17][23];
    ele[17][13] != ele[17][24];
    ele[17][13] != ele[18][10];
    ele[17][13] != ele[18][11];
    ele[17][13] != ele[18][12];
    ele[17][13] != ele[18][13];
    ele[17][13] != ele[18][14];
    ele[17][13] != ele[19][10];
    ele[17][13] != ele[19][11];
    ele[17][13] != ele[19][12];
    ele[17][13] != ele[19][13];
    ele[17][13] != ele[19][14];
    ele[17][13] != ele[20][13];
    ele[17][13] != ele[21][13];
    ele[17][13] != ele[22][13];
    ele[17][13] != ele[23][13];
    ele[17][13] != ele[24][13];
    ele[17][14] != ele[17][15];
    ele[17][14] != ele[17][16];
    ele[17][14] != ele[17][17];
    ele[17][14] != ele[17][18];
    ele[17][14] != ele[17][19];
    ele[17][14] != ele[17][20];
    ele[17][14] != ele[17][21];
    ele[17][14] != ele[17][22];
    ele[17][14] != ele[17][23];
    ele[17][14] != ele[17][24];
    ele[17][14] != ele[18][10];
    ele[17][14] != ele[18][11];
    ele[17][14] != ele[18][12];
    ele[17][14] != ele[18][13];
    ele[17][14] != ele[18][14];
    ele[17][14] != ele[19][10];
    ele[17][14] != ele[19][11];
    ele[17][14] != ele[19][12];
    ele[17][14] != ele[19][13];
    ele[17][14] != ele[19][14];
    ele[17][14] != ele[20][14];
    ele[17][14] != ele[21][14];
    ele[17][14] != ele[22][14];
    ele[17][14] != ele[23][14];
    ele[17][14] != ele[24][14];
    ele[17][15] != ele[17][16];
    ele[17][15] != ele[17][17];
    ele[17][15] != ele[17][18];
    ele[17][15] != ele[17][19];
    ele[17][15] != ele[17][20];
    ele[17][15] != ele[17][21];
    ele[17][15] != ele[17][22];
    ele[17][15] != ele[17][23];
    ele[17][15] != ele[17][24];
    ele[17][15] != ele[18][15];
    ele[17][15] != ele[18][16];
    ele[17][15] != ele[18][17];
    ele[17][15] != ele[18][18];
    ele[17][15] != ele[18][19];
    ele[17][15] != ele[19][15];
    ele[17][15] != ele[19][16];
    ele[17][15] != ele[19][17];
    ele[17][15] != ele[19][18];
    ele[17][15] != ele[19][19];
    ele[17][15] != ele[20][15];
    ele[17][15] != ele[21][15];
    ele[17][15] != ele[22][15];
    ele[17][15] != ele[23][15];
    ele[17][15] != ele[24][15];
    ele[17][16] != ele[17][17];
    ele[17][16] != ele[17][18];
    ele[17][16] != ele[17][19];
    ele[17][16] != ele[17][20];
    ele[17][16] != ele[17][21];
    ele[17][16] != ele[17][22];
    ele[17][16] != ele[17][23];
    ele[17][16] != ele[17][24];
    ele[17][16] != ele[18][15];
    ele[17][16] != ele[18][16];
    ele[17][16] != ele[18][17];
    ele[17][16] != ele[18][18];
    ele[17][16] != ele[18][19];
    ele[17][16] != ele[19][15];
    ele[17][16] != ele[19][16];
    ele[17][16] != ele[19][17];
    ele[17][16] != ele[19][18];
    ele[17][16] != ele[19][19];
    ele[17][16] != ele[20][16];
    ele[17][16] != ele[21][16];
    ele[17][16] != ele[22][16];
    ele[17][16] != ele[23][16];
    ele[17][16] != ele[24][16];
    ele[17][17] != ele[17][18];
    ele[17][17] != ele[17][19];
    ele[17][17] != ele[17][20];
    ele[17][17] != ele[17][21];
    ele[17][17] != ele[17][22];
    ele[17][17] != ele[17][23];
    ele[17][17] != ele[17][24];
    ele[17][17] != ele[18][15];
    ele[17][17] != ele[18][16];
    ele[17][17] != ele[18][17];
    ele[17][17] != ele[18][18];
    ele[17][17] != ele[18][19];
    ele[17][17] != ele[19][15];
    ele[17][17] != ele[19][16];
    ele[17][17] != ele[19][17];
    ele[17][17] != ele[19][18];
    ele[17][17] != ele[19][19];
    ele[17][17] != ele[20][17];
    ele[17][17] != ele[21][17];
    ele[17][17] != ele[22][17];
    ele[17][17] != ele[23][17];
    ele[17][17] != ele[24][17];
    ele[17][18] != ele[17][19];
    ele[17][18] != ele[17][20];
    ele[17][18] != ele[17][21];
    ele[17][18] != ele[17][22];
    ele[17][18] != ele[17][23];
    ele[17][18] != ele[17][24];
    ele[17][18] != ele[18][15];
    ele[17][18] != ele[18][16];
    ele[17][18] != ele[18][17];
    ele[17][18] != ele[18][18];
    ele[17][18] != ele[18][19];
    ele[17][18] != ele[19][15];
    ele[17][18] != ele[19][16];
    ele[17][18] != ele[19][17];
    ele[17][18] != ele[19][18];
    ele[17][18] != ele[19][19];
    ele[17][18] != ele[20][18];
    ele[17][18] != ele[21][18];
    ele[17][18] != ele[22][18];
    ele[17][18] != ele[23][18];
    ele[17][18] != ele[24][18];
    ele[17][19] != ele[17][20];
    ele[17][19] != ele[17][21];
    ele[17][19] != ele[17][22];
    ele[17][19] != ele[17][23];
    ele[17][19] != ele[17][24];
    ele[17][19] != ele[18][15];
    ele[17][19] != ele[18][16];
    ele[17][19] != ele[18][17];
    ele[17][19] != ele[18][18];
    ele[17][19] != ele[18][19];
    ele[17][19] != ele[19][15];
    ele[17][19] != ele[19][16];
    ele[17][19] != ele[19][17];
    ele[17][19] != ele[19][18];
    ele[17][19] != ele[19][19];
    ele[17][19] != ele[20][19];
    ele[17][19] != ele[21][19];
    ele[17][19] != ele[22][19];
    ele[17][19] != ele[23][19];
    ele[17][19] != ele[24][19];
    ele[17][2] != ele[17][10];
    ele[17][2] != ele[17][11];
    ele[17][2] != ele[17][12];
    ele[17][2] != ele[17][13];
    ele[17][2] != ele[17][14];
    ele[17][2] != ele[17][15];
    ele[17][2] != ele[17][16];
    ele[17][2] != ele[17][17];
    ele[17][2] != ele[17][18];
    ele[17][2] != ele[17][19];
    ele[17][2] != ele[17][20];
    ele[17][2] != ele[17][21];
    ele[17][2] != ele[17][22];
    ele[17][2] != ele[17][23];
    ele[17][2] != ele[17][24];
    ele[17][2] != ele[17][3];
    ele[17][2] != ele[17][4];
    ele[17][2] != ele[17][5];
    ele[17][2] != ele[17][6];
    ele[17][2] != ele[17][7];
    ele[17][2] != ele[17][8];
    ele[17][2] != ele[17][9];
    ele[17][2] != ele[18][0];
    ele[17][2] != ele[18][1];
    ele[17][2] != ele[18][2];
    ele[17][2] != ele[18][3];
    ele[17][2] != ele[18][4];
    ele[17][2] != ele[19][0];
    ele[17][2] != ele[19][1];
    ele[17][2] != ele[19][2];
    ele[17][2] != ele[19][3];
    ele[17][2] != ele[19][4];
    ele[17][2] != ele[20][2];
    ele[17][2] != ele[21][2];
    ele[17][2] != ele[22][2];
    ele[17][2] != ele[23][2];
    ele[17][2] != ele[24][2];
    ele[17][20] != ele[17][21];
    ele[17][20] != ele[17][22];
    ele[17][20] != ele[17][23];
    ele[17][20] != ele[17][24];
    ele[17][20] != ele[18][20];
    ele[17][20] != ele[18][21];
    ele[17][20] != ele[18][22];
    ele[17][20] != ele[18][23];
    ele[17][20] != ele[18][24];
    ele[17][20] != ele[19][20];
    ele[17][20] != ele[19][21];
    ele[17][20] != ele[19][22];
    ele[17][20] != ele[19][23];
    ele[17][20] != ele[19][24];
    ele[17][20] != ele[20][20];
    ele[17][20] != ele[21][20];
    ele[17][20] != ele[22][20];
    ele[17][20] != ele[23][20];
    ele[17][20] != ele[24][20];
    ele[17][21] != ele[17][22];
    ele[17][21] != ele[17][23];
    ele[17][21] != ele[17][24];
    ele[17][21] != ele[18][20];
    ele[17][21] != ele[18][21];
    ele[17][21] != ele[18][22];
    ele[17][21] != ele[18][23];
    ele[17][21] != ele[18][24];
    ele[17][21] != ele[19][20];
    ele[17][21] != ele[19][21];
    ele[17][21] != ele[19][22];
    ele[17][21] != ele[19][23];
    ele[17][21] != ele[19][24];
    ele[17][21] != ele[20][21];
    ele[17][21] != ele[21][21];
    ele[17][21] != ele[22][21];
    ele[17][21] != ele[23][21];
    ele[17][21] != ele[24][21];
    ele[17][22] != ele[17][23];
    ele[17][22] != ele[17][24];
    ele[17][22] != ele[18][20];
    ele[17][22] != ele[18][21];
    ele[17][22] != ele[18][22];
    ele[17][22] != ele[18][23];
    ele[17][22] != ele[18][24];
    ele[17][22] != ele[19][20];
    ele[17][22] != ele[19][21];
    ele[17][22] != ele[19][22];
    ele[17][22] != ele[19][23];
    ele[17][22] != ele[19][24];
    ele[17][22] != ele[20][22];
    ele[17][22] != ele[21][22];
    ele[17][22] != ele[22][22];
    ele[17][22] != ele[23][22];
    ele[17][22] != ele[24][22];
    ele[17][23] != ele[17][24];
    ele[17][23] != ele[18][20];
    ele[17][23] != ele[18][21];
    ele[17][23] != ele[18][22];
    ele[17][23] != ele[18][23];
    ele[17][23] != ele[18][24];
    ele[17][23] != ele[19][20];
    ele[17][23] != ele[19][21];
    ele[17][23] != ele[19][22];
    ele[17][23] != ele[19][23];
    ele[17][23] != ele[19][24];
    ele[17][23] != ele[20][23];
    ele[17][23] != ele[21][23];
    ele[17][23] != ele[22][23];
    ele[17][23] != ele[23][23];
    ele[17][23] != ele[24][23];
    ele[17][24] != ele[18][20];
    ele[17][24] != ele[18][21];
    ele[17][24] != ele[18][22];
    ele[17][24] != ele[18][23];
    ele[17][24] != ele[18][24];
    ele[17][24] != ele[19][20];
    ele[17][24] != ele[19][21];
    ele[17][24] != ele[19][22];
    ele[17][24] != ele[19][23];
    ele[17][24] != ele[19][24];
    ele[17][24] != ele[20][24];
    ele[17][24] != ele[21][24];
    ele[17][24] != ele[22][24];
    ele[17][24] != ele[23][24];
    ele[17][24] != ele[24][24];
    ele[17][3] != ele[17][10];
    ele[17][3] != ele[17][11];
    ele[17][3] != ele[17][12];
    ele[17][3] != ele[17][13];
    ele[17][3] != ele[17][14];
    ele[17][3] != ele[17][15];
    ele[17][3] != ele[17][16];
    ele[17][3] != ele[17][17];
    ele[17][3] != ele[17][18];
    ele[17][3] != ele[17][19];
    ele[17][3] != ele[17][20];
    ele[17][3] != ele[17][21];
    ele[17][3] != ele[17][22];
    ele[17][3] != ele[17][23];
    ele[17][3] != ele[17][24];
    ele[17][3] != ele[17][4];
    ele[17][3] != ele[17][5];
    ele[17][3] != ele[17][6];
    ele[17][3] != ele[17][7];
    ele[17][3] != ele[17][8];
    ele[17][3] != ele[17][9];
    ele[17][3] != ele[18][0];
    ele[17][3] != ele[18][1];
    ele[17][3] != ele[18][2];
    ele[17][3] != ele[18][3];
    ele[17][3] != ele[18][4];
    ele[17][3] != ele[19][0];
    ele[17][3] != ele[19][1];
    ele[17][3] != ele[19][2];
    ele[17][3] != ele[19][3];
    ele[17][3] != ele[19][4];
    ele[17][3] != ele[20][3];
    ele[17][3] != ele[21][3];
    ele[17][3] != ele[22][3];
    ele[17][3] != ele[23][3];
    ele[17][3] != ele[24][3];
    ele[17][4] != ele[17][10];
    ele[17][4] != ele[17][11];
    ele[17][4] != ele[17][12];
    ele[17][4] != ele[17][13];
    ele[17][4] != ele[17][14];
    ele[17][4] != ele[17][15];
    ele[17][4] != ele[17][16];
    ele[17][4] != ele[17][17];
    ele[17][4] != ele[17][18];
    ele[17][4] != ele[17][19];
    ele[17][4] != ele[17][20];
    ele[17][4] != ele[17][21];
    ele[17][4] != ele[17][22];
    ele[17][4] != ele[17][23];
    ele[17][4] != ele[17][24];
    ele[17][4] != ele[17][5];
    ele[17][4] != ele[17][6];
    ele[17][4] != ele[17][7];
    ele[17][4] != ele[17][8];
    ele[17][4] != ele[17][9];
    ele[17][4] != ele[18][0];
    ele[17][4] != ele[18][1];
    ele[17][4] != ele[18][2];
    ele[17][4] != ele[18][3];
    ele[17][4] != ele[18][4];
    ele[17][4] != ele[19][0];
    ele[17][4] != ele[19][1];
    ele[17][4] != ele[19][2];
    ele[17][4] != ele[19][3];
    ele[17][4] != ele[19][4];
    ele[17][4] != ele[20][4];
    ele[17][4] != ele[21][4];
    ele[17][4] != ele[22][4];
    ele[17][4] != ele[23][4];
    ele[17][4] != ele[24][4];
    ele[17][5] != ele[17][10];
    ele[17][5] != ele[17][11];
    ele[17][5] != ele[17][12];
    ele[17][5] != ele[17][13];
    ele[17][5] != ele[17][14];
    ele[17][5] != ele[17][15];
    ele[17][5] != ele[17][16];
    ele[17][5] != ele[17][17];
    ele[17][5] != ele[17][18];
    ele[17][5] != ele[17][19];
    ele[17][5] != ele[17][20];
    ele[17][5] != ele[17][21];
    ele[17][5] != ele[17][22];
    ele[17][5] != ele[17][23];
    ele[17][5] != ele[17][24];
    ele[17][5] != ele[17][6];
    ele[17][5] != ele[17][7];
    ele[17][5] != ele[17][8];
    ele[17][5] != ele[17][9];
    ele[17][5] != ele[18][5];
    ele[17][5] != ele[18][6];
    ele[17][5] != ele[18][7];
    ele[17][5] != ele[18][8];
    ele[17][5] != ele[18][9];
    ele[17][5] != ele[19][5];
    ele[17][5] != ele[19][6];
    ele[17][5] != ele[19][7];
    ele[17][5] != ele[19][8];
    ele[17][5] != ele[19][9];
    ele[17][5] != ele[20][5];
    ele[17][5] != ele[21][5];
    ele[17][5] != ele[22][5];
    ele[17][5] != ele[23][5];
    ele[17][5] != ele[24][5];
    ele[17][6] != ele[17][10];
    ele[17][6] != ele[17][11];
    ele[17][6] != ele[17][12];
    ele[17][6] != ele[17][13];
    ele[17][6] != ele[17][14];
    ele[17][6] != ele[17][15];
    ele[17][6] != ele[17][16];
    ele[17][6] != ele[17][17];
    ele[17][6] != ele[17][18];
    ele[17][6] != ele[17][19];
    ele[17][6] != ele[17][20];
    ele[17][6] != ele[17][21];
    ele[17][6] != ele[17][22];
    ele[17][6] != ele[17][23];
    ele[17][6] != ele[17][24];
    ele[17][6] != ele[17][7];
    ele[17][6] != ele[17][8];
    ele[17][6] != ele[17][9];
    ele[17][6] != ele[18][5];
    ele[17][6] != ele[18][6];
    ele[17][6] != ele[18][7];
    ele[17][6] != ele[18][8];
    ele[17][6] != ele[18][9];
    ele[17][6] != ele[19][5];
    ele[17][6] != ele[19][6];
    ele[17][6] != ele[19][7];
    ele[17][6] != ele[19][8];
    ele[17][6] != ele[19][9];
    ele[17][6] != ele[20][6];
    ele[17][6] != ele[21][6];
    ele[17][6] != ele[22][6];
    ele[17][6] != ele[23][6];
    ele[17][6] != ele[24][6];
    ele[17][7] != ele[17][10];
    ele[17][7] != ele[17][11];
    ele[17][7] != ele[17][12];
    ele[17][7] != ele[17][13];
    ele[17][7] != ele[17][14];
    ele[17][7] != ele[17][15];
    ele[17][7] != ele[17][16];
    ele[17][7] != ele[17][17];
    ele[17][7] != ele[17][18];
    ele[17][7] != ele[17][19];
    ele[17][7] != ele[17][20];
    ele[17][7] != ele[17][21];
    ele[17][7] != ele[17][22];
    ele[17][7] != ele[17][23];
    ele[17][7] != ele[17][24];
    ele[17][7] != ele[17][8];
    ele[17][7] != ele[17][9];
    ele[17][7] != ele[18][5];
    ele[17][7] != ele[18][6];
    ele[17][7] != ele[18][7];
    ele[17][7] != ele[18][8];
    ele[17][7] != ele[18][9];
    ele[17][7] != ele[19][5];
    ele[17][7] != ele[19][6];
    ele[17][7] != ele[19][7];
    ele[17][7] != ele[19][8];
    ele[17][7] != ele[19][9];
    ele[17][7] != ele[20][7];
    ele[17][7] != ele[21][7];
    ele[17][7] != ele[22][7];
    ele[17][7] != ele[23][7];
    ele[17][7] != ele[24][7];
    ele[17][8] != ele[17][10];
    ele[17][8] != ele[17][11];
    ele[17][8] != ele[17][12];
    ele[17][8] != ele[17][13];
    ele[17][8] != ele[17][14];
    ele[17][8] != ele[17][15];
    ele[17][8] != ele[17][16];
    ele[17][8] != ele[17][17];
    ele[17][8] != ele[17][18];
    ele[17][8] != ele[17][19];
    ele[17][8] != ele[17][20];
    ele[17][8] != ele[17][21];
    ele[17][8] != ele[17][22];
    ele[17][8] != ele[17][23];
    ele[17][8] != ele[17][24];
    ele[17][8] != ele[17][9];
    ele[17][8] != ele[18][5];
    ele[17][8] != ele[18][6];
    ele[17][8] != ele[18][7];
    ele[17][8] != ele[18][8];
    ele[17][8] != ele[18][9];
    ele[17][8] != ele[19][5];
    ele[17][8] != ele[19][6];
    ele[17][8] != ele[19][7];
    ele[17][8] != ele[19][8];
    ele[17][8] != ele[19][9];
    ele[17][8] != ele[20][8];
    ele[17][8] != ele[21][8];
    ele[17][8] != ele[22][8];
    ele[17][8] != ele[23][8];
    ele[17][8] != ele[24][8];
    ele[17][9] != ele[17][10];
    ele[17][9] != ele[17][11];
    ele[17][9] != ele[17][12];
    ele[17][9] != ele[17][13];
    ele[17][9] != ele[17][14];
    ele[17][9] != ele[17][15];
    ele[17][9] != ele[17][16];
    ele[17][9] != ele[17][17];
    ele[17][9] != ele[17][18];
    ele[17][9] != ele[17][19];
    ele[17][9] != ele[17][20];
    ele[17][9] != ele[17][21];
    ele[17][9] != ele[17][22];
    ele[17][9] != ele[17][23];
    ele[17][9] != ele[17][24];
    ele[17][9] != ele[18][5];
    ele[17][9] != ele[18][6];
    ele[17][9] != ele[18][7];
    ele[17][9] != ele[18][8];
    ele[17][9] != ele[18][9];
    ele[17][9] != ele[19][5];
    ele[17][9] != ele[19][6];
    ele[17][9] != ele[19][7];
    ele[17][9] != ele[19][8];
    ele[17][9] != ele[19][9];
    ele[17][9] != ele[20][9];
    ele[17][9] != ele[21][9];
    ele[17][9] != ele[22][9];
    ele[17][9] != ele[23][9];
    ele[17][9] != ele[24][9];
    ele[18][0] != ele[18][1];
    ele[18][0] != ele[18][10];
    ele[18][0] != ele[18][11];
    ele[18][0] != ele[18][12];
    ele[18][0] != ele[18][13];
    ele[18][0] != ele[18][14];
    ele[18][0] != ele[18][15];
    ele[18][0] != ele[18][16];
    ele[18][0] != ele[18][17];
    ele[18][0] != ele[18][18];
    ele[18][0] != ele[18][19];
    ele[18][0] != ele[18][2];
    ele[18][0] != ele[18][20];
    ele[18][0] != ele[18][21];
    ele[18][0] != ele[18][22];
    ele[18][0] != ele[18][23];
    ele[18][0] != ele[18][24];
    ele[18][0] != ele[18][3];
    ele[18][0] != ele[18][4];
    ele[18][0] != ele[18][5];
    ele[18][0] != ele[18][6];
    ele[18][0] != ele[18][7];
    ele[18][0] != ele[18][8];
    ele[18][0] != ele[18][9];
    ele[18][0] != ele[19][0];
    ele[18][0] != ele[19][1];
    ele[18][0] != ele[19][2];
    ele[18][0] != ele[19][3];
    ele[18][0] != ele[19][4];
    ele[18][0] != ele[20][0];
    ele[18][0] != ele[21][0];
    ele[18][0] != ele[22][0];
    ele[18][0] != ele[23][0];
    ele[18][0] != ele[24][0];
    ele[18][1] != ele[18][10];
    ele[18][1] != ele[18][11];
    ele[18][1] != ele[18][12];
    ele[18][1] != ele[18][13];
    ele[18][1] != ele[18][14];
    ele[18][1] != ele[18][15];
    ele[18][1] != ele[18][16];
    ele[18][1] != ele[18][17];
    ele[18][1] != ele[18][18];
    ele[18][1] != ele[18][19];
    ele[18][1] != ele[18][2];
    ele[18][1] != ele[18][20];
    ele[18][1] != ele[18][21];
    ele[18][1] != ele[18][22];
    ele[18][1] != ele[18][23];
    ele[18][1] != ele[18][24];
    ele[18][1] != ele[18][3];
    ele[18][1] != ele[18][4];
    ele[18][1] != ele[18][5];
    ele[18][1] != ele[18][6];
    ele[18][1] != ele[18][7];
    ele[18][1] != ele[18][8];
    ele[18][1] != ele[18][9];
    ele[18][1] != ele[19][0];
    ele[18][1] != ele[19][1];
    ele[18][1] != ele[19][2];
    ele[18][1] != ele[19][3];
    ele[18][1] != ele[19][4];
    ele[18][1] != ele[20][1];
    ele[18][1] != ele[21][1];
    ele[18][1] != ele[22][1];
    ele[18][1] != ele[23][1];
    ele[18][1] != ele[24][1];
    ele[18][10] != ele[18][11];
    ele[18][10] != ele[18][12];
    ele[18][10] != ele[18][13];
    ele[18][10] != ele[18][14];
    ele[18][10] != ele[18][15];
    ele[18][10] != ele[18][16];
    ele[18][10] != ele[18][17];
    ele[18][10] != ele[18][18];
    ele[18][10] != ele[18][19];
    ele[18][10] != ele[18][20];
    ele[18][10] != ele[18][21];
    ele[18][10] != ele[18][22];
    ele[18][10] != ele[18][23];
    ele[18][10] != ele[18][24];
    ele[18][10] != ele[19][10];
    ele[18][10] != ele[19][11];
    ele[18][10] != ele[19][12];
    ele[18][10] != ele[19][13];
    ele[18][10] != ele[19][14];
    ele[18][10] != ele[20][10];
    ele[18][10] != ele[21][10];
    ele[18][10] != ele[22][10];
    ele[18][10] != ele[23][10];
    ele[18][10] != ele[24][10];
    ele[18][11] != ele[18][12];
    ele[18][11] != ele[18][13];
    ele[18][11] != ele[18][14];
    ele[18][11] != ele[18][15];
    ele[18][11] != ele[18][16];
    ele[18][11] != ele[18][17];
    ele[18][11] != ele[18][18];
    ele[18][11] != ele[18][19];
    ele[18][11] != ele[18][20];
    ele[18][11] != ele[18][21];
    ele[18][11] != ele[18][22];
    ele[18][11] != ele[18][23];
    ele[18][11] != ele[18][24];
    ele[18][11] != ele[19][10];
    ele[18][11] != ele[19][11];
    ele[18][11] != ele[19][12];
    ele[18][11] != ele[19][13];
    ele[18][11] != ele[19][14];
    ele[18][11] != ele[20][11];
    ele[18][11] != ele[21][11];
    ele[18][11] != ele[22][11];
    ele[18][11] != ele[23][11];
    ele[18][11] != ele[24][11];
    ele[18][12] != ele[18][13];
    ele[18][12] != ele[18][14];
    ele[18][12] != ele[18][15];
    ele[18][12] != ele[18][16];
    ele[18][12] != ele[18][17];
    ele[18][12] != ele[18][18];
    ele[18][12] != ele[18][19];
    ele[18][12] != ele[18][20];
    ele[18][12] != ele[18][21];
    ele[18][12] != ele[18][22];
    ele[18][12] != ele[18][23];
    ele[18][12] != ele[18][24];
    ele[18][12] != ele[19][10];
    ele[18][12] != ele[19][11];
    ele[18][12] != ele[19][12];
    ele[18][12] != ele[19][13];
    ele[18][12] != ele[19][14];
    ele[18][12] != ele[20][12];
    ele[18][12] != ele[21][12];
    ele[18][12] != ele[22][12];
    ele[18][12] != ele[23][12];
    ele[18][12] != ele[24][12];
    ele[18][13] != ele[18][14];
    ele[18][13] != ele[18][15];
    ele[18][13] != ele[18][16];
    ele[18][13] != ele[18][17];
    ele[18][13] != ele[18][18];
    ele[18][13] != ele[18][19];
    ele[18][13] != ele[18][20];
    ele[18][13] != ele[18][21];
    ele[18][13] != ele[18][22];
    ele[18][13] != ele[18][23];
    ele[18][13] != ele[18][24];
    ele[18][13] != ele[19][10];
    ele[18][13] != ele[19][11];
    ele[18][13] != ele[19][12];
    ele[18][13] != ele[19][13];
    ele[18][13] != ele[19][14];
    ele[18][13] != ele[20][13];
    ele[18][13] != ele[21][13];
    ele[18][13] != ele[22][13];
    ele[18][13] != ele[23][13];
    ele[18][13] != ele[24][13];
    ele[18][14] != ele[18][15];
    ele[18][14] != ele[18][16];
    ele[18][14] != ele[18][17];
    ele[18][14] != ele[18][18];
    ele[18][14] != ele[18][19];
    ele[18][14] != ele[18][20];
    ele[18][14] != ele[18][21];
    ele[18][14] != ele[18][22];
    ele[18][14] != ele[18][23];
    ele[18][14] != ele[18][24];
    ele[18][14] != ele[19][10];
    ele[18][14] != ele[19][11];
    ele[18][14] != ele[19][12];
    ele[18][14] != ele[19][13];
    ele[18][14] != ele[19][14];
    ele[18][14] != ele[20][14];
    ele[18][14] != ele[21][14];
    ele[18][14] != ele[22][14];
    ele[18][14] != ele[23][14];
    ele[18][14] != ele[24][14];
    ele[18][15] != ele[18][16];
    ele[18][15] != ele[18][17];
    ele[18][15] != ele[18][18];
    ele[18][15] != ele[18][19];
    ele[18][15] != ele[18][20];
    ele[18][15] != ele[18][21];
    ele[18][15] != ele[18][22];
    ele[18][15] != ele[18][23];
    ele[18][15] != ele[18][24];
    ele[18][15] != ele[19][15];
    ele[18][15] != ele[19][16];
    ele[18][15] != ele[19][17];
    ele[18][15] != ele[19][18];
    ele[18][15] != ele[19][19];
    ele[18][15] != ele[20][15];
    ele[18][15] != ele[21][15];
    ele[18][15] != ele[22][15];
    ele[18][15] != ele[23][15];
    ele[18][15] != ele[24][15];
    ele[18][16] != ele[18][17];
    ele[18][16] != ele[18][18];
    ele[18][16] != ele[18][19];
    ele[18][16] != ele[18][20];
    ele[18][16] != ele[18][21];
    ele[18][16] != ele[18][22];
    ele[18][16] != ele[18][23];
    ele[18][16] != ele[18][24];
    ele[18][16] != ele[19][15];
    ele[18][16] != ele[19][16];
    ele[18][16] != ele[19][17];
    ele[18][16] != ele[19][18];
    ele[18][16] != ele[19][19];
    ele[18][16] != ele[20][16];
    ele[18][16] != ele[21][16];
    ele[18][16] != ele[22][16];
    ele[18][16] != ele[23][16];
    ele[18][16] != ele[24][16];
    ele[18][17] != ele[18][18];
    ele[18][17] != ele[18][19];
    ele[18][17] != ele[18][20];
    ele[18][17] != ele[18][21];
    ele[18][17] != ele[18][22];
    ele[18][17] != ele[18][23];
    ele[18][17] != ele[18][24];
    ele[18][17] != ele[19][15];
    ele[18][17] != ele[19][16];
    ele[18][17] != ele[19][17];
    ele[18][17] != ele[19][18];
    ele[18][17] != ele[19][19];
    ele[18][17] != ele[20][17];
    ele[18][17] != ele[21][17];
    ele[18][17] != ele[22][17];
    ele[18][17] != ele[23][17];
    ele[18][17] != ele[24][17];
    ele[18][18] != ele[18][19];
    ele[18][18] != ele[18][20];
    ele[18][18] != ele[18][21];
    ele[18][18] != ele[18][22];
    ele[18][18] != ele[18][23];
    ele[18][18] != ele[18][24];
    ele[18][18] != ele[19][15];
    ele[18][18] != ele[19][16];
    ele[18][18] != ele[19][17];
    ele[18][18] != ele[19][18];
    ele[18][18] != ele[19][19];
    ele[18][18] != ele[20][18];
    ele[18][18] != ele[21][18];
    ele[18][18] != ele[22][18];
    ele[18][18] != ele[23][18];
    ele[18][18] != ele[24][18];
    ele[18][19] != ele[18][20];
    ele[18][19] != ele[18][21];
    ele[18][19] != ele[18][22];
    ele[18][19] != ele[18][23];
    ele[18][19] != ele[18][24];
    ele[18][19] != ele[19][15];
    ele[18][19] != ele[19][16];
    ele[18][19] != ele[19][17];
    ele[18][19] != ele[19][18];
    ele[18][19] != ele[19][19];
    ele[18][19] != ele[20][19];
    ele[18][19] != ele[21][19];
    ele[18][19] != ele[22][19];
    ele[18][19] != ele[23][19];
    ele[18][19] != ele[24][19];
    ele[18][2] != ele[18][10];
    ele[18][2] != ele[18][11];
    ele[18][2] != ele[18][12];
    ele[18][2] != ele[18][13];
    ele[18][2] != ele[18][14];
    ele[18][2] != ele[18][15];
    ele[18][2] != ele[18][16];
    ele[18][2] != ele[18][17];
    ele[18][2] != ele[18][18];
    ele[18][2] != ele[18][19];
    ele[18][2] != ele[18][20];
    ele[18][2] != ele[18][21];
    ele[18][2] != ele[18][22];
    ele[18][2] != ele[18][23];
    ele[18][2] != ele[18][24];
    ele[18][2] != ele[18][3];
    ele[18][2] != ele[18][4];
    ele[18][2] != ele[18][5];
    ele[18][2] != ele[18][6];
    ele[18][2] != ele[18][7];
    ele[18][2] != ele[18][8];
    ele[18][2] != ele[18][9];
    ele[18][2] != ele[19][0];
    ele[18][2] != ele[19][1];
    ele[18][2] != ele[19][2];
    ele[18][2] != ele[19][3];
    ele[18][2] != ele[19][4];
    ele[18][2] != ele[20][2];
    ele[18][2] != ele[21][2];
    ele[18][2] != ele[22][2];
    ele[18][2] != ele[23][2];
    ele[18][2] != ele[24][2];
    ele[18][20] != ele[18][21];
    ele[18][20] != ele[18][22];
    ele[18][20] != ele[18][23];
    ele[18][20] != ele[18][24];
    ele[18][20] != ele[19][20];
    ele[18][20] != ele[19][21];
    ele[18][20] != ele[19][22];
    ele[18][20] != ele[19][23];
    ele[18][20] != ele[19][24];
    ele[18][20] != ele[20][20];
    ele[18][20] != ele[21][20];
    ele[18][20] != ele[22][20];
    ele[18][20] != ele[23][20];
    ele[18][20] != ele[24][20];
    ele[18][21] != ele[18][22];
    ele[18][21] != ele[18][23];
    ele[18][21] != ele[18][24];
    ele[18][21] != ele[19][20];
    ele[18][21] != ele[19][21];
    ele[18][21] != ele[19][22];
    ele[18][21] != ele[19][23];
    ele[18][21] != ele[19][24];
    ele[18][21] != ele[20][21];
    ele[18][21] != ele[21][21];
    ele[18][21] != ele[22][21];
    ele[18][21] != ele[23][21];
    ele[18][21] != ele[24][21];
    ele[18][22] != ele[18][23];
    ele[18][22] != ele[18][24];
    ele[18][22] != ele[19][20];
    ele[18][22] != ele[19][21];
    ele[18][22] != ele[19][22];
    ele[18][22] != ele[19][23];
    ele[18][22] != ele[19][24];
    ele[18][22] != ele[20][22];
    ele[18][22] != ele[21][22];
    ele[18][22] != ele[22][22];
    ele[18][22] != ele[23][22];
    ele[18][22] != ele[24][22];
    ele[18][23] != ele[18][24];
    ele[18][23] != ele[19][20];
    ele[18][23] != ele[19][21];
    ele[18][23] != ele[19][22];
    ele[18][23] != ele[19][23];
    ele[18][23] != ele[19][24];
    ele[18][23] != ele[20][23];
    ele[18][23] != ele[21][23];
    ele[18][23] != ele[22][23];
    ele[18][23] != ele[23][23];
    ele[18][23] != ele[24][23];
    ele[18][24] != ele[19][20];
    ele[18][24] != ele[19][21];
    ele[18][24] != ele[19][22];
    ele[18][24] != ele[19][23];
    ele[18][24] != ele[19][24];
    ele[18][24] != ele[20][24];
    ele[18][24] != ele[21][24];
    ele[18][24] != ele[22][24];
    ele[18][24] != ele[23][24];
    ele[18][24] != ele[24][24];
    ele[18][3] != ele[18][10];
    ele[18][3] != ele[18][11];
    ele[18][3] != ele[18][12];
    ele[18][3] != ele[18][13];
    ele[18][3] != ele[18][14];
    ele[18][3] != ele[18][15];
    ele[18][3] != ele[18][16];
    ele[18][3] != ele[18][17];
    ele[18][3] != ele[18][18];
    ele[18][3] != ele[18][19];
    ele[18][3] != ele[18][20];
    ele[18][3] != ele[18][21];
    ele[18][3] != ele[18][22];
    ele[18][3] != ele[18][23];
    ele[18][3] != ele[18][24];
    ele[18][3] != ele[18][4];
    ele[18][3] != ele[18][5];
    ele[18][3] != ele[18][6];
    ele[18][3] != ele[18][7];
    ele[18][3] != ele[18][8];
    ele[18][3] != ele[18][9];
    ele[18][3] != ele[19][0];
    ele[18][3] != ele[19][1];
    ele[18][3] != ele[19][2];
    ele[18][3] != ele[19][3];
    ele[18][3] != ele[19][4];
    ele[18][3] != ele[20][3];
    ele[18][3] != ele[21][3];
    ele[18][3] != ele[22][3];
    ele[18][3] != ele[23][3];
    ele[18][3] != ele[24][3];
    ele[18][4] != ele[18][10];
    ele[18][4] != ele[18][11];
    ele[18][4] != ele[18][12];
    ele[18][4] != ele[18][13];
    ele[18][4] != ele[18][14];
    ele[18][4] != ele[18][15];
    ele[18][4] != ele[18][16];
    ele[18][4] != ele[18][17];
    ele[18][4] != ele[18][18];
    ele[18][4] != ele[18][19];
    ele[18][4] != ele[18][20];
    ele[18][4] != ele[18][21];
    ele[18][4] != ele[18][22];
    ele[18][4] != ele[18][23];
    ele[18][4] != ele[18][24];
    ele[18][4] != ele[18][5];
    ele[18][4] != ele[18][6];
    ele[18][4] != ele[18][7];
    ele[18][4] != ele[18][8];
    ele[18][4] != ele[18][9];
    ele[18][4] != ele[19][0];
    ele[18][4] != ele[19][1];
    ele[18][4] != ele[19][2];
    ele[18][4] != ele[19][3];
    ele[18][4] != ele[19][4];
    ele[18][4] != ele[20][4];
    ele[18][4] != ele[21][4];
    ele[18][4] != ele[22][4];
    ele[18][4] != ele[23][4];
    ele[18][4] != ele[24][4];
    ele[18][5] != ele[18][10];
    ele[18][5] != ele[18][11];
    ele[18][5] != ele[18][12];
    ele[18][5] != ele[18][13];
    ele[18][5] != ele[18][14];
    ele[18][5] != ele[18][15];
    ele[18][5] != ele[18][16];
    ele[18][5] != ele[18][17];
    ele[18][5] != ele[18][18];
    ele[18][5] != ele[18][19];
    ele[18][5] != ele[18][20];
    ele[18][5] != ele[18][21];
    ele[18][5] != ele[18][22];
    ele[18][5] != ele[18][23];
    ele[18][5] != ele[18][24];
    ele[18][5] != ele[18][6];
    ele[18][5] != ele[18][7];
    ele[18][5] != ele[18][8];
    ele[18][5] != ele[18][9];
    ele[18][5] != ele[19][5];
    ele[18][5] != ele[19][6];
    ele[18][5] != ele[19][7];
    ele[18][5] != ele[19][8];
    ele[18][5] != ele[19][9];
    ele[18][5] != ele[20][5];
    ele[18][5] != ele[21][5];
    ele[18][5] != ele[22][5];
    ele[18][5] != ele[23][5];
    ele[18][5] != ele[24][5];
    ele[18][6] != ele[18][10];
    ele[18][6] != ele[18][11];
    ele[18][6] != ele[18][12];
    ele[18][6] != ele[18][13];
    ele[18][6] != ele[18][14];
    ele[18][6] != ele[18][15];
    ele[18][6] != ele[18][16];
    ele[18][6] != ele[18][17];
    ele[18][6] != ele[18][18];
    ele[18][6] != ele[18][19];
    ele[18][6] != ele[18][20];
    ele[18][6] != ele[18][21];
    ele[18][6] != ele[18][22];
    ele[18][6] != ele[18][23];
    ele[18][6] != ele[18][24];
    ele[18][6] != ele[18][7];
    ele[18][6] != ele[18][8];
    ele[18][6] != ele[18][9];
    ele[18][6] != ele[19][5];
    ele[18][6] != ele[19][6];
    ele[18][6] != ele[19][7];
    ele[18][6] != ele[19][8];
    ele[18][6] != ele[19][9];
    ele[18][6] != ele[20][6];
    ele[18][6] != ele[21][6];
    ele[18][6] != ele[22][6];
    ele[18][6] != ele[23][6];
    ele[18][6] != ele[24][6];
    ele[18][7] != ele[18][10];
    ele[18][7] != ele[18][11];
    ele[18][7] != ele[18][12];
    ele[18][7] != ele[18][13];
    ele[18][7] != ele[18][14];
    ele[18][7] != ele[18][15];
    ele[18][7] != ele[18][16];
    ele[18][7] != ele[18][17];
    ele[18][7] != ele[18][18];
    ele[18][7] != ele[18][19];
    ele[18][7] != ele[18][20];
    ele[18][7] != ele[18][21];
    ele[18][7] != ele[18][22];
    ele[18][7] != ele[18][23];
    ele[18][7] != ele[18][24];
    ele[18][7] != ele[18][8];
    ele[18][7] != ele[18][9];
    ele[18][7] != ele[19][5];
    ele[18][7] != ele[19][6];
    ele[18][7] != ele[19][7];
    ele[18][7] != ele[19][8];
    ele[18][7] != ele[19][9];
    ele[18][7] != ele[20][7];
    ele[18][7] != ele[21][7];
    ele[18][7] != ele[22][7];
    ele[18][7] != ele[23][7];
    ele[18][7] != ele[24][7];
    ele[18][8] != ele[18][10];
    ele[18][8] != ele[18][11];
    ele[18][8] != ele[18][12];
    ele[18][8] != ele[18][13];
    ele[18][8] != ele[18][14];
    ele[18][8] != ele[18][15];
    ele[18][8] != ele[18][16];
    ele[18][8] != ele[18][17];
    ele[18][8] != ele[18][18];
    ele[18][8] != ele[18][19];
    ele[18][8] != ele[18][20];
    ele[18][8] != ele[18][21];
    ele[18][8] != ele[18][22];
    ele[18][8] != ele[18][23];
    ele[18][8] != ele[18][24];
    ele[18][8] != ele[18][9];
    ele[18][8] != ele[19][5];
    ele[18][8] != ele[19][6];
    ele[18][8] != ele[19][7];
    ele[18][8] != ele[19][8];
    ele[18][8] != ele[19][9];
    ele[18][8] != ele[20][8];
    ele[18][8] != ele[21][8];
    ele[18][8] != ele[22][8];
    ele[18][8] != ele[23][8];
    ele[18][8] != ele[24][8];
    ele[18][9] != ele[18][10];
    ele[18][9] != ele[18][11];
    ele[18][9] != ele[18][12];
    ele[18][9] != ele[18][13];
    ele[18][9] != ele[18][14];
    ele[18][9] != ele[18][15];
    ele[18][9] != ele[18][16];
    ele[18][9] != ele[18][17];
    ele[18][9] != ele[18][18];
    ele[18][9] != ele[18][19];
    ele[18][9] != ele[18][20];
    ele[18][9] != ele[18][21];
    ele[18][9] != ele[18][22];
    ele[18][9] != ele[18][23];
    ele[18][9] != ele[18][24];
    ele[18][9] != ele[19][5];
    ele[18][9] != ele[19][6];
    ele[18][9] != ele[19][7];
    ele[18][9] != ele[19][8];
    ele[18][9] != ele[19][9];
    ele[18][9] != ele[20][9];
    ele[18][9] != ele[21][9];
    ele[18][9] != ele[22][9];
    ele[18][9] != ele[23][9];
    ele[18][9] != ele[24][9];
    ele[19][0] != ele[19][1];
    ele[19][0] != ele[19][10];
    ele[19][0] != ele[19][11];
    ele[19][0] != ele[19][12];
    ele[19][0] != ele[19][13];
    ele[19][0] != ele[19][14];
    ele[19][0] != ele[19][15];
    ele[19][0] != ele[19][16];
    ele[19][0] != ele[19][17];
    ele[19][0] != ele[19][18];
    ele[19][0] != ele[19][19];
    ele[19][0] != ele[19][2];
    ele[19][0] != ele[19][20];
    ele[19][0] != ele[19][21];
    ele[19][0] != ele[19][22];
    ele[19][0] != ele[19][23];
    ele[19][0] != ele[19][24];
    ele[19][0] != ele[19][3];
    ele[19][0] != ele[19][4];
    ele[19][0] != ele[19][5];
    ele[19][0] != ele[19][6];
    ele[19][0] != ele[19][7];
    ele[19][0] != ele[19][8];
    ele[19][0] != ele[19][9];
    ele[19][0] != ele[20][0];
    ele[19][0] != ele[21][0];
    ele[19][0] != ele[22][0];
    ele[19][0] != ele[23][0];
    ele[19][0] != ele[24][0];
    ele[19][1] != ele[19][10];
    ele[19][1] != ele[19][11];
    ele[19][1] != ele[19][12];
    ele[19][1] != ele[19][13];
    ele[19][1] != ele[19][14];
    ele[19][1] != ele[19][15];
    ele[19][1] != ele[19][16];
    ele[19][1] != ele[19][17];
    ele[19][1] != ele[19][18];
    ele[19][1] != ele[19][19];
    ele[19][1] != ele[19][2];
    ele[19][1] != ele[19][20];
    ele[19][1] != ele[19][21];
    ele[19][1] != ele[19][22];
    ele[19][1] != ele[19][23];
    ele[19][1] != ele[19][24];
    ele[19][1] != ele[19][3];
    ele[19][1] != ele[19][4];
    ele[19][1] != ele[19][5];
    ele[19][1] != ele[19][6];
    ele[19][1] != ele[19][7];
    ele[19][1] != ele[19][8];
    ele[19][1] != ele[19][9];
    ele[19][1] != ele[20][1];
    ele[19][1] != ele[21][1];
    ele[19][1] != ele[22][1];
    ele[19][1] != ele[23][1];
    ele[19][1] != ele[24][1];
    ele[19][10] != ele[19][11];
    ele[19][10] != ele[19][12];
    ele[19][10] != ele[19][13];
    ele[19][10] != ele[19][14];
    ele[19][10] != ele[19][15];
    ele[19][10] != ele[19][16];
    ele[19][10] != ele[19][17];
    ele[19][10] != ele[19][18];
    ele[19][10] != ele[19][19];
    ele[19][10] != ele[19][20];
    ele[19][10] != ele[19][21];
    ele[19][10] != ele[19][22];
    ele[19][10] != ele[19][23];
    ele[19][10] != ele[19][24];
    ele[19][10] != ele[20][10];
    ele[19][10] != ele[21][10];
    ele[19][10] != ele[22][10];
    ele[19][10] != ele[23][10];
    ele[19][10] != ele[24][10];
    ele[19][11] != ele[19][12];
    ele[19][11] != ele[19][13];
    ele[19][11] != ele[19][14];
    ele[19][11] != ele[19][15];
    ele[19][11] != ele[19][16];
    ele[19][11] != ele[19][17];
    ele[19][11] != ele[19][18];
    ele[19][11] != ele[19][19];
    ele[19][11] != ele[19][20];
    ele[19][11] != ele[19][21];
    ele[19][11] != ele[19][22];
    ele[19][11] != ele[19][23];
    ele[19][11] != ele[19][24];
    ele[19][11] != ele[20][11];
    ele[19][11] != ele[21][11];
    ele[19][11] != ele[22][11];
    ele[19][11] != ele[23][11];
    ele[19][11] != ele[24][11];
    ele[19][12] != ele[19][13];
    ele[19][12] != ele[19][14];
    ele[19][12] != ele[19][15];
    ele[19][12] != ele[19][16];
    ele[19][12] != ele[19][17];
    ele[19][12] != ele[19][18];
    ele[19][12] != ele[19][19];
    ele[19][12] != ele[19][20];
    ele[19][12] != ele[19][21];
    ele[19][12] != ele[19][22];
    ele[19][12] != ele[19][23];
    ele[19][12] != ele[19][24];
    ele[19][12] != ele[20][12];
    ele[19][12] != ele[21][12];
    ele[19][12] != ele[22][12];
    ele[19][12] != ele[23][12];
    ele[19][12] != ele[24][12];
    ele[19][13] != ele[19][14];
    ele[19][13] != ele[19][15];
    ele[19][13] != ele[19][16];
    ele[19][13] != ele[19][17];
    ele[19][13] != ele[19][18];
    ele[19][13] != ele[19][19];
    ele[19][13] != ele[19][20];
    ele[19][13] != ele[19][21];
    ele[19][13] != ele[19][22];
    ele[19][13] != ele[19][23];
    ele[19][13] != ele[19][24];
    ele[19][13] != ele[20][13];
    ele[19][13] != ele[21][13];
    ele[19][13] != ele[22][13];
    ele[19][13] != ele[23][13];
    ele[19][13] != ele[24][13];
    ele[19][14] != ele[19][15];
    ele[19][14] != ele[19][16];
    ele[19][14] != ele[19][17];
    ele[19][14] != ele[19][18];
    ele[19][14] != ele[19][19];
    ele[19][14] != ele[19][20];
    ele[19][14] != ele[19][21];
    ele[19][14] != ele[19][22];
    ele[19][14] != ele[19][23];
    ele[19][14] != ele[19][24];
    ele[19][14] != ele[20][14];
    ele[19][14] != ele[21][14];
    ele[19][14] != ele[22][14];
    ele[19][14] != ele[23][14];
    ele[19][14] != ele[24][14];
    ele[19][15] != ele[19][16];
    ele[19][15] != ele[19][17];
    ele[19][15] != ele[19][18];
    ele[19][15] != ele[19][19];
    ele[19][15] != ele[19][20];
    ele[19][15] != ele[19][21];
    ele[19][15] != ele[19][22];
    ele[19][15] != ele[19][23];
    ele[19][15] != ele[19][24];
    ele[19][15] != ele[20][15];
    ele[19][15] != ele[21][15];
    ele[19][15] != ele[22][15];
    ele[19][15] != ele[23][15];
    ele[19][15] != ele[24][15];
    ele[19][16] != ele[19][17];
    ele[19][16] != ele[19][18];
    ele[19][16] != ele[19][19];
    ele[19][16] != ele[19][20];
    ele[19][16] != ele[19][21];
    ele[19][16] != ele[19][22];
    ele[19][16] != ele[19][23];
    ele[19][16] != ele[19][24];
    ele[19][16] != ele[20][16];
    ele[19][16] != ele[21][16];
    ele[19][16] != ele[22][16];
    ele[19][16] != ele[23][16];
    ele[19][16] != ele[24][16];
    ele[19][17] != ele[19][18];
    ele[19][17] != ele[19][19];
    ele[19][17] != ele[19][20];
    ele[19][17] != ele[19][21];
    ele[19][17] != ele[19][22];
    ele[19][17] != ele[19][23];
    ele[19][17] != ele[19][24];
    ele[19][17] != ele[20][17];
    ele[19][17] != ele[21][17];
    ele[19][17] != ele[22][17];
    ele[19][17] != ele[23][17];
    ele[19][17] != ele[24][17];
    ele[19][18] != ele[19][19];
    ele[19][18] != ele[19][20];
    ele[19][18] != ele[19][21];
    ele[19][18] != ele[19][22];
    ele[19][18] != ele[19][23];
    ele[19][18] != ele[19][24];
    ele[19][18] != ele[20][18];
    ele[19][18] != ele[21][18];
    ele[19][18] != ele[22][18];
    ele[19][18] != ele[23][18];
    ele[19][18] != ele[24][18];
    ele[19][19] != ele[19][20];
    ele[19][19] != ele[19][21];
    ele[19][19] != ele[19][22];
    ele[19][19] != ele[19][23];
    ele[19][19] != ele[19][24];
    ele[19][19] != ele[20][19];
    ele[19][19] != ele[21][19];
    ele[19][19] != ele[22][19];
    ele[19][19] != ele[23][19];
    ele[19][19] != ele[24][19];
    ele[19][2] != ele[19][10];
    ele[19][2] != ele[19][11];
    ele[19][2] != ele[19][12];
    ele[19][2] != ele[19][13];
    ele[19][2] != ele[19][14];
    ele[19][2] != ele[19][15];
    ele[19][2] != ele[19][16];
    ele[19][2] != ele[19][17];
    ele[19][2] != ele[19][18];
    ele[19][2] != ele[19][19];
    ele[19][2] != ele[19][20];
    ele[19][2] != ele[19][21];
    ele[19][2] != ele[19][22];
    ele[19][2] != ele[19][23];
    ele[19][2] != ele[19][24];
    ele[19][2] != ele[19][3];
    ele[19][2] != ele[19][4];
    ele[19][2] != ele[19][5];
    ele[19][2] != ele[19][6];
    ele[19][2] != ele[19][7];
    ele[19][2] != ele[19][8];
    ele[19][2] != ele[19][9];
    ele[19][2] != ele[20][2];
    ele[19][2] != ele[21][2];
    ele[19][2] != ele[22][2];
    ele[19][2] != ele[23][2];
    ele[19][2] != ele[24][2];
    ele[19][20] != ele[19][21];
    ele[19][20] != ele[19][22];
    ele[19][20] != ele[19][23];
    ele[19][20] != ele[19][24];
    ele[19][20] != ele[20][20];
    ele[19][20] != ele[21][20];
    ele[19][20] != ele[22][20];
    ele[19][20] != ele[23][20];
    ele[19][20] != ele[24][20];
    ele[19][21] != ele[19][22];
    ele[19][21] != ele[19][23];
    ele[19][21] != ele[19][24];
    ele[19][21] != ele[20][21];
    ele[19][21] != ele[21][21];
    ele[19][21] != ele[22][21];
    ele[19][21] != ele[23][21];
    ele[19][21] != ele[24][21];
    ele[19][22] != ele[19][23];
    ele[19][22] != ele[19][24];
    ele[19][22] != ele[20][22];
    ele[19][22] != ele[21][22];
    ele[19][22] != ele[22][22];
    ele[19][22] != ele[23][22];
    ele[19][22] != ele[24][22];
    ele[19][23] != ele[19][24];
    ele[19][23] != ele[20][23];
    ele[19][23] != ele[21][23];
    ele[19][23] != ele[22][23];
    ele[19][23] != ele[23][23];
    ele[19][23] != ele[24][23];
    ele[19][24] != ele[20][24];
    ele[19][24] != ele[21][24];
    ele[19][24] != ele[22][24];
    ele[19][24] != ele[23][24];
    ele[19][24] != ele[24][24];
    ele[19][3] != ele[19][10];
    ele[19][3] != ele[19][11];
    ele[19][3] != ele[19][12];
    ele[19][3] != ele[19][13];
    ele[19][3] != ele[19][14];
    ele[19][3] != ele[19][15];
    ele[19][3] != ele[19][16];
    ele[19][3] != ele[19][17];
    ele[19][3] != ele[19][18];
    ele[19][3] != ele[19][19];
    ele[19][3] != ele[19][20];
    ele[19][3] != ele[19][21];
    ele[19][3] != ele[19][22];
    ele[19][3] != ele[19][23];
    ele[19][3] != ele[19][24];
    ele[19][3] != ele[19][4];
    ele[19][3] != ele[19][5];
    ele[19][3] != ele[19][6];
    ele[19][3] != ele[19][7];
    ele[19][3] != ele[19][8];
    ele[19][3] != ele[19][9];
    ele[19][3] != ele[20][3];
    ele[19][3] != ele[21][3];
    ele[19][3] != ele[22][3];
    ele[19][3] != ele[23][3];
    ele[19][3] != ele[24][3];
    ele[19][4] != ele[19][10];
    ele[19][4] != ele[19][11];
    ele[19][4] != ele[19][12];
    ele[19][4] != ele[19][13];
    ele[19][4] != ele[19][14];
    ele[19][4] != ele[19][15];
    ele[19][4] != ele[19][16];
    ele[19][4] != ele[19][17];
    ele[19][4] != ele[19][18];
    ele[19][4] != ele[19][19];
    ele[19][4] != ele[19][20];
    ele[19][4] != ele[19][21];
    ele[19][4] != ele[19][22];
    ele[19][4] != ele[19][23];
    ele[19][4] != ele[19][24];
    ele[19][4] != ele[19][5];
    ele[19][4] != ele[19][6];
    ele[19][4] != ele[19][7];
    ele[19][4] != ele[19][8];
    ele[19][4] != ele[19][9];
    ele[19][4] != ele[20][4];
    ele[19][4] != ele[21][4];
    ele[19][4] != ele[22][4];
    ele[19][4] != ele[23][4];
    ele[19][4] != ele[24][4];
    ele[19][5] != ele[19][10];
    ele[19][5] != ele[19][11];
    ele[19][5] != ele[19][12];
    ele[19][5] != ele[19][13];
    ele[19][5] != ele[19][14];
    ele[19][5] != ele[19][15];
    ele[19][5] != ele[19][16];
    ele[19][5] != ele[19][17];
    ele[19][5] != ele[19][18];
    ele[19][5] != ele[19][19];
    ele[19][5] != ele[19][20];
    ele[19][5] != ele[19][21];
    ele[19][5] != ele[19][22];
    ele[19][5] != ele[19][23];
    ele[19][5] != ele[19][24];
    ele[19][5] != ele[19][6];
    ele[19][5] != ele[19][7];
    ele[19][5] != ele[19][8];
    ele[19][5] != ele[19][9];
    ele[19][5] != ele[20][5];
    ele[19][5] != ele[21][5];
    ele[19][5] != ele[22][5];
    ele[19][5] != ele[23][5];
    ele[19][5] != ele[24][5];
    ele[19][6] != ele[19][10];
    ele[19][6] != ele[19][11];
    ele[19][6] != ele[19][12];
    ele[19][6] != ele[19][13];
    ele[19][6] != ele[19][14];
    ele[19][6] != ele[19][15];
    ele[19][6] != ele[19][16];
    ele[19][6] != ele[19][17];
    ele[19][6] != ele[19][18];
    ele[19][6] != ele[19][19];
    ele[19][6] != ele[19][20];
    ele[19][6] != ele[19][21];
    ele[19][6] != ele[19][22];
    ele[19][6] != ele[19][23];
    ele[19][6] != ele[19][24];
    ele[19][6] != ele[19][7];
    ele[19][6] != ele[19][8];
    ele[19][6] != ele[19][9];
    ele[19][6] != ele[20][6];
    ele[19][6] != ele[21][6];
    ele[19][6] != ele[22][6];
    ele[19][6] != ele[23][6];
    ele[19][6] != ele[24][6];
    ele[19][7] != ele[19][10];
    ele[19][7] != ele[19][11];
    ele[19][7] != ele[19][12];
    ele[19][7] != ele[19][13];
    ele[19][7] != ele[19][14];
    ele[19][7] != ele[19][15];
    ele[19][7] != ele[19][16];
    ele[19][7] != ele[19][17];
    ele[19][7] != ele[19][18];
    ele[19][7] != ele[19][19];
    ele[19][7] != ele[19][20];
    ele[19][7] != ele[19][21];
    ele[19][7] != ele[19][22];
    ele[19][7] != ele[19][23];
    ele[19][7] != ele[19][24];
    ele[19][7] != ele[19][8];
    ele[19][7] != ele[19][9];
    ele[19][7] != ele[20][7];
    ele[19][7] != ele[21][7];
    ele[19][7] != ele[22][7];
    ele[19][7] != ele[23][7];
    ele[19][7] != ele[24][7];
    ele[19][8] != ele[19][10];
    ele[19][8] != ele[19][11];
    ele[19][8] != ele[19][12];
    ele[19][8] != ele[19][13];
    ele[19][8] != ele[19][14];
    ele[19][8] != ele[19][15];
    ele[19][8] != ele[19][16];
    ele[19][8] != ele[19][17];
    ele[19][8] != ele[19][18];
    ele[19][8] != ele[19][19];
    ele[19][8] != ele[19][20];
    ele[19][8] != ele[19][21];
    ele[19][8] != ele[19][22];
    ele[19][8] != ele[19][23];
    ele[19][8] != ele[19][24];
    ele[19][8] != ele[19][9];
    ele[19][8] != ele[20][8];
    ele[19][8] != ele[21][8];
    ele[19][8] != ele[22][8];
    ele[19][8] != ele[23][8];
    ele[19][8] != ele[24][8];
    ele[19][9] != ele[19][10];
    ele[19][9] != ele[19][11];
    ele[19][9] != ele[19][12];
    ele[19][9] != ele[19][13];
    ele[19][9] != ele[19][14];
    ele[19][9] != ele[19][15];
    ele[19][9] != ele[19][16];
    ele[19][9] != ele[19][17];
    ele[19][9] != ele[19][18];
    ele[19][9] != ele[19][19];
    ele[19][9] != ele[19][20];
    ele[19][9] != ele[19][21];
    ele[19][9] != ele[19][22];
    ele[19][9] != ele[19][23];
    ele[19][9] != ele[19][24];
    ele[19][9] != ele[20][9];
    ele[19][9] != ele[21][9];
    ele[19][9] != ele[22][9];
    ele[19][9] != ele[23][9];
    ele[19][9] != ele[24][9];
    ele[2][0] != ele[10][0];
    ele[2][0] != ele[11][0];
    ele[2][0] != ele[12][0];
    ele[2][0] != ele[13][0];
    ele[2][0] != ele[14][0];
    ele[2][0] != ele[15][0];
    ele[2][0] != ele[16][0];
    ele[2][0] != ele[17][0];
    ele[2][0] != ele[18][0];
    ele[2][0] != ele[19][0];
    ele[2][0] != ele[2][1];
    ele[2][0] != ele[2][10];
    ele[2][0] != ele[2][11];
    ele[2][0] != ele[2][12];
    ele[2][0] != ele[2][13];
    ele[2][0] != ele[2][14];
    ele[2][0] != ele[2][15];
    ele[2][0] != ele[2][16];
    ele[2][0] != ele[2][17];
    ele[2][0] != ele[2][18];
    ele[2][0] != ele[2][19];
    ele[2][0] != ele[2][2];
    ele[2][0] != ele[2][20];
    ele[2][0] != ele[2][21];
    ele[2][0] != ele[2][22];
    ele[2][0] != ele[2][23];
    ele[2][0] != ele[2][24];
    ele[2][0] != ele[2][3];
    ele[2][0] != ele[2][4];
    ele[2][0] != ele[2][5];
    ele[2][0] != ele[2][6];
    ele[2][0] != ele[2][7];
    ele[2][0] != ele[2][8];
    ele[2][0] != ele[2][9];
    ele[2][0] != ele[20][0];
    ele[2][0] != ele[21][0];
    ele[2][0] != ele[22][0];
    ele[2][0] != ele[23][0];
    ele[2][0] != ele[24][0];
    ele[2][0] != ele[3][0];
    ele[2][0] != ele[3][1];
    ele[2][0] != ele[3][2];
    ele[2][0] != ele[3][3];
    ele[2][0] != ele[3][4];
    ele[2][0] != ele[4][0];
    ele[2][0] != ele[4][1];
    ele[2][0] != ele[4][2];
    ele[2][0] != ele[4][3];
    ele[2][0] != ele[4][4];
    ele[2][0] != ele[5][0];
    ele[2][0] != ele[6][0];
    ele[2][0] != ele[7][0];
    ele[2][0] != ele[8][0];
    ele[2][0] != ele[9][0];
    ele[2][1] != ele[10][1];
    ele[2][1] != ele[11][1];
    ele[2][1] != ele[12][1];
    ele[2][1] != ele[13][1];
    ele[2][1] != ele[14][1];
    ele[2][1] != ele[15][1];
    ele[2][1] != ele[16][1];
    ele[2][1] != ele[17][1];
    ele[2][1] != ele[18][1];
    ele[2][1] != ele[19][1];
    ele[2][1] != ele[2][10];
    ele[2][1] != ele[2][11];
    ele[2][1] != ele[2][12];
    ele[2][1] != ele[2][13];
    ele[2][1] != ele[2][14];
    ele[2][1] != ele[2][15];
    ele[2][1] != ele[2][16];
    ele[2][1] != ele[2][17];
    ele[2][1] != ele[2][18];
    ele[2][1] != ele[2][19];
    ele[2][1] != ele[2][2];
    ele[2][1] != ele[2][20];
    ele[2][1] != ele[2][21];
    ele[2][1] != ele[2][22];
    ele[2][1] != ele[2][23];
    ele[2][1] != ele[2][24];
    ele[2][1] != ele[2][3];
    ele[2][1] != ele[2][4];
    ele[2][1] != ele[2][5];
    ele[2][1] != ele[2][6];
    ele[2][1] != ele[2][7];
    ele[2][1] != ele[2][8];
    ele[2][1] != ele[2][9];
    ele[2][1] != ele[20][1];
    ele[2][1] != ele[21][1];
    ele[2][1] != ele[22][1];
    ele[2][1] != ele[23][1];
    ele[2][1] != ele[24][1];
    ele[2][1] != ele[3][0];
    ele[2][1] != ele[3][1];
    ele[2][1] != ele[3][2];
    ele[2][1] != ele[3][3];
    ele[2][1] != ele[3][4];
    ele[2][1] != ele[4][0];
    ele[2][1] != ele[4][1];
    ele[2][1] != ele[4][2];
    ele[2][1] != ele[4][3];
    ele[2][1] != ele[4][4];
    ele[2][1] != ele[5][1];
    ele[2][1] != ele[6][1];
    ele[2][1] != ele[7][1];
    ele[2][1] != ele[8][1];
    ele[2][1] != ele[9][1];
    ele[2][10] != ele[10][10];
    ele[2][10] != ele[11][10];
    ele[2][10] != ele[12][10];
    ele[2][10] != ele[13][10];
    ele[2][10] != ele[14][10];
    ele[2][10] != ele[15][10];
    ele[2][10] != ele[16][10];
    ele[2][10] != ele[17][10];
    ele[2][10] != ele[18][10];
    ele[2][10] != ele[19][10];
    ele[2][10] != ele[2][11];
    ele[2][10] != ele[2][12];
    ele[2][10] != ele[2][13];
    ele[2][10] != ele[2][14];
    ele[2][10] != ele[2][15];
    ele[2][10] != ele[2][16];
    ele[2][10] != ele[2][17];
    ele[2][10] != ele[2][18];
    ele[2][10] != ele[2][19];
    ele[2][10] != ele[2][20];
    ele[2][10] != ele[2][21];
    ele[2][10] != ele[2][22];
    ele[2][10] != ele[2][23];
    ele[2][10] != ele[2][24];
    ele[2][10] != ele[20][10];
    ele[2][10] != ele[21][10];
    ele[2][10] != ele[22][10];
    ele[2][10] != ele[23][10];
    ele[2][10] != ele[24][10];
    ele[2][10] != ele[3][10];
    ele[2][10] != ele[3][11];
    ele[2][10] != ele[3][12];
    ele[2][10] != ele[3][13];
    ele[2][10] != ele[3][14];
    ele[2][10] != ele[4][10];
    ele[2][10] != ele[4][11];
    ele[2][10] != ele[4][12];
    ele[2][10] != ele[4][13];
    ele[2][10] != ele[4][14];
    ele[2][10] != ele[5][10];
    ele[2][10] != ele[6][10];
    ele[2][10] != ele[7][10];
    ele[2][10] != ele[8][10];
    ele[2][10] != ele[9][10];
    ele[2][11] != ele[10][11];
    ele[2][11] != ele[11][11];
    ele[2][11] != ele[12][11];
    ele[2][11] != ele[13][11];
    ele[2][11] != ele[14][11];
    ele[2][11] != ele[15][11];
    ele[2][11] != ele[16][11];
    ele[2][11] != ele[17][11];
    ele[2][11] != ele[18][11];
    ele[2][11] != ele[19][11];
    ele[2][11] != ele[2][12];
    ele[2][11] != ele[2][13];
    ele[2][11] != ele[2][14];
    ele[2][11] != ele[2][15];
    ele[2][11] != ele[2][16];
    ele[2][11] != ele[2][17];
    ele[2][11] != ele[2][18];
    ele[2][11] != ele[2][19];
    ele[2][11] != ele[2][20];
    ele[2][11] != ele[2][21];
    ele[2][11] != ele[2][22];
    ele[2][11] != ele[2][23];
    ele[2][11] != ele[2][24];
    ele[2][11] != ele[20][11];
    ele[2][11] != ele[21][11];
    ele[2][11] != ele[22][11];
    ele[2][11] != ele[23][11];
    ele[2][11] != ele[24][11];
    ele[2][11] != ele[3][10];
    ele[2][11] != ele[3][11];
    ele[2][11] != ele[3][12];
    ele[2][11] != ele[3][13];
    ele[2][11] != ele[3][14];
    ele[2][11] != ele[4][10];
    ele[2][11] != ele[4][11];
    ele[2][11] != ele[4][12];
    ele[2][11] != ele[4][13];
    ele[2][11] != ele[4][14];
    ele[2][11] != ele[5][11];
    ele[2][11] != ele[6][11];
    ele[2][11] != ele[7][11];
    ele[2][11] != ele[8][11];
    ele[2][11] != ele[9][11];
    ele[2][12] != ele[10][12];
    ele[2][12] != ele[11][12];
    ele[2][12] != ele[12][12];
    ele[2][12] != ele[13][12];
    ele[2][12] != ele[14][12];
    ele[2][12] != ele[15][12];
    ele[2][12] != ele[16][12];
    ele[2][12] != ele[17][12];
    ele[2][12] != ele[18][12];
    ele[2][12] != ele[19][12];
    ele[2][12] != ele[2][13];
    ele[2][12] != ele[2][14];
    ele[2][12] != ele[2][15];
    ele[2][12] != ele[2][16];
    ele[2][12] != ele[2][17];
    ele[2][12] != ele[2][18];
    ele[2][12] != ele[2][19];
    ele[2][12] != ele[2][20];
    ele[2][12] != ele[2][21];
    ele[2][12] != ele[2][22];
    ele[2][12] != ele[2][23];
    ele[2][12] != ele[2][24];
    ele[2][12] != ele[20][12];
    ele[2][12] != ele[21][12];
    ele[2][12] != ele[22][12];
    ele[2][12] != ele[23][12];
    ele[2][12] != ele[24][12];
    ele[2][12] != ele[3][10];
    ele[2][12] != ele[3][11];
    ele[2][12] != ele[3][12];
    ele[2][12] != ele[3][13];
    ele[2][12] != ele[3][14];
    ele[2][12] != ele[4][10];
    ele[2][12] != ele[4][11];
    ele[2][12] != ele[4][12];
    ele[2][12] != ele[4][13];
    ele[2][12] != ele[4][14];
    ele[2][12] != ele[5][12];
    ele[2][12] != ele[6][12];
    ele[2][12] != ele[7][12];
    ele[2][12] != ele[8][12];
    ele[2][12] != ele[9][12];
    ele[2][13] != ele[10][13];
    ele[2][13] != ele[11][13];
    ele[2][13] != ele[12][13];
    ele[2][13] != ele[13][13];
    ele[2][13] != ele[14][13];
    ele[2][13] != ele[15][13];
    ele[2][13] != ele[16][13];
    ele[2][13] != ele[17][13];
    ele[2][13] != ele[18][13];
    ele[2][13] != ele[19][13];
    ele[2][13] != ele[2][14];
    ele[2][13] != ele[2][15];
    ele[2][13] != ele[2][16];
    ele[2][13] != ele[2][17];
    ele[2][13] != ele[2][18];
    ele[2][13] != ele[2][19];
    ele[2][13] != ele[2][20];
    ele[2][13] != ele[2][21];
    ele[2][13] != ele[2][22];
    ele[2][13] != ele[2][23];
    ele[2][13] != ele[2][24];
    ele[2][13] != ele[20][13];
    ele[2][13] != ele[21][13];
    ele[2][13] != ele[22][13];
    ele[2][13] != ele[23][13];
    ele[2][13] != ele[24][13];
    ele[2][13] != ele[3][10];
    ele[2][13] != ele[3][11];
    ele[2][13] != ele[3][12];
    ele[2][13] != ele[3][13];
    ele[2][13] != ele[3][14];
    ele[2][13] != ele[4][10];
    ele[2][13] != ele[4][11];
    ele[2][13] != ele[4][12];
    ele[2][13] != ele[4][13];
    ele[2][13] != ele[4][14];
    ele[2][13] != ele[5][13];
    ele[2][13] != ele[6][13];
    ele[2][13] != ele[7][13];
    ele[2][13] != ele[8][13];
    ele[2][13] != ele[9][13];
    ele[2][14] != ele[10][14];
    ele[2][14] != ele[11][14];
    ele[2][14] != ele[12][14];
    ele[2][14] != ele[13][14];
    ele[2][14] != ele[14][14];
    ele[2][14] != ele[15][14];
    ele[2][14] != ele[16][14];
    ele[2][14] != ele[17][14];
    ele[2][14] != ele[18][14];
    ele[2][14] != ele[19][14];
    ele[2][14] != ele[2][15];
    ele[2][14] != ele[2][16];
    ele[2][14] != ele[2][17];
    ele[2][14] != ele[2][18];
    ele[2][14] != ele[2][19];
    ele[2][14] != ele[2][20];
    ele[2][14] != ele[2][21];
    ele[2][14] != ele[2][22];
    ele[2][14] != ele[2][23];
    ele[2][14] != ele[2][24];
    ele[2][14] != ele[20][14];
    ele[2][14] != ele[21][14];
    ele[2][14] != ele[22][14];
    ele[2][14] != ele[23][14];
    ele[2][14] != ele[24][14];
    ele[2][14] != ele[3][10];
    ele[2][14] != ele[3][11];
    ele[2][14] != ele[3][12];
    ele[2][14] != ele[3][13];
    ele[2][14] != ele[3][14];
    ele[2][14] != ele[4][10];
    ele[2][14] != ele[4][11];
    ele[2][14] != ele[4][12];
    ele[2][14] != ele[4][13];
    ele[2][14] != ele[4][14];
    ele[2][14] != ele[5][14];
    ele[2][14] != ele[6][14];
    ele[2][14] != ele[7][14];
    ele[2][14] != ele[8][14];
    ele[2][14] != ele[9][14];
    ele[2][15] != ele[10][15];
    ele[2][15] != ele[11][15];
    ele[2][15] != ele[12][15];
    ele[2][15] != ele[13][15];
    ele[2][15] != ele[14][15];
    ele[2][15] != ele[15][15];
    ele[2][15] != ele[16][15];
    ele[2][15] != ele[17][15];
    ele[2][15] != ele[18][15];
    ele[2][15] != ele[19][15];
    ele[2][15] != ele[2][16];
    ele[2][15] != ele[2][17];
    ele[2][15] != ele[2][18];
    ele[2][15] != ele[2][19];
    ele[2][15] != ele[2][20];
    ele[2][15] != ele[2][21];
    ele[2][15] != ele[2][22];
    ele[2][15] != ele[2][23];
    ele[2][15] != ele[2][24];
    ele[2][15] != ele[20][15];
    ele[2][15] != ele[21][15];
    ele[2][15] != ele[22][15];
    ele[2][15] != ele[23][15];
    ele[2][15] != ele[24][15];
    ele[2][15] != ele[3][15];
    ele[2][15] != ele[3][16];
    ele[2][15] != ele[3][17];
    ele[2][15] != ele[3][18];
    ele[2][15] != ele[3][19];
    ele[2][15] != ele[4][15];
    ele[2][15] != ele[4][16];
    ele[2][15] != ele[4][17];
    ele[2][15] != ele[4][18];
    ele[2][15] != ele[4][19];
    ele[2][15] != ele[5][15];
    ele[2][15] != ele[6][15];
    ele[2][15] != ele[7][15];
    ele[2][15] != ele[8][15];
    ele[2][15] != ele[9][15];
    ele[2][16] != ele[10][16];
    ele[2][16] != ele[11][16];
    ele[2][16] != ele[12][16];
    ele[2][16] != ele[13][16];
    ele[2][16] != ele[14][16];
    ele[2][16] != ele[15][16];
    ele[2][16] != ele[16][16];
    ele[2][16] != ele[17][16];
    ele[2][16] != ele[18][16];
    ele[2][16] != ele[19][16];
    ele[2][16] != ele[2][17];
    ele[2][16] != ele[2][18];
    ele[2][16] != ele[2][19];
    ele[2][16] != ele[2][20];
    ele[2][16] != ele[2][21];
    ele[2][16] != ele[2][22];
    ele[2][16] != ele[2][23];
    ele[2][16] != ele[2][24];
    ele[2][16] != ele[20][16];
    ele[2][16] != ele[21][16];
    ele[2][16] != ele[22][16];
    ele[2][16] != ele[23][16];
    ele[2][16] != ele[24][16];
    ele[2][16] != ele[3][15];
    ele[2][16] != ele[3][16];
    ele[2][16] != ele[3][17];
    ele[2][16] != ele[3][18];
    ele[2][16] != ele[3][19];
    ele[2][16] != ele[4][15];
    ele[2][16] != ele[4][16];
    ele[2][16] != ele[4][17];
    ele[2][16] != ele[4][18];
    ele[2][16] != ele[4][19];
    ele[2][16] != ele[5][16];
    ele[2][16] != ele[6][16];
    ele[2][16] != ele[7][16];
    ele[2][16] != ele[8][16];
    ele[2][16] != ele[9][16];
    ele[2][17] != ele[10][17];
    ele[2][17] != ele[11][17];
    ele[2][17] != ele[12][17];
    ele[2][17] != ele[13][17];
    ele[2][17] != ele[14][17];
    ele[2][17] != ele[15][17];
    ele[2][17] != ele[16][17];
    ele[2][17] != ele[17][17];
    ele[2][17] != ele[18][17];
    ele[2][17] != ele[19][17];
    ele[2][17] != ele[2][18];
    ele[2][17] != ele[2][19];
    ele[2][17] != ele[2][20];
    ele[2][17] != ele[2][21];
    ele[2][17] != ele[2][22];
    ele[2][17] != ele[2][23];
    ele[2][17] != ele[2][24];
    ele[2][17] != ele[20][17];
    ele[2][17] != ele[21][17];
    ele[2][17] != ele[22][17];
    ele[2][17] != ele[23][17];
    ele[2][17] != ele[24][17];
    ele[2][17] != ele[3][15];
    ele[2][17] != ele[3][16];
    ele[2][17] != ele[3][17];
    ele[2][17] != ele[3][18];
    ele[2][17] != ele[3][19];
    ele[2][17] != ele[4][15];
    ele[2][17] != ele[4][16];
    ele[2][17] != ele[4][17];
    ele[2][17] != ele[4][18];
    ele[2][17] != ele[4][19];
    ele[2][17] != ele[5][17];
    ele[2][17] != ele[6][17];
    ele[2][17] != ele[7][17];
    ele[2][17] != ele[8][17];
    ele[2][17] != ele[9][17];
    ele[2][18] != ele[10][18];
    ele[2][18] != ele[11][18];
    ele[2][18] != ele[12][18];
    ele[2][18] != ele[13][18];
    ele[2][18] != ele[14][18];
    ele[2][18] != ele[15][18];
    ele[2][18] != ele[16][18];
    ele[2][18] != ele[17][18];
    ele[2][18] != ele[18][18];
    ele[2][18] != ele[19][18];
    ele[2][18] != ele[2][19];
    ele[2][18] != ele[2][20];
    ele[2][18] != ele[2][21];
    ele[2][18] != ele[2][22];
    ele[2][18] != ele[2][23];
    ele[2][18] != ele[2][24];
    ele[2][18] != ele[20][18];
    ele[2][18] != ele[21][18];
    ele[2][18] != ele[22][18];
    ele[2][18] != ele[23][18];
    ele[2][18] != ele[24][18];
    ele[2][18] != ele[3][15];
    ele[2][18] != ele[3][16];
    ele[2][18] != ele[3][17];
    ele[2][18] != ele[3][18];
    ele[2][18] != ele[3][19];
    ele[2][18] != ele[4][15];
    ele[2][18] != ele[4][16];
    ele[2][18] != ele[4][17];
    ele[2][18] != ele[4][18];
    ele[2][18] != ele[4][19];
    ele[2][18] != ele[5][18];
    ele[2][18] != ele[6][18];
    ele[2][18] != ele[7][18];
    ele[2][18] != ele[8][18];
    ele[2][18] != ele[9][18];
    ele[2][19] != ele[10][19];
    ele[2][19] != ele[11][19];
    ele[2][19] != ele[12][19];
    ele[2][19] != ele[13][19];
    ele[2][19] != ele[14][19];
    ele[2][19] != ele[15][19];
    ele[2][19] != ele[16][19];
    ele[2][19] != ele[17][19];
    ele[2][19] != ele[18][19];
    ele[2][19] != ele[19][19];
    ele[2][19] != ele[2][20];
    ele[2][19] != ele[2][21];
    ele[2][19] != ele[2][22];
    ele[2][19] != ele[2][23];
    ele[2][19] != ele[2][24];
    ele[2][19] != ele[20][19];
    ele[2][19] != ele[21][19];
    ele[2][19] != ele[22][19];
    ele[2][19] != ele[23][19];
    ele[2][19] != ele[24][19];
    ele[2][19] != ele[3][15];
    ele[2][19] != ele[3][16];
    ele[2][19] != ele[3][17];
    ele[2][19] != ele[3][18];
    ele[2][19] != ele[3][19];
    ele[2][19] != ele[4][15];
    ele[2][19] != ele[4][16];
    ele[2][19] != ele[4][17];
    ele[2][19] != ele[4][18];
    ele[2][19] != ele[4][19];
    ele[2][19] != ele[5][19];
    ele[2][19] != ele[6][19];
    ele[2][19] != ele[7][19];
    ele[2][19] != ele[8][19];
    ele[2][19] != ele[9][19];
    ele[2][2] != ele[10][2];
    ele[2][2] != ele[11][2];
    ele[2][2] != ele[12][2];
    ele[2][2] != ele[13][2];
    ele[2][2] != ele[14][2];
    ele[2][2] != ele[15][2];
    ele[2][2] != ele[16][2];
    ele[2][2] != ele[17][2];
    ele[2][2] != ele[18][2];
    ele[2][2] != ele[19][2];
    ele[2][2] != ele[2][10];
    ele[2][2] != ele[2][11];
    ele[2][2] != ele[2][12];
    ele[2][2] != ele[2][13];
    ele[2][2] != ele[2][14];
    ele[2][2] != ele[2][15];
    ele[2][2] != ele[2][16];
    ele[2][2] != ele[2][17];
    ele[2][2] != ele[2][18];
    ele[2][2] != ele[2][19];
    ele[2][2] != ele[2][20];
    ele[2][2] != ele[2][21];
    ele[2][2] != ele[2][22];
    ele[2][2] != ele[2][23];
    ele[2][2] != ele[2][24];
    ele[2][2] != ele[2][3];
    ele[2][2] != ele[2][4];
    ele[2][2] != ele[2][5];
    ele[2][2] != ele[2][6];
    ele[2][2] != ele[2][7];
    ele[2][2] != ele[2][8];
    ele[2][2] != ele[2][9];
    ele[2][2] != ele[20][2];
    ele[2][2] != ele[21][2];
    ele[2][2] != ele[22][2];
    ele[2][2] != ele[23][2];
    ele[2][2] != ele[24][2];
    ele[2][2] != ele[3][0];
    ele[2][2] != ele[3][1];
    ele[2][2] != ele[3][2];
    ele[2][2] != ele[3][3];
    ele[2][2] != ele[3][4];
    ele[2][2] != ele[4][0];
    ele[2][2] != ele[4][1];
    ele[2][2] != ele[4][2];
    ele[2][2] != ele[4][3];
    ele[2][2] != ele[4][4];
    ele[2][2] != ele[5][2];
    ele[2][2] != ele[6][2];
    ele[2][2] != ele[7][2];
    ele[2][2] != ele[8][2];
    ele[2][2] != ele[9][2];
    ele[2][20] != ele[10][20];
    ele[2][20] != ele[11][20];
    ele[2][20] != ele[12][20];
    ele[2][20] != ele[13][20];
    ele[2][20] != ele[14][20];
    ele[2][20] != ele[15][20];
    ele[2][20] != ele[16][20];
    ele[2][20] != ele[17][20];
    ele[2][20] != ele[18][20];
    ele[2][20] != ele[19][20];
    ele[2][20] != ele[2][21];
    ele[2][20] != ele[2][22];
    ele[2][20] != ele[2][23];
    ele[2][20] != ele[2][24];
    ele[2][20] != ele[20][20];
    ele[2][20] != ele[21][20];
    ele[2][20] != ele[22][20];
    ele[2][20] != ele[23][20];
    ele[2][20] != ele[24][20];
    ele[2][20] != ele[3][20];
    ele[2][20] != ele[3][21];
    ele[2][20] != ele[3][22];
    ele[2][20] != ele[3][23];
    ele[2][20] != ele[3][24];
    ele[2][20] != ele[4][20];
    ele[2][20] != ele[4][21];
    ele[2][20] != ele[4][22];
    ele[2][20] != ele[4][23];
    ele[2][20] != ele[4][24];
    ele[2][20] != ele[5][20];
    ele[2][20] != ele[6][20];
    ele[2][20] != ele[7][20];
    ele[2][20] != ele[8][20];
    ele[2][20] != ele[9][20];
    ele[2][21] != ele[10][21];
    ele[2][21] != ele[11][21];
    ele[2][21] != ele[12][21];
    ele[2][21] != ele[13][21];
    ele[2][21] != ele[14][21];
    ele[2][21] != ele[15][21];
    ele[2][21] != ele[16][21];
    ele[2][21] != ele[17][21];
    ele[2][21] != ele[18][21];
    ele[2][21] != ele[19][21];
    ele[2][21] != ele[2][22];
    ele[2][21] != ele[2][23];
    ele[2][21] != ele[2][24];
    ele[2][21] != ele[20][21];
    ele[2][21] != ele[21][21];
    ele[2][21] != ele[22][21];
    ele[2][21] != ele[23][21];
    ele[2][21] != ele[24][21];
    ele[2][21] != ele[3][20];
    ele[2][21] != ele[3][21];
    ele[2][21] != ele[3][22];
    ele[2][21] != ele[3][23];
    ele[2][21] != ele[3][24];
    ele[2][21] != ele[4][20];
    ele[2][21] != ele[4][21];
    ele[2][21] != ele[4][22];
    ele[2][21] != ele[4][23];
    ele[2][21] != ele[4][24];
    ele[2][21] != ele[5][21];
    ele[2][21] != ele[6][21];
    ele[2][21] != ele[7][21];
    ele[2][21] != ele[8][21];
    ele[2][21] != ele[9][21];
    ele[2][22] != ele[10][22];
    ele[2][22] != ele[11][22];
    ele[2][22] != ele[12][22];
    ele[2][22] != ele[13][22];
    ele[2][22] != ele[14][22];
    ele[2][22] != ele[15][22];
    ele[2][22] != ele[16][22];
    ele[2][22] != ele[17][22];
    ele[2][22] != ele[18][22];
    ele[2][22] != ele[19][22];
    ele[2][22] != ele[2][23];
    ele[2][22] != ele[2][24];
    ele[2][22] != ele[20][22];
    ele[2][22] != ele[21][22];
    ele[2][22] != ele[22][22];
    ele[2][22] != ele[23][22];
    ele[2][22] != ele[24][22];
    ele[2][22] != ele[3][20];
    ele[2][22] != ele[3][21];
    ele[2][22] != ele[3][22];
    ele[2][22] != ele[3][23];
    ele[2][22] != ele[3][24];
    ele[2][22] != ele[4][20];
    ele[2][22] != ele[4][21];
    ele[2][22] != ele[4][22];
    ele[2][22] != ele[4][23];
    ele[2][22] != ele[4][24];
    ele[2][22] != ele[5][22];
    ele[2][22] != ele[6][22];
    ele[2][22] != ele[7][22];
    ele[2][22] != ele[8][22];
    ele[2][22] != ele[9][22];
    ele[2][23] != ele[10][23];
    ele[2][23] != ele[11][23];
    ele[2][23] != ele[12][23];
    ele[2][23] != ele[13][23];
    ele[2][23] != ele[14][23];
    ele[2][23] != ele[15][23];
    ele[2][23] != ele[16][23];
    ele[2][23] != ele[17][23];
    ele[2][23] != ele[18][23];
    ele[2][23] != ele[19][23];
    ele[2][23] != ele[2][24];
    ele[2][23] != ele[20][23];
    ele[2][23] != ele[21][23];
    ele[2][23] != ele[22][23];
    ele[2][23] != ele[23][23];
    ele[2][23] != ele[24][23];
    ele[2][23] != ele[3][20];
    ele[2][23] != ele[3][21];
    ele[2][23] != ele[3][22];
    ele[2][23] != ele[3][23];
    ele[2][23] != ele[3][24];
    ele[2][23] != ele[4][20];
    ele[2][23] != ele[4][21];
    ele[2][23] != ele[4][22];
    ele[2][23] != ele[4][23];
    ele[2][23] != ele[4][24];
    ele[2][23] != ele[5][23];
    ele[2][23] != ele[6][23];
    ele[2][23] != ele[7][23];
    ele[2][23] != ele[8][23];
    ele[2][23] != ele[9][23];
    ele[2][24] != ele[10][24];
    ele[2][24] != ele[11][24];
    ele[2][24] != ele[12][24];
    ele[2][24] != ele[13][24];
    ele[2][24] != ele[14][24];
    ele[2][24] != ele[15][24];
    ele[2][24] != ele[16][24];
    ele[2][24] != ele[17][24];
    ele[2][24] != ele[18][24];
    ele[2][24] != ele[19][24];
    ele[2][24] != ele[20][24];
    ele[2][24] != ele[21][24];
    ele[2][24] != ele[22][24];
    ele[2][24] != ele[23][24];
    ele[2][24] != ele[24][24];
    ele[2][24] != ele[3][20];
    ele[2][24] != ele[3][21];
    ele[2][24] != ele[3][22];
    ele[2][24] != ele[3][23];
    ele[2][24] != ele[3][24];
    ele[2][24] != ele[4][20];
    ele[2][24] != ele[4][21];
    ele[2][24] != ele[4][22];
    ele[2][24] != ele[4][23];
    ele[2][24] != ele[4][24];
    ele[2][24] != ele[5][24];
    ele[2][24] != ele[6][24];
    ele[2][24] != ele[7][24];
    ele[2][24] != ele[8][24];
    ele[2][24] != ele[9][24];
    ele[2][3] != ele[10][3];
    ele[2][3] != ele[11][3];
    ele[2][3] != ele[12][3];
    ele[2][3] != ele[13][3];
    ele[2][3] != ele[14][3];
    ele[2][3] != ele[15][3];
    ele[2][3] != ele[16][3];
    ele[2][3] != ele[17][3];
    ele[2][3] != ele[18][3];
    ele[2][3] != ele[19][3];
    ele[2][3] != ele[2][10];
    ele[2][3] != ele[2][11];
    ele[2][3] != ele[2][12];
    ele[2][3] != ele[2][13];
    ele[2][3] != ele[2][14];
    ele[2][3] != ele[2][15];
    ele[2][3] != ele[2][16];
    ele[2][3] != ele[2][17];
    ele[2][3] != ele[2][18];
    ele[2][3] != ele[2][19];
    ele[2][3] != ele[2][20];
    ele[2][3] != ele[2][21];
    ele[2][3] != ele[2][22];
    ele[2][3] != ele[2][23];
    ele[2][3] != ele[2][24];
    ele[2][3] != ele[2][4];
    ele[2][3] != ele[2][5];
    ele[2][3] != ele[2][6];
    ele[2][3] != ele[2][7];
    ele[2][3] != ele[2][8];
    ele[2][3] != ele[2][9];
    ele[2][3] != ele[20][3];
    ele[2][3] != ele[21][3];
    ele[2][3] != ele[22][3];
    ele[2][3] != ele[23][3];
    ele[2][3] != ele[24][3];
    ele[2][3] != ele[3][0];
    ele[2][3] != ele[3][1];
    ele[2][3] != ele[3][2];
    ele[2][3] != ele[3][3];
    ele[2][3] != ele[3][4];
    ele[2][3] != ele[4][0];
    ele[2][3] != ele[4][1];
    ele[2][3] != ele[4][2];
    ele[2][3] != ele[4][3];
    ele[2][3] != ele[4][4];
    ele[2][3] != ele[5][3];
    ele[2][3] != ele[6][3];
    ele[2][3] != ele[7][3];
    ele[2][3] != ele[8][3];
    ele[2][3] != ele[9][3];
    ele[2][4] != ele[10][4];
    ele[2][4] != ele[11][4];
    ele[2][4] != ele[12][4];
    ele[2][4] != ele[13][4];
    ele[2][4] != ele[14][4];
    ele[2][4] != ele[15][4];
    ele[2][4] != ele[16][4];
    ele[2][4] != ele[17][4];
    ele[2][4] != ele[18][4];
    ele[2][4] != ele[19][4];
    ele[2][4] != ele[2][10];
    ele[2][4] != ele[2][11];
    ele[2][4] != ele[2][12];
    ele[2][4] != ele[2][13];
    ele[2][4] != ele[2][14];
    ele[2][4] != ele[2][15];
    ele[2][4] != ele[2][16];
    ele[2][4] != ele[2][17];
    ele[2][4] != ele[2][18];
    ele[2][4] != ele[2][19];
    ele[2][4] != ele[2][20];
    ele[2][4] != ele[2][21];
    ele[2][4] != ele[2][22];
    ele[2][4] != ele[2][23];
    ele[2][4] != ele[2][24];
    ele[2][4] != ele[2][5];
    ele[2][4] != ele[2][6];
    ele[2][4] != ele[2][7];
    ele[2][4] != ele[2][8];
    ele[2][4] != ele[2][9];
    ele[2][4] != ele[20][4];
    ele[2][4] != ele[21][4];
    ele[2][4] != ele[22][4];
    ele[2][4] != ele[23][4];
    ele[2][4] != ele[24][4];
    ele[2][4] != ele[3][0];
    ele[2][4] != ele[3][1];
    ele[2][4] != ele[3][2];
    ele[2][4] != ele[3][3];
    ele[2][4] != ele[3][4];
    ele[2][4] != ele[4][0];
    ele[2][4] != ele[4][1];
    ele[2][4] != ele[4][2];
    ele[2][4] != ele[4][3];
    ele[2][4] != ele[4][4];
    ele[2][4] != ele[5][4];
    ele[2][4] != ele[6][4];
    ele[2][4] != ele[7][4];
    ele[2][4] != ele[8][4];
    ele[2][4] != ele[9][4];
    ele[2][5] != ele[10][5];
    ele[2][5] != ele[11][5];
    ele[2][5] != ele[12][5];
    ele[2][5] != ele[13][5];
    ele[2][5] != ele[14][5];
    ele[2][5] != ele[15][5];
    ele[2][5] != ele[16][5];
    ele[2][5] != ele[17][5];
    ele[2][5] != ele[18][5];
    ele[2][5] != ele[19][5];
    ele[2][5] != ele[2][10];
    ele[2][5] != ele[2][11];
    ele[2][5] != ele[2][12];
    ele[2][5] != ele[2][13];
    ele[2][5] != ele[2][14];
    ele[2][5] != ele[2][15];
    ele[2][5] != ele[2][16];
    ele[2][5] != ele[2][17];
    ele[2][5] != ele[2][18];
    ele[2][5] != ele[2][19];
    ele[2][5] != ele[2][20];
    ele[2][5] != ele[2][21];
    ele[2][5] != ele[2][22];
    ele[2][5] != ele[2][23];
    ele[2][5] != ele[2][24];
    ele[2][5] != ele[2][6];
    ele[2][5] != ele[2][7];
    ele[2][5] != ele[2][8];
    ele[2][5] != ele[2][9];
    ele[2][5] != ele[20][5];
    ele[2][5] != ele[21][5];
    ele[2][5] != ele[22][5];
    ele[2][5] != ele[23][5];
    ele[2][5] != ele[24][5];
    ele[2][5] != ele[3][5];
    ele[2][5] != ele[3][6];
    ele[2][5] != ele[3][7];
    ele[2][5] != ele[3][8];
    ele[2][5] != ele[3][9];
    ele[2][5] != ele[4][5];
    ele[2][5] != ele[4][6];
    ele[2][5] != ele[4][7];
    ele[2][5] != ele[4][8];
    ele[2][5] != ele[4][9];
    ele[2][5] != ele[5][5];
    ele[2][5] != ele[6][5];
    ele[2][5] != ele[7][5];
    ele[2][5] != ele[8][5];
    ele[2][5] != ele[9][5];
    ele[2][6] != ele[10][6];
    ele[2][6] != ele[11][6];
    ele[2][6] != ele[12][6];
    ele[2][6] != ele[13][6];
    ele[2][6] != ele[14][6];
    ele[2][6] != ele[15][6];
    ele[2][6] != ele[16][6];
    ele[2][6] != ele[17][6];
    ele[2][6] != ele[18][6];
    ele[2][6] != ele[19][6];
    ele[2][6] != ele[2][10];
    ele[2][6] != ele[2][11];
    ele[2][6] != ele[2][12];
    ele[2][6] != ele[2][13];
    ele[2][6] != ele[2][14];
    ele[2][6] != ele[2][15];
    ele[2][6] != ele[2][16];
    ele[2][6] != ele[2][17];
    ele[2][6] != ele[2][18];
    ele[2][6] != ele[2][19];
    ele[2][6] != ele[2][20];
    ele[2][6] != ele[2][21];
    ele[2][6] != ele[2][22];
    ele[2][6] != ele[2][23];
    ele[2][6] != ele[2][24];
    ele[2][6] != ele[2][7];
    ele[2][6] != ele[2][8];
    ele[2][6] != ele[2][9];
    ele[2][6] != ele[20][6];
    ele[2][6] != ele[21][6];
    ele[2][6] != ele[22][6];
    ele[2][6] != ele[23][6];
    ele[2][6] != ele[24][6];
    ele[2][6] != ele[3][5];
    ele[2][6] != ele[3][6];
    ele[2][6] != ele[3][7];
    ele[2][6] != ele[3][8];
    ele[2][6] != ele[3][9];
    ele[2][6] != ele[4][5];
    ele[2][6] != ele[4][6];
    ele[2][6] != ele[4][7];
    ele[2][6] != ele[4][8];
    ele[2][6] != ele[4][9];
    ele[2][6] != ele[5][6];
    ele[2][6] != ele[6][6];
    ele[2][6] != ele[7][6];
    ele[2][6] != ele[8][6];
    ele[2][6] != ele[9][6];
    ele[2][7] != ele[10][7];
    ele[2][7] != ele[11][7];
    ele[2][7] != ele[12][7];
    ele[2][7] != ele[13][7];
    ele[2][7] != ele[14][7];
    ele[2][7] != ele[15][7];
    ele[2][7] != ele[16][7];
    ele[2][7] != ele[17][7];
    ele[2][7] != ele[18][7];
    ele[2][7] != ele[19][7];
    ele[2][7] != ele[2][10];
    ele[2][7] != ele[2][11];
    ele[2][7] != ele[2][12];
    ele[2][7] != ele[2][13];
    ele[2][7] != ele[2][14];
    ele[2][7] != ele[2][15];
    ele[2][7] != ele[2][16];
    ele[2][7] != ele[2][17];
    ele[2][7] != ele[2][18];
    ele[2][7] != ele[2][19];
    ele[2][7] != ele[2][20];
    ele[2][7] != ele[2][21];
    ele[2][7] != ele[2][22];
    ele[2][7] != ele[2][23];
    ele[2][7] != ele[2][24];
    ele[2][7] != ele[2][8];
    ele[2][7] != ele[2][9];
    ele[2][7] != ele[20][7];
    ele[2][7] != ele[21][7];
    ele[2][7] != ele[22][7];
    ele[2][7] != ele[23][7];
    ele[2][7] != ele[24][7];
    ele[2][7] != ele[3][5];
    ele[2][7] != ele[3][6];
    ele[2][7] != ele[3][7];
    ele[2][7] != ele[3][8];
    ele[2][7] != ele[3][9];
    ele[2][7] != ele[4][5];
    ele[2][7] != ele[4][6];
    ele[2][7] != ele[4][7];
    ele[2][7] != ele[4][8];
    ele[2][7] != ele[4][9];
    ele[2][7] != ele[5][7];
    ele[2][7] != ele[6][7];
    ele[2][7] != ele[7][7];
    ele[2][7] != ele[8][7];
    ele[2][7] != ele[9][7];
    ele[2][8] != ele[10][8];
    ele[2][8] != ele[11][8];
    ele[2][8] != ele[12][8];
    ele[2][8] != ele[13][8];
    ele[2][8] != ele[14][8];
    ele[2][8] != ele[15][8];
    ele[2][8] != ele[16][8];
    ele[2][8] != ele[17][8];
    ele[2][8] != ele[18][8];
    ele[2][8] != ele[19][8];
    ele[2][8] != ele[2][10];
    ele[2][8] != ele[2][11];
    ele[2][8] != ele[2][12];
    ele[2][8] != ele[2][13];
    ele[2][8] != ele[2][14];
    ele[2][8] != ele[2][15];
    ele[2][8] != ele[2][16];
    ele[2][8] != ele[2][17];
    ele[2][8] != ele[2][18];
    ele[2][8] != ele[2][19];
    ele[2][8] != ele[2][20];
    ele[2][8] != ele[2][21];
    ele[2][8] != ele[2][22];
    ele[2][8] != ele[2][23];
    ele[2][8] != ele[2][24];
    ele[2][8] != ele[2][9];
    ele[2][8] != ele[20][8];
    ele[2][8] != ele[21][8];
    ele[2][8] != ele[22][8];
    ele[2][8] != ele[23][8];
    ele[2][8] != ele[24][8];
    ele[2][8] != ele[3][5];
    ele[2][8] != ele[3][6];
    ele[2][8] != ele[3][7];
    ele[2][8] != ele[3][8];
    ele[2][8] != ele[3][9];
    ele[2][8] != ele[4][5];
    ele[2][8] != ele[4][6];
    ele[2][8] != ele[4][7];
    ele[2][8] != ele[4][8];
    ele[2][8] != ele[4][9];
    ele[2][8] != ele[5][8];
    ele[2][8] != ele[6][8];
    ele[2][8] != ele[7][8];
    ele[2][8] != ele[8][8];
    ele[2][8] != ele[9][8];
    ele[2][9] != ele[10][9];
    ele[2][9] != ele[11][9];
    ele[2][9] != ele[12][9];
    ele[2][9] != ele[13][9];
    ele[2][9] != ele[14][9];
    ele[2][9] != ele[15][9];
    ele[2][9] != ele[16][9];
    ele[2][9] != ele[17][9];
    ele[2][9] != ele[18][9];
    ele[2][9] != ele[19][9];
    ele[2][9] != ele[2][10];
    ele[2][9] != ele[2][11];
    ele[2][9] != ele[2][12];
    ele[2][9] != ele[2][13];
    ele[2][9] != ele[2][14];
    ele[2][9] != ele[2][15];
    ele[2][9] != ele[2][16];
    ele[2][9] != ele[2][17];
    ele[2][9] != ele[2][18];
    ele[2][9] != ele[2][19];
    ele[2][9] != ele[2][20];
    ele[2][9] != ele[2][21];
    ele[2][9] != ele[2][22];
    ele[2][9] != ele[2][23];
    ele[2][9] != ele[2][24];
    ele[2][9] != ele[20][9];
    ele[2][9] != ele[21][9];
    ele[2][9] != ele[22][9];
    ele[2][9] != ele[23][9];
    ele[2][9] != ele[24][9];
    ele[2][9] != ele[3][5];
    ele[2][9] != ele[3][6];
    ele[2][9] != ele[3][7];
    ele[2][9] != ele[3][8];
    ele[2][9] != ele[3][9];
    ele[2][9] != ele[4][5];
    ele[2][9] != ele[4][6];
    ele[2][9] != ele[4][7];
    ele[2][9] != ele[4][8];
    ele[2][9] != ele[4][9];
    ele[2][9] != ele[5][9];
    ele[2][9] != ele[6][9];
    ele[2][9] != ele[7][9];
    ele[2][9] != ele[8][9];
    ele[2][9] != ele[9][9];
    ele[20][0] != ele[20][1];
    ele[20][0] != ele[20][10];
    ele[20][0] != ele[20][11];
    ele[20][0] != ele[20][12];
    ele[20][0] != ele[20][13];
    ele[20][0] != ele[20][14];
    ele[20][0] != ele[20][15];
    ele[20][0] != ele[20][16];
    ele[20][0] != ele[20][17];
    ele[20][0] != ele[20][18];
    ele[20][0] != ele[20][19];
    ele[20][0] != ele[20][2];
    ele[20][0] != ele[20][20];
    ele[20][0] != ele[20][21];
    ele[20][0] != ele[20][22];
    ele[20][0] != ele[20][23];
    ele[20][0] != ele[20][24];
    ele[20][0] != ele[20][3];
    ele[20][0] != ele[20][4];
    ele[20][0] != ele[20][5];
    ele[20][0] != ele[20][6];
    ele[20][0] != ele[20][7];
    ele[20][0] != ele[20][8];
    ele[20][0] != ele[20][9];
    ele[20][0] != ele[21][0];
    ele[20][0] != ele[21][1];
    ele[20][0] != ele[21][2];
    ele[20][0] != ele[21][3];
    ele[20][0] != ele[21][4];
    ele[20][0] != ele[22][0];
    ele[20][0] != ele[22][1];
    ele[20][0] != ele[22][2];
    ele[20][0] != ele[22][3];
    ele[20][0] != ele[22][4];
    ele[20][0] != ele[23][0];
    ele[20][0] != ele[23][1];
    ele[20][0] != ele[23][2];
    ele[20][0] != ele[23][3];
    ele[20][0] != ele[23][4];
    ele[20][0] != ele[24][0];
    ele[20][0] != ele[24][1];
    ele[20][0] != ele[24][2];
    ele[20][0] != ele[24][3];
    ele[20][0] != ele[24][4];
    ele[20][1] != ele[20][10];
    ele[20][1] != ele[20][11];
    ele[20][1] != ele[20][12];
    ele[20][1] != ele[20][13];
    ele[20][1] != ele[20][14];
    ele[20][1] != ele[20][15];
    ele[20][1] != ele[20][16];
    ele[20][1] != ele[20][17];
    ele[20][1] != ele[20][18];
    ele[20][1] != ele[20][19];
    ele[20][1] != ele[20][2];
    ele[20][1] != ele[20][20];
    ele[20][1] != ele[20][21];
    ele[20][1] != ele[20][22];
    ele[20][1] != ele[20][23];
    ele[20][1] != ele[20][24];
    ele[20][1] != ele[20][3];
    ele[20][1] != ele[20][4];
    ele[20][1] != ele[20][5];
    ele[20][1] != ele[20][6];
    ele[20][1] != ele[20][7];
    ele[20][1] != ele[20][8];
    ele[20][1] != ele[20][9];
    ele[20][1] != ele[21][0];
    ele[20][1] != ele[21][1];
    ele[20][1] != ele[21][2];
    ele[20][1] != ele[21][3];
    ele[20][1] != ele[21][4];
    ele[20][1] != ele[22][0];
    ele[20][1] != ele[22][1];
    ele[20][1] != ele[22][2];
    ele[20][1] != ele[22][3];
    ele[20][1] != ele[22][4];
    ele[20][1] != ele[23][0];
    ele[20][1] != ele[23][1];
    ele[20][1] != ele[23][2];
    ele[20][1] != ele[23][3];
    ele[20][1] != ele[23][4];
    ele[20][1] != ele[24][0];
    ele[20][1] != ele[24][1];
    ele[20][1] != ele[24][2];
    ele[20][1] != ele[24][3];
    ele[20][1] != ele[24][4];
    ele[20][10] != ele[20][11];
    ele[20][10] != ele[20][12];
    ele[20][10] != ele[20][13];
    ele[20][10] != ele[20][14];
    ele[20][10] != ele[20][15];
    ele[20][10] != ele[20][16];
    ele[20][10] != ele[20][17];
    ele[20][10] != ele[20][18];
    ele[20][10] != ele[20][19];
    ele[20][10] != ele[20][20];
    ele[20][10] != ele[20][21];
    ele[20][10] != ele[20][22];
    ele[20][10] != ele[20][23];
    ele[20][10] != ele[20][24];
    ele[20][10] != ele[21][10];
    ele[20][10] != ele[21][11];
    ele[20][10] != ele[21][12];
    ele[20][10] != ele[21][13];
    ele[20][10] != ele[21][14];
    ele[20][10] != ele[22][10];
    ele[20][10] != ele[22][11];
    ele[20][10] != ele[22][12];
    ele[20][10] != ele[22][13];
    ele[20][10] != ele[22][14];
    ele[20][10] != ele[23][10];
    ele[20][10] != ele[23][11];
    ele[20][10] != ele[23][12];
    ele[20][10] != ele[23][13];
    ele[20][10] != ele[23][14];
    ele[20][10] != ele[24][10];
    ele[20][10] != ele[24][11];
    ele[20][10] != ele[24][12];
    ele[20][10] != ele[24][13];
    ele[20][10] != ele[24][14];
    ele[20][11] != ele[20][12];
    ele[20][11] != ele[20][13];
    ele[20][11] != ele[20][14];
    ele[20][11] != ele[20][15];
    ele[20][11] != ele[20][16];
    ele[20][11] != ele[20][17];
    ele[20][11] != ele[20][18];
    ele[20][11] != ele[20][19];
    ele[20][11] != ele[20][20];
    ele[20][11] != ele[20][21];
    ele[20][11] != ele[20][22];
    ele[20][11] != ele[20][23];
    ele[20][11] != ele[20][24];
    ele[20][11] != ele[21][10];
    ele[20][11] != ele[21][11];
    ele[20][11] != ele[21][12];
    ele[20][11] != ele[21][13];
    ele[20][11] != ele[21][14];
    ele[20][11] != ele[22][10];
    ele[20][11] != ele[22][11];
    ele[20][11] != ele[22][12];
    ele[20][11] != ele[22][13];
    ele[20][11] != ele[22][14];
    ele[20][11] != ele[23][10];
    ele[20][11] != ele[23][11];
    ele[20][11] != ele[23][12];
    ele[20][11] != ele[23][13];
    ele[20][11] != ele[23][14];
    ele[20][11] != ele[24][10];
    ele[20][11] != ele[24][11];
    ele[20][11] != ele[24][12];
    ele[20][11] != ele[24][13];
    ele[20][11] != ele[24][14];
    ele[20][12] != ele[20][13];
    ele[20][12] != ele[20][14];
    ele[20][12] != ele[20][15];
    ele[20][12] != ele[20][16];
    ele[20][12] != ele[20][17];
    ele[20][12] != ele[20][18];
    ele[20][12] != ele[20][19];
    ele[20][12] != ele[20][20];
    ele[20][12] != ele[20][21];
    ele[20][12] != ele[20][22];
    ele[20][12] != ele[20][23];
    ele[20][12] != ele[20][24];
    ele[20][12] != ele[21][10];
    ele[20][12] != ele[21][11];
    ele[20][12] != ele[21][12];
    ele[20][12] != ele[21][13];
    ele[20][12] != ele[21][14];
    ele[20][12] != ele[22][10];
    ele[20][12] != ele[22][11];
    ele[20][12] != ele[22][12];
    ele[20][12] != ele[22][13];
    ele[20][12] != ele[22][14];
    ele[20][12] != ele[23][10];
    ele[20][12] != ele[23][11];
    ele[20][12] != ele[23][12];
    ele[20][12] != ele[23][13];
    ele[20][12] != ele[23][14];
    ele[20][12] != ele[24][10];
    ele[20][12] != ele[24][11];
    ele[20][12] != ele[24][12];
    ele[20][12] != ele[24][13];
    ele[20][12] != ele[24][14];
    ele[20][13] != ele[20][14];
    ele[20][13] != ele[20][15];
    ele[20][13] != ele[20][16];
    ele[20][13] != ele[20][17];
    ele[20][13] != ele[20][18];
    ele[20][13] != ele[20][19];
    ele[20][13] != ele[20][20];
    ele[20][13] != ele[20][21];
    ele[20][13] != ele[20][22];
    ele[20][13] != ele[20][23];
    ele[20][13] != ele[20][24];
    ele[20][13] != ele[21][10];
    ele[20][13] != ele[21][11];
    ele[20][13] != ele[21][12];
    ele[20][13] != ele[21][13];
    ele[20][13] != ele[21][14];
    ele[20][13] != ele[22][10];
    ele[20][13] != ele[22][11];
    ele[20][13] != ele[22][12];
    ele[20][13] != ele[22][13];
    ele[20][13] != ele[22][14];
    ele[20][13] != ele[23][10];
    ele[20][13] != ele[23][11];
    ele[20][13] != ele[23][12];
    ele[20][13] != ele[23][13];
    ele[20][13] != ele[23][14];
    ele[20][13] != ele[24][10];
    ele[20][13] != ele[24][11];
    ele[20][13] != ele[24][12];
    ele[20][13] != ele[24][13];
    ele[20][13] != ele[24][14];
    ele[20][14] != ele[20][15];
    ele[20][14] != ele[20][16];
    ele[20][14] != ele[20][17];
    ele[20][14] != ele[20][18];
    ele[20][14] != ele[20][19];
    ele[20][14] != ele[20][20];
    ele[20][14] != ele[20][21];
    ele[20][14] != ele[20][22];
    ele[20][14] != ele[20][23];
    ele[20][14] != ele[20][24];
    ele[20][14] != ele[21][10];
    ele[20][14] != ele[21][11];
    ele[20][14] != ele[21][12];
    ele[20][14] != ele[21][13];
    ele[20][14] != ele[21][14];
    ele[20][14] != ele[22][10];
    ele[20][14] != ele[22][11];
    ele[20][14] != ele[22][12];
    ele[20][14] != ele[22][13];
    ele[20][14] != ele[22][14];
    ele[20][14] != ele[23][10];
    ele[20][14] != ele[23][11];
    ele[20][14] != ele[23][12];
    ele[20][14] != ele[23][13];
    ele[20][14] != ele[23][14];
    ele[20][14] != ele[24][10];
    ele[20][14] != ele[24][11];
    ele[20][14] != ele[24][12];
    ele[20][14] != ele[24][13];
    ele[20][14] != ele[24][14];
    ele[20][15] != ele[20][16];
    ele[20][15] != ele[20][17];
    ele[20][15] != ele[20][18];
    ele[20][15] != ele[20][19];
    ele[20][15] != ele[20][20];
    ele[20][15] != ele[20][21];
    ele[20][15] != ele[20][22];
    ele[20][15] != ele[20][23];
    ele[20][15] != ele[20][24];
    ele[20][15] != ele[21][15];
    ele[20][15] != ele[21][16];
    ele[20][15] != ele[21][17];
    ele[20][15] != ele[21][18];
    ele[20][15] != ele[21][19];
    ele[20][15] != ele[22][15];
    ele[20][15] != ele[22][16];
    ele[20][15] != ele[22][17];
    ele[20][15] != ele[22][18];
    ele[20][15] != ele[22][19];
    ele[20][15] != ele[23][15];
    ele[20][15] != ele[23][16];
    ele[20][15] != ele[23][17];
    ele[20][15] != ele[23][18];
    ele[20][15] != ele[23][19];
    ele[20][15] != ele[24][15];
    ele[20][15] != ele[24][16];
    ele[20][15] != ele[24][17];
    ele[20][15] != ele[24][18];
    ele[20][15] != ele[24][19];
    ele[20][16] != ele[20][17];
    ele[20][16] != ele[20][18];
    ele[20][16] != ele[20][19];
    ele[20][16] != ele[20][20];
    ele[20][16] != ele[20][21];
    ele[20][16] != ele[20][22];
    ele[20][16] != ele[20][23];
    ele[20][16] != ele[20][24];
    ele[20][16] != ele[21][15];
    ele[20][16] != ele[21][16];
    ele[20][16] != ele[21][17];
    ele[20][16] != ele[21][18];
    ele[20][16] != ele[21][19];
    ele[20][16] != ele[22][15];
    ele[20][16] != ele[22][16];
    ele[20][16] != ele[22][17];
    ele[20][16] != ele[22][18];
    ele[20][16] != ele[22][19];
    ele[20][16] != ele[23][15];
    ele[20][16] != ele[23][16];
    ele[20][16] != ele[23][17];
    ele[20][16] != ele[23][18];
    ele[20][16] != ele[23][19];
    ele[20][16] != ele[24][15];
    ele[20][16] != ele[24][16];
    ele[20][16] != ele[24][17];
    ele[20][16] != ele[24][18];
    ele[20][16] != ele[24][19];
    ele[20][17] != ele[20][18];
    ele[20][17] != ele[20][19];
    ele[20][17] != ele[20][20];
    ele[20][17] != ele[20][21];
    ele[20][17] != ele[20][22];
    ele[20][17] != ele[20][23];
    ele[20][17] != ele[20][24];
    ele[20][17] != ele[21][15];
    ele[20][17] != ele[21][16];
    ele[20][17] != ele[21][17];
    ele[20][17] != ele[21][18];
    ele[20][17] != ele[21][19];
    ele[20][17] != ele[22][15];
    ele[20][17] != ele[22][16];
    ele[20][17] != ele[22][17];
    ele[20][17] != ele[22][18];
    ele[20][17] != ele[22][19];
    ele[20][17] != ele[23][15];
    ele[20][17] != ele[23][16];
    ele[20][17] != ele[23][17];
    ele[20][17] != ele[23][18];
    ele[20][17] != ele[23][19];
    ele[20][17] != ele[24][15];
    ele[20][17] != ele[24][16];
    ele[20][17] != ele[24][17];
    ele[20][17] != ele[24][18];
    ele[20][17] != ele[24][19];
    ele[20][18] != ele[20][19];
    ele[20][18] != ele[20][20];
    ele[20][18] != ele[20][21];
    ele[20][18] != ele[20][22];
    ele[20][18] != ele[20][23];
    ele[20][18] != ele[20][24];
    ele[20][18] != ele[21][15];
    ele[20][18] != ele[21][16];
    ele[20][18] != ele[21][17];
    ele[20][18] != ele[21][18];
    ele[20][18] != ele[21][19];
    ele[20][18] != ele[22][15];
    ele[20][18] != ele[22][16];
    ele[20][18] != ele[22][17];
    ele[20][18] != ele[22][18];
    ele[20][18] != ele[22][19];
    ele[20][18] != ele[23][15];
    ele[20][18] != ele[23][16];
    ele[20][18] != ele[23][17];
    ele[20][18] != ele[23][18];
    ele[20][18] != ele[23][19];
    ele[20][18] != ele[24][15];
    ele[20][18] != ele[24][16];
    ele[20][18] != ele[24][17];
    ele[20][18] != ele[24][18];
    ele[20][18] != ele[24][19];
    ele[20][19] != ele[20][20];
    ele[20][19] != ele[20][21];
    ele[20][19] != ele[20][22];
    ele[20][19] != ele[20][23];
    ele[20][19] != ele[20][24];
    ele[20][19] != ele[21][15];
    ele[20][19] != ele[21][16];
    ele[20][19] != ele[21][17];
    ele[20][19] != ele[21][18];
    ele[20][19] != ele[21][19];
    ele[20][19] != ele[22][15];
    ele[20][19] != ele[22][16];
    ele[20][19] != ele[22][17];
    ele[20][19] != ele[22][18];
    ele[20][19] != ele[22][19];
    ele[20][19] != ele[23][15];
    ele[20][19] != ele[23][16];
    ele[20][19] != ele[23][17];
    ele[20][19] != ele[23][18];
    ele[20][19] != ele[23][19];
    ele[20][19] != ele[24][15];
    ele[20][19] != ele[24][16];
    ele[20][19] != ele[24][17];
    ele[20][19] != ele[24][18];
    ele[20][19] != ele[24][19];
    ele[20][2] != ele[20][10];
    ele[20][2] != ele[20][11];
    ele[20][2] != ele[20][12];
    ele[20][2] != ele[20][13];
    ele[20][2] != ele[20][14];
    ele[20][2] != ele[20][15];
    ele[20][2] != ele[20][16];
    ele[20][2] != ele[20][17];
    ele[20][2] != ele[20][18];
    ele[20][2] != ele[20][19];
    ele[20][2] != ele[20][20];
    ele[20][2] != ele[20][21];
    ele[20][2] != ele[20][22];
    ele[20][2] != ele[20][23];
    ele[20][2] != ele[20][24];
    ele[20][2] != ele[20][3];
    ele[20][2] != ele[20][4];
    ele[20][2] != ele[20][5];
    ele[20][2] != ele[20][6];
    ele[20][2] != ele[20][7];
    ele[20][2] != ele[20][8];
    ele[20][2] != ele[20][9];
    ele[20][2] != ele[21][0];
    ele[20][2] != ele[21][1];
    ele[20][2] != ele[21][2];
    ele[20][2] != ele[21][3];
    ele[20][2] != ele[21][4];
    ele[20][2] != ele[22][0];
    ele[20][2] != ele[22][1];
    ele[20][2] != ele[22][2];
    ele[20][2] != ele[22][3];
    ele[20][2] != ele[22][4];
    ele[20][2] != ele[23][0];
    ele[20][2] != ele[23][1];
    ele[20][2] != ele[23][2];
    ele[20][2] != ele[23][3];
    ele[20][2] != ele[23][4];
    ele[20][2] != ele[24][0];
    ele[20][2] != ele[24][1];
    ele[20][2] != ele[24][2];
    ele[20][2] != ele[24][3];
    ele[20][2] != ele[24][4];
    ele[20][20] != ele[20][21];
    ele[20][20] != ele[20][22];
    ele[20][20] != ele[20][23];
    ele[20][20] != ele[20][24];
    ele[20][20] != ele[21][20];
    ele[20][20] != ele[21][21];
    ele[20][20] != ele[21][22];
    ele[20][20] != ele[21][23];
    ele[20][20] != ele[21][24];
    ele[20][20] != ele[22][20];
    ele[20][20] != ele[22][21];
    ele[20][20] != ele[22][22];
    ele[20][20] != ele[22][23];
    ele[20][20] != ele[22][24];
    ele[20][20] != ele[23][20];
    ele[20][20] != ele[23][21];
    ele[20][20] != ele[23][22];
    ele[20][20] != ele[23][23];
    ele[20][20] != ele[23][24];
    ele[20][20] != ele[24][20];
    ele[20][20] != ele[24][21];
    ele[20][20] != ele[24][22];
    ele[20][20] != ele[24][23];
    ele[20][20] != ele[24][24];
    ele[20][21] != ele[20][22];
    ele[20][21] != ele[20][23];
    ele[20][21] != ele[20][24];
    ele[20][21] != ele[21][20];
    ele[20][21] != ele[21][21];
    ele[20][21] != ele[21][22];
    ele[20][21] != ele[21][23];
    ele[20][21] != ele[21][24];
    ele[20][21] != ele[22][20];
    ele[20][21] != ele[22][21];
    ele[20][21] != ele[22][22];
    ele[20][21] != ele[22][23];
    ele[20][21] != ele[22][24];
    ele[20][21] != ele[23][20];
    ele[20][21] != ele[23][21];
    ele[20][21] != ele[23][22];
    ele[20][21] != ele[23][23];
    ele[20][21] != ele[23][24];
    ele[20][21] != ele[24][20];
    ele[20][21] != ele[24][21];
    ele[20][21] != ele[24][22];
    ele[20][21] != ele[24][23];
    ele[20][21] != ele[24][24];
    ele[20][22] != ele[20][23];
    ele[20][22] != ele[20][24];
    ele[20][22] != ele[21][20];
    ele[20][22] != ele[21][21];
    ele[20][22] != ele[21][22];
    ele[20][22] != ele[21][23];
    ele[20][22] != ele[21][24];
    ele[20][22] != ele[22][20];
    ele[20][22] != ele[22][21];
    ele[20][22] != ele[22][22];
    ele[20][22] != ele[22][23];
    ele[20][22] != ele[22][24];
    ele[20][22] != ele[23][20];
    ele[20][22] != ele[23][21];
    ele[20][22] != ele[23][22];
    ele[20][22] != ele[23][23];
    ele[20][22] != ele[23][24];
    ele[20][22] != ele[24][20];
    ele[20][22] != ele[24][21];
    ele[20][22] != ele[24][22];
    ele[20][22] != ele[24][23];
    ele[20][22] != ele[24][24];
    ele[20][23] != ele[20][24];
    ele[20][23] != ele[21][20];
    ele[20][23] != ele[21][21];
    ele[20][23] != ele[21][22];
    ele[20][23] != ele[21][23];
    ele[20][23] != ele[21][24];
    ele[20][23] != ele[22][20];
    ele[20][23] != ele[22][21];
    ele[20][23] != ele[22][22];
    ele[20][23] != ele[22][23];
    ele[20][23] != ele[22][24];
    ele[20][23] != ele[23][20];
    ele[20][23] != ele[23][21];
    ele[20][23] != ele[23][22];
    ele[20][23] != ele[23][23];
    ele[20][23] != ele[23][24];
    ele[20][23] != ele[24][20];
    ele[20][23] != ele[24][21];
    ele[20][23] != ele[24][22];
    ele[20][23] != ele[24][23];
    ele[20][23] != ele[24][24];
    ele[20][24] != ele[21][20];
    ele[20][24] != ele[21][21];
    ele[20][24] != ele[21][22];
    ele[20][24] != ele[21][23];
    ele[20][24] != ele[21][24];
    ele[20][24] != ele[22][20];
    ele[20][24] != ele[22][21];
    ele[20][24] != ele[22][22];
    ele[20][24] != ele[22][23];
    ele[20][24] != ele[22][24];
    ele[20][24] != ele[23][20];
    ele[20][24] != ele[23][21];
    ele[20][24] != ele[23][22];
    ele[20][24] != ele[23][23];
    ele[20][24] != ele[23][24];
    ele[20][24] != ele[24][20];
    ele[20][24] != ele[24][21];
    ele[20][24] != ele[24][22];
    ele[20][24] != ele[24][23];
    ele[20][24] != ele[24][24];
    ele[20][3] != ele[20][10];
    ele[20][3] != ele[20][11];
    ele[20][3] != ele[20][12];
    ele[20][3] != ele[20][13];
    ele[20][3] != ele[20][14];
    ele[20][3] != ele[20][15];
    ele[20][3] != ele[20][16];
    ele[20][3] != ele[20][17];
    ele[20][3] != ele[20][18];
    ele[20][3] != ele[20][19];
    ele[20][3] != ele[20][20];
    ele[20][3] != ele[20][21];
    ele[20][3] != ele[20][22];
    ele[20][3] != ele[20][23];
    ele[20][3] != ele[20][24];
    ele[20][3] != ele[20][4];
    ele[20][3] != ele[20][5];
    ele[20][3] != ele[20][6];
    ele[20][3] != ele[20][7];
    ele[20][3] != ele[20][8];
    ele[20][3] != ele[20][9];
    ele[20][3] != ele[21][0];
    ele[20][3] != ele[21][1];
    ele[20][3] != ele[21][2];
    ele[20][3] != ele[21][3];
    ele[20][3] != ele[21][4];
    ele[20][3] != ele[22][0];
    ele[20][3] != ele[22][1];
    ele[20][3] != ele[22][2];
    ele[20][3] != ele[22][3];
    ele[20][3] != ele[22][4];
    ele[20][3] != ele[23][0];
    ele[20][3] != ele[23][1];
    ele[20][3] != ele[23][2];
    ele[20][3] != ele[23][3];
    ele[20][3] != ele[23][4];
    ele[20][3] != ele[24][0];
    ele[20][3] != ele[24][1];
    ele[20][3] != ele[24][2];
    ele[20][3] != ele[24][3];
    ele[20][3] != ele[24][4];
    ele[20][4] != ele[20][10];
    ele[20][4] != ele[20][11];
    ele[20][4] != ele[20][12];
    ele[20][4] != ele[20][13];
    ele[20][4] != ele[20][14];
    ele[20][4] != ele[20][15];
    ele[20][4] != ele[20][16];
    ele[20][4] != ele[20][17];
    ele[20][4] != ele[20][18];
    ele[20][4] != ele[20][19];
    ele[20][4] != ele[20][20];
    ele[20][4] != ele[20][21];
    ele[20][4] != ele[20][22];
    ele[20][4] != ele[20][23];
    ele[20][4] != ele[20][24];
    ele[20][4] != ele[20][5];
    ele[20][4] != ele[20][6];
    ele[20][4] != ele[20][7];
    ele[20][4] != ele[20][8];
    ele[20][4] != ele[20][9];
    ele[20][4] != ele[21][0];
    ele[20][4] != ele[21][1];
    ele[20][4] != ele[21][2];
    ele[20][4] != ele[21][3];
    ele[20][4] != ele[21][4];
    ele[20][4] != ele[22][0];
    ele[20][4] != ele[22][1];
    ele[20][4] != ele[22][2];
    ele[20][4] != ele[22][3];
    ele[20][4] != ele[22][4];
    ele[20][4] != ele[23][0];
    ele[20][4] != ele[23][1];
    ele[20][4] != ele[23][2];
    ele[20][4] != ele[23][3];
    ele[20][4] != ele[23][4];
    ele[20][4] != ele[24][0];
    ele[20][4] != ele[24][1];
    ele[20][4] != ele[24][2];
    ele[20][4] != ele[24][3];
    ele[20][4] != ele[24][4];
    ele[20][5] != ele[20][10];
    ele[20][5] != ele[20][11];
    ele[20][5] != ele[20][12];
    ele[20][5] != ele[20][13];
    ele[20][5] != ele[20][14];
    ele[20][5] != ele[20][15];
    ele[20][5] != ele[20][16];
    ele[20][5] != ele[20][17];
    ele[20][5] != ele[20][18];
    ele[20][5] != ele[20][19];
    ele[20][5] != ele[20][20];
    ele[20][5] != ele[20][21];
    ele[20][5] != ele[20][22];
    ele[20][5] != ele[20][23];
    ele[20][5] != ele[20][24];
    ele[20][5] != ele[20][6];
    ele[20][5] != ele[20][7];
    ele[20][5] != ele[20][8];
    ele[20][5] != ele[20][9];
    ele[20][5] != ele[21][5];
    ele[20][5] != ele[21][6];
    ele[20][5] != ele[21][7];
    ele[20][5] != ele[21][8];
    ele[20][5] != ele[21][9];
    ele[20][5] != ele[22][5];
    ele[20][5] != ele[22][6];
    ele[20][5] != ele[22][7];
    ele[20][5] != ele[22][8];
    ele[20][5] != ele[22][9];
    ele[20][5] != ele[23][5];
    ele[20][5] != ele[23][6];
    ele[20][5] != ele[23][7];
    ele[20][5] != ele[23][8];
    ele[20][5] != ele[23][9];
    ele[20][5] != ele[24][5];
    ele[20][5] != ele[24][6];
    ele[20][5] != ele[24][7];
    ele[20][5] != ele[24][8];
    ele[20][5] != ele[24][9];
    ele[20][6] != ele[20][10];
    ele[20][6] != ele[20][11];
    ele[20][6] != ele[20][12];
    ele[20][6] != ele[20][13];
    ele[20][6] != ele[20][14];
    ele[20][6] != ele[20][15];
    ele[20][6] != ele[20][16];
    ele[20][6] != ele[20][17];
    ele[20][6] != ele[20][18];
    ele[20][6] != ele[20][19];
    ele[20][6] != ele[20][20];
    ele[20][6] != ele[20][21];
    ele[20][6] != ele[20][22];
    ele[20][6] != ele[20][23];
    ele[20][6] != ele[20][24];
    ele[20][6] != ele[20][7];
    ele[20][6] != ele[20][8];
    ele[20][6] != ele[20][9];
    ele[20][6] != ele[21][5];
    ele[20][6] != ele[21][6];
    ele[20][6] != ele[21][7];
    ele[20][6] != ele[21][8];
    ele[20][6] != ele[21][9];
    ele[20][6] != ele[22][5];
    ele[20][6] != ele[22][6];
    ele[20][6] != ele[22][7];
    ele[20][6] != ele[22][8];
    ele[20][6] != ele[22][9];
    ele[20][6] != ele[23][5];
    ele[20][6] != ele[23][6];
    ele[20][6] != ele[23][7];
    ele[20][6] != ele[23][8];
    ele[20][6] != ele[23][9];
    ele[20][6] != ele[24][5];
    ele[20][6] != ele[24][6];
    ele[20][6] != ele[24][7];
    ele[20][6] != ele[24][8];
    ele[20][6] != ele[24][9];
    ele[20][7] != ele[20][10];
    ele[20][7] != ele[20][11];
    ele[20][7] != ele[20][12];
    ele[20][7] != ele[20][13];
    ele[20][7] != ele[20][14];
    ele[20][7] != ele[20][15];
    ele[20][7] != ele[20][16];
    ele[20][7] != ele[20][17];
    ele[20][7] != ele[20][18];
    ele[20][7] != ele[20][19];
    ele[20][7] != ele[20][20];
    ele[20][7] != ele[20][21];
    ele[20][7] != ele[20][22];
    ele[20][7] != ele[20][23];
    ele[20][7] != ele[20][24];
    ele[20][7] != ele[20][8];
    ele[20][7] != ele[20][9];
    ele[20][7] != ele[21][5];
    ele[20][7] != ele[21][6];
    ele[20][7] != ele[21][7];
    ele[20][7] != ele[21][8];
    ele[20][7] != ele[21][9];
    ele[20][7] != ele[22][5];
    ele[20][7] != ele[22][6];
    ele[20][7] != ele[22][7];
    ele[20][7] != ele[22][8];
    ele[20][7] != ele[22][9];
    ele[20][7] != ele[23][5];
    ele[20][7] != ele[23][6];
    ele[20][7] != ele[23][7];
    ele[20][7] != ele[23][8];
    ele[20][7] != ele[23][9];
    ele[20][7] != ele[24][5];
    ele[20][7] != ele[24][6];
    ele[20][7] != ele[24][7];
    ele[20][7] != ele[24][8];
    ele[20][7] != ele[24][9];
    ele[20][8] != ele[20][10];
    ele[20][8] != ele[20][11];
    ele[20][8] != ele[20][12];
    ele[20][8] != ele[20][13];
    ele[20][8] != ele[20][14];
    ele[20][8] != ele[20][15];
    ele[20][8] != ele[20][16];
    ele[20][8] != ele[20][17];
    ele[20][8] != ele[20][18];
    ele[20][8] != ele[20][19];
    ele[20][8] != ele[20][20];
    ele[20][8] != ele[20][21];
    ele[20][8] != ele[20][22];
    ele[20][8] != ele[20][23];
    ele[20][8] != ele[20][24];
    ele[20][8] != ele[20][9];
    ele[20][8] != ele[21][5];
    ele[20][8] != ele[21][6];
    ele[20][8] != ele[21][7];
    ele[20][8] != ele[21][8];
    ele[20][8] != ele[21][9];
    ele[20][8] != ele[22][5];
    ele[20][8] != ele[22][6];
    ele[20][8] != ele[22][7];
    ele[20][8] != ele[22][8];
    ele[20][8] != ele[22][9];
    ele[20][8] != ele[23][5];
    ele[20][8] != ele[23][6];
    ele[20][8] != ele[23][7];
    ele[20][8] != ele[23][8];
    ele[20][8] != ele[23][9];
    ele[20][8] != ele[24][5];
    ele[20][8] != ele[24][6];
    ele[20][8] != ele[24][7];
    ele[20][8] != ele[24][8];
    ele[20][8] != ele[24][9];
    ele[20][9] != ele[20][10];
    ele[20][9] != ele[20][11];
    ele[20][9] != ele[20][12];
    ele[20][9] != ele[20][13];
    ele[20][9] != ele[20][14];
    ele[20][9] != ele[20][15];
    ele[20][9] != ele[20][16];
    ele[20][9] != ele[20][17];
    ele[20][9] != ele[20][18];
    ele[20][9] != ele[20][19];
    ele[20][9] != ele[20][20];
    ele[20][9] != ele[20][21];
    ele[20][9] != ele[20][22];
    ele[20][9] != ele[20][23];
    ele[20][9] != ele[20][24];
    ele[20][9] != ele[21][5];
    ele[20][9] != ele[21][6];
    ele[20][9] != ele[21][7];
    ele[20][9] != ele[21][8];
    ele[20][9] != ele[21][9];
    ele[20][9] != ele[22][5];
    ele[20][9] != ele[22][6];
    ele[20][9] != ele[22][7];
    ele[20][9] != ele[22][8];
    ele[20][9] != ele[22][9];
    ele[20][9] != ele[23][5];
    ele[20][9] != ele[23][6];
    ele[20][9] != ele[23][7];
    ele[20][9] != ele[23][8];
    ele[20][9] != ele[23][9];
    ele[20][9] != ele[24][5];
    ele[20][9] != ele[24][6];
    ele[20][9] != ele[24][7];
    ele[20][9] != ele[24][8];
    ele[20][9] != ele[24][9];
    ele[21][0] != ele[21][1];
    ele[21][0] != ele[21][10];
    ele[21][0] != ele[21][11];
    ele[21][0] != ele[21][12];
    ele[21][0] != ele[21][13];
    ele[21][0] != ele[21][14];
    ele[21][0] != ele[21][15];
    ele[21][0] != ele[21][16];
    ele[21][0] != ele[21][17];
    ele[21][0] != ele[21][18];
    ele[21][0] != ele[21][19];
    ele[21][0] != ele[21][2];
    ele[21][0] != ele[21][20];
    ele[21][0] != ele[21][21];
    ele[21][0] != ele[21][22];
    ele[21][0] != ele[21][23];
    ele[21][0] != ele[21][24];
    ele[21][0] != ele[21][3];
    ele[21][0] != ele[21][4];
    ele[21][0] != ele[21][5];
    ele[21][0] != ele[21][6];
    ele[21][0] != ele[21][7];
    ele[21][0] != ele[21][8];
    ele[21][0] != ele[21][9];
    ele[21][0] != ele[22][0];
    ele[21][0] != ele[22][1];
    ele[21][0] != ele[22][2];
    ele[21][0] != ele[22][3];
    ele[21][0] != ele[22][4];
    ele[21][0] != ele[23][0];
    ele[21][0] != ele[23][1];
    ele[21][0] != ele[23][2];
    ele[21][0] != ele[23][3];
    ele[21][0] != ele[23][4];
    ele[21][0] != ele[24][0];
    ele[21][0] != ele[24][1];
    ele[21][0] != ele[24][2];
    ele[21][0] != ele[24][3];
    ele[21][0] != ele[24][4];
    ele[21][1] != ele[21][10];
    ele[21][1] != ele[21][11];
    ele[21][1] != ele[21][12];
    ele[21][1] != ele[21][13];
    ele[21][1] != ele[21][14];
    ele[21][1] != ele[21][15];
    ele[21][1] != ele[21][16];
    ele[21][1] != ele[21][17];
    ele[21][1] != ele[21][18];
    ele[21][1] != ele[21][19];
    ele[21][1] != ele[21][2];
    ele[21][1] != ele[21][20];
    ele[21][1] != ele[21][21];
    ele[21][1] != ele[21][22];
    ele[21][1] != ele[21][23];
    ele[21][1] != ele[21][24];
    ele[21][1] != ele[21][3];
    ele[21][1] != ele[21][4];
    ele[21][1] != ele[21][5];
    ele[21][1] != ele[21][6];
    ele[21][1] != ele[21][7];
    ele[21][1] != ele[21][8];
    ele[21][1] != ele[21][9];
    ele[21][1] != ele[22][0];
    ele[21][1] != ele[22][1];
    ele[21][1] != ele[22][2];
    ele[21][1] != ele[22][3];
    ele[21][1] != ele[22][4];
    ele[21][1] != ele[23][0];
    ele[21][1] != ele[23][1];
    ele[21][1] != ele[23][2];
    ele[21][1] != ele[23][3];
    ele[21][1] != ele[23][4];
    ele[21][1] != ele[24][0];
    ele[21][1] != ele[24][1];
    ele[21][1] != ele[24][2];
    ele[21][1] != ele[24][3];
    ele[21][1] != ele[24][4];
    ele[21][10] != ele[21][11];
    ele[21][10] != ele[21][12];
    ele[21][10] != ele[21][13];
    ele[21][10] != ele[21][14];
    ele[21][10] != ele[21][15];
    ele[21][10] != ele[21][16];
    ele[21][10] != ele[21][17];
    ele[21][10] != ele[21][18];
    ele[21][10] != ele[21][19];
    ele[21][10] != ele[21][20];
    ele[21][10] != ele[21][21];
    ele[21][10] != ele[21][22];
    ele[21][10] != ele[21][23];
    ele[21][10] != ele[21][24];
    ele[21][10] != ele[22][10];
    ele[21][10] != ele[22][11];
    ele[21][10] != ele[22][12];
    ele[21][10] != ele[22][13];
    ele[21][10] != ele[22][14];
    ele[21][10] != ele[23][10];
    ele[21][10] != ele[23][11];
    ele[21][10] != ele[23][12];
    ele[21][10] != ele[23][13];
    ele[21][10] != ele[23][14];
    ele[21][10] != ele[24][10];
    ele[21][10] != ele[24][11];
    ele[21][10] != ele[24][12];
    ele[21][10] != ele[24][13];
    ele[21][10] != ele[24][14];
    ele[21][11] != ele[21][12];
    ele[21][11] != ele[21][13];
    ele[21][11] != ele[21][14];
    ele[21][11] != ele[21][15];
    ele[21][11] != ele[21][16];
    ele[21][11] != ele[21][17];
    ele[21][11] != ele[21][18];
    ele[21][11] != ele[21][19];
    ele[21][11] != ele[21][20];
    ele[21][11] != ele[21][21];
    ele[21][11] != ele[21][22];
    ele[21][11] != ele[21][23];
    ele[21][11] != ele[21][24];
    ele[21][11] != ele[22][10];
    ele[21][11] != ele[22][11];
    ele[21][11] != ele[22][12];
    ele[21][11] != ele[22][13];
    ele[21][11] != ele[22][14];
    ele[21][11] != ele[23][10];
    ele[21][11] != ele[23][11];
    ele[21][11] != ele[23][12];
    ele[21][11] != ele[23][13];
    ele[21][11] != ele[23][14];
    ele[21][11] != ele[24][10];
    ele[21][11] != ele[24][11];
    ele[21][11] != ele[24][12];
    ele[21][11] != ele[24][13];
    ele[21][11] != ele[24][14];
    ele[21][12] != ele[21][13];
    ele[21][12] != ele[21][14];
    ele[21][12] != ele[21][15];
    ele[21][12] != ele[21][16];
    ele[21][12] != ele[21][17];
    ele[21][12] != ele[21][18];
    ele[21][12] != ele[21][19];
    ele[21][12] != ele[21][20];
    ele[21][12] != ele[21][21];
    ele[21][12] != ele[21][22];
    ele[21][12] != ele[21][23];
    ele[21][12] != ele[21][24];
    ele[21][12] != ele[22][10];
    ele[21][12] != ele[22][11];
    ele[21][12] != ele[22][12];
    ele[21][12] != ele[22][13];
    ele[21][12] != ele[22][14];
    ele[21][12] != ele[23][10];
    ele[21][12] != ele[23][11];
    ele[21][12] != ele[23][12];
    ele[21][12] != ele[23][13];
    ele[21][12] != ele[23][14];
    ele[21][12] != ele[24][10];
    ele[21][12] != ele[24][11];
    ele[21][12] != ele[24][12];
    ele[21][12] != ele[24][13];
    ele[21][12] != ele[24][14];
    ele[21][13] != ele[21][14];
    ele[21][13] != ele[21][15];
    ele[21][13] != ele[21][16];
    ele[21][13] != ele[21][17];
    ele[21][13] != ele[21][18];
    ele[21][13] != ele[21][19];
    ele[21][13] != ele[21][20];
    ele[21][13] != ele[21][21];
    ele[21][13] != ele[21][22];
    ele[21][13] != ele[21][23];
    ele[21][13] != ele[21][24];
    ele[21][13] != ele[22][10];
    ele[21][13] != ele[22][11];
    ele[21][13] != ele[22][12];
    ele[21][13] != ele[22][13];
    ele[21][13] != ele[22][14];
    ele[21][13] != ele[23][10];
    ele[21][13] != ele[23][11];
    ele[21][13] != ele[23][12];
    ele[21][13] != ele[23][13];
    ele[21][13] != ele[23][14];
    ele[21][13] != ele[24][10];
    ele[21][13] != ele[24][11];
    ele[21][13] != ele[24][12];
    ele[21][13] != ele[24][13];
    ele[21][13] != ele[24][14];
    ele[21][14] != ele[21][15];
    ele[21][14] != ele[21][16];
    ele[21][14] != ele[21][17];
    ele[21][14] != ele[21][18];
    ele[21][14] != ele[21][19];
    ele[21][14] != ele[21][20];
    ele[21][14] != ele[21][21];
    ele[21][14] != ele[21][22];
    ele[21][14] != ele[21][23];
    ele[21][14] != ele[21][24];
    ele[21][14] != ele[22][10];
    ele[21][14] != ele[22][11];
    ele[21][14] != ele[22][12];
    ele[21][14] != ele[22][13];
    ele[21][14] != ele[22][14];
    ele[21][14] != ele[23][10];
    ele[21][14] != ele[23][11];
    ele[21][14] != ele[23][12];
    ele[21][14] != ele[23][13];
    ele[21][14] != ele[23][14];
    ele[21][14] != ele[24][10];
    ele[21][14] != ele[24][11];
    ele[21][14] != ele[24][12];
    ele[21][14] != ele[24][13];
    ele[21][14] != ele[24][14];
    ele[21][15] != ele[21][16];
    ele[21][15] != ele[21][17];
    ele[21][15] != ele[21][18];
    ele[21][15] != ele[21][19];
    ele[21][15] != ele[21][20];
    ele[21][15] != ele[21][21];
    ele[21][15] != ele[21][22];
    ele[21][15] != ele[21][23];
    ele[21][15] != ele[21][24];
    ele[21][15] != ele[22][15];
    ele[21][15] != ele[22][16];
    ele[21][15] != ele[22][17];
    ele[21][15] != ele[22][18];
    ele[21][15] != ele[22][19];
    ele[21][15] != ele[23][15];
    ele[21][15] != ele[23][16];
    ele[21][15] != ele[23][17];
    ele[21][15] != ele[23][18];
    ele[21][15] != ele[23][19];
    ele[21][15] != ele[24][15];
    ele[21][15] != ele[24][16];
    ele[21][15] != ele[24][17];
    ele[21][15] != ele[24][18];
    ele[21][15] != ele[24][19];
    ele[21][16] != ele[21][17];
    ele[21][16] != ele[21][18];
    ele[21][16] != ele[21][19];
    ele[21][16] != ele[21][20];
    ele[21][16] != ele[21][21];
    ele[21][16] != ele[21][22];
    ele[21][16] != ele[21][23];
    ele[21][16] != ele[21][24];
    ele[21][16] != ele[22][15];
    ele[21][16] != ele[22][16];
    ele[21][16] != ele[22][17];
    ele[21][16] != ele[22][18];
    ele[21][16] != ele[22][19];
    ele[21][16] != ele[23][15];
    ele[21][16] != ele[23][16];
    ele[21][16] != ele[23][17];
    ele[21][16] != ele[23][18];
    ele[21][16] != ele[23][19];
    ele[21][16] != ele[24][15];
    ele[21][16] != ele[24][16];
    ele[21][16] != ele[24][17];
    ele[21][16] != ele[24][18];
    ele[21][16] != ele[24][19];
    ele[21][17] != ele[21][18];
    ele[21][17] != ele[21][19];
    ele[21][17] != ele[21][20];
    ele[21][17] != ele[21][21];
    ele[21][17] != ele[21][22];
    ele[21][17] != ele[21][23];
    ele[21][17] != ele[21][24];
    ele[21][17] != ele[22][15];
    ele[21][17] != ele[22][16];
    ele[21][17] != ele[22][17];
    ele[21][17] != ele[22][18];
    ele[21][17] != ele[22][19];
    ele[21][17] != ele[23][15];
    ele[21][17] != ele[23][16];
    ele[21][17] != ele[23][17];
    ele[21][17] != ele[23][18];
    ele[21][17] != ele[23][19];
    ele[21][17] != ele[24][15];
    ele[21][17] != ele[24][16];
    ele[21][17] != ele[24][17];
    ele[21][17] != ele[24][18];
    ele[21][17] != ele[24][19];
    ele[21][18] != ele[21][19];
    ele[21][18] != ele[21][20];
    ele[21][18] != ele[21][21];
    ele[21][18] != ele[21][22];
    ele[21][18] != ele[21][23];
    ele[21][18] != ele[21][24];
    ele[21][18] != ele[22][15];
    ele[21][18] != ele[22][16];
    ele[21][18] != ele[22][17];
    ele[21][18] != ele[22][18];
    ele[21][18] != ele[22][19];
    ele[21][18] != ele[23][15];
    ele[21][18] != ele[23][16];
    ele[21][18] != ele[23][17];
    ele[21][18] != ele[23][18];
    ele[21][18] != ele[23][19];
    ele[21][18] != ele[24][15];
    ele[21][18] != ele[24][16];
    ele[21][18] != ele[24][17];
    ele[21][18] != ele[24][18];
    ele[21][18] != ele[24][19];
    ele[21][19] != ele[21][20];
    ele[21][19] != ele[21][21];
    ele[21][19] != ele[21][22];
    ele[21][19] != ele[21][23];
    ele[21][19] != ele[21][24];
    ele[21][19] != ele[22][15];
    ele[21][19] != ele[22][16];
    ele[21][19] != ele[22][17];
    ele[21][19] != ele[22][18];
    ele[21][19] != ele[22][19];
    ele[21][19] != ele[23][15];
    ele[21][19] != ele[23][16];
    ele[21][19] != ele[23][17];
    ele[21][19] != ele[23][18];
    ele[21][19] != ele[23][19];
    ele[21][19] != ele[24][15];
    ele[21][19] != ele[24][16];
    ele[21][19] != ele[24][17];
    ele[21][19] != ele[24][18];
    ele[21][19] != ele[24][19];
    ele[21][2] != ele[21][10];
    ele[21][2] != ele[21][11];
    ele[21][2] != ele[21][12];
    ele[21][2] != ele[21][13];
    ele[21][2] != ele[21][14];
    ele[21][2] != ele[21][15];
    ele[21][2] != ele[21][16];
    ele[21][2] != ele[21][17];
    ele[21][2] != ele[21][18];
    ele[21][2] != ele[21][19];
    ele[21][2] != ele[21][20];
    ele[21][2] != ele[21][21];
    ele[21][2] != ele[21][22];
    ele[21][2] != ele[21][23];
    ele[21][2] != ele[21][24];
    ele[21][2] != ele[21][3];
    ele[21][2] != ele[21][4];
    ele[21][2] != ele[21][5];
    ele[21][2] != ele[21][6];
    ele[21][2] != ele[21][7];
    ele[21][2] != ele[21][8];
    ele[21][2] != ele[21][9];
    ele[21][2] != ele[22][0];
    ele[21][2] != ele[22][1];
    ele[21][2] != ele[22][2];
    ele[21][2] != ele[22][3];
    ele[21][2] != ele[22][4];
    ele[21][2] != ele[23][0];
    ele[21][2] != ele[23][1];
    ele[21][2] != ele[23][2];
    ele[21][2] != ele[23][3];
    ele[21][2] != ele[23][4];
    ele[21][2] != ele[24][0];
    ele[21][2] != ele[24][1];
    ele[21][2] != ele[24][2];
    ele[21][2] != ele[24][3];
    ele[21][2] != ele[24][4];
    ele[21][20] != ele[21][21];
    ele[21][20] != ele[21][22];
    ele[21][20] != ele[21][23];
    ele[21][20] != ele[21][24];
    ele[21][20] != ele[22][20];
    ele[21][20] != ele[22][21];
    ele[21][20] != ele[22][22];
    ele[21][20] != ele[22][23];
    ele[21][20] != ele[22][24];
    ele[21][20] != ele[23][20];
    ele[21][20] != ele[23][21];
    ele[21][20] != ele[23][22];
    ele[21][20] != ele[23][23];
    ele[21][20] != ele[23][24];
    ele[21][20] != ele[24][20];
    ele[21][20] != ele[24][21];
    ele[21][20] != ele[24][22];
    ele[21][20] != ele[24][23];
    ele[21][20] != ele[24][24];
    ele[21][21] != ele[21][22];
    ele[21][21] != ele[21][23];
    ele[21][21] != ele[21][24];
    ele[21][21] != ele[22][20];
    ele[21][21] != ele[22][21];
    ele[21][21] != ele[22][22];
    ele[21][21] != ele[22][23];
    ele[21][21] != ele[22][24];
    ele[21][21] != ele[23][20];
    ele[21][21] != ele[23][21];
    ele[21][21] != ele[23][22];
    ele[21][21] != ele[23][23];
    ele[21][21] != ele[23][24];
    ele[21][21] != ele[24][20];
    ele[21][21] != ele[24][21];
    ele[21][21] != ele[24][22];
    ele[21][21] != ele[24][23];
    ele[21][21] != ele[24][24];
    ele[21][22] != ele[21][23];
    ele[21][22] != ele[21][24];
    ele[21][22] != ele[22][20];
    ele[21][22] != ele[22][21];
    ele[21][22] != ele[22][22];
    ele[21][22] != ele[22][23];
    ele[21][22] != ele[22][24];
    ele[21][22] != ele[23][20];
    ele[21][22] != ele[23][21];
    ele[21][22] != ele[23][22];
    ele[21][22] != ele[23][23];
    ele[21][22] != ele[23][24];
    ele[21][22] != ele[24][20];
    ele[21][22] != ele[24][21];
    ele[21][22] != ele[24][22];
    ele[21][22] != ele[24][23];
    ele[21][22] != ele[24][24];
    ele[21][23] != ele[21][24];
    ele[21][23] != ele[22][20];
    ele[21][23] != ele[22][21];
    ele[21][23] != ele[22][22];
    ele[21][23] != ele[22][23];
    ele[21][23] != ele[22][24];
    ele[21][23] != ele[23][20];
    ele[21][23] != ele[23][21];
    ele[21][23] != ele[23][22];
    ele[21][23] != ele[23][23];
    ele[21][23] != ele[23][24];
    ele[21][23] != ele[24][20];
    ele[21][23] != ele[24][21];
    ele[21][23] != ele[24][22];
    ele[21][23] != ele[24][23];
    ele[21][23] != ele[24][24];
    ele[21][24] != ele[22][20];
    ele[21][24] != ele[22][21];
    ele[21][24] != ele[22][22];
    ele[21][24] != ele[22][23];
    ele[21][24] != ele[22][24];
    ele[21][24] != ele[23][20];
    ele[21][24] != ele[23][21];
    ele[21][24] != ele[23][22];
    ele[21][24] != ele[23][23];
    ele[21][24] != ele[23][24];
    ele[21][24] != ele[24][20];
    ele[21][24] != ele[24][21];
    ele[21][24] != ele[24][22];
    ele[21][24] != ele[24][23];
    ele[21][24] != ele[24][24];
    ele[21][3] != ele[21][10];
    ele[21][3] != ele[21][11];
    ele[21][3] != ele[21][12];
    ele[21][3] != ele[21][13];
    ele[21][3] != ele[21][14];
    ele[21][3] != ele[21][15];
    ele[21][3] != ele[21][16];
    ele[21][3] != ele[21][17];
    ele[21][3] != ele[21][18];
    ele[21][3] != ele[21][19];
    ele[21][3] != ele[21][20];
    ele[21][3] != ele[21][21];
    ele[21][3] != ele[21][22];
    ele[21][3] != ele[21][23];
    ele[21][3] != ele[21][24];
    ele[21][3] != ele[21][4];
    ele[21][3] != ele[21][5];
    ele[21][3] != ele[21][6];
    ele[21][3] != ele[21][7];
    ele[21][3] != ele[21][8];
    ele[21][3] != ele[21][9];
    ele[21][3] != ele[22][0];
    ele[21][3] != ele[22][1];
    ele[21][3] != ele[22][2];
    ele[21][3] != ele[22][3];
    ele[21][3] != ele[22][4];
    ele[21][3] != ele[23][0];
    ele[21][3] != ele[23][1];
    ele[21][3] != ele[23][2];
    ele[21][3] != ele[23][3];
    ele[21][3] != ele[23][4];
    ele[21][3] != ele[24][0];
    ele[21][3] != ele[24][1];
    ele[21][3] != ele[24][2];
    ele[21][3] != ele[24][3];
    ele[21][3] != ele[24][4];
    ele[21][4] != ele[21][10];
    ele[21][4] != ele[21][11];
    ele[21][4] != ele[21][12];
    ele[21][4] != ele[21][13];
    ele[21][4] != ele[21][14];
    ele[21][4] != ele[21][15];
    ele[21][4] != ele[21][16];
    ele[21][4] != ele[21][17];
    ele[21][4] != ele[21][18];
    ele[21][4] != ele[21][19];
    ele[21][4] != ele[21][20];
    ele[21][4] != ele[21][21];
    ele[21][4] != ele[21][22];
    ele[21][4] != ele[21][23];
    ele[21][4] != ele[21][24];
    ele[21][4] != ele[21][5];
    ele[21][4] != ele[21][6];
    ele[21][4] != ele[21][7];
    ele[21][4] != ele[21][8];
    ele[21][4] != ele[21][9];
    ele[21][4] != ele[22][0];
    ele[21][4] != ele[22][1];
    ele[21][4] != ele[22][2];
    ele[21][4] != ele[22][3];
    ele[21][4] != ele[22][4];
    ele[21][4] != ele[23][0];
    ele[21][4] != ele[23][1];
    ele[21][4] != ele[23][2];
    ele[21][4] != ele[23][3];
    ele[21][4] != ele[23][4];
    ele[21][4] != ele[24][0];
    ele[21][4] != ele[24][1];
    ele[21][4] != ele[24][2];
    ele[21][4] != ele[24][3];
    ele[21][4] != ele[24][4];
    ele[21][5] != ele[21][10];
    ele[21][5] != ele[21][11];
    ele[21][5] != ele[21][12];
    ele[21][5] != ele[21][13];
    ele[21][5] != ele[21][14];
    ele[21][5] != ele[21][15];
    ele[21][5] != ele[21][16];
    ele[21][5] != ele[21][17];
    ele[21][5] != ele[21][18];
    ele[21][5] != ele[21][19];
    ele[21][5] != ele[21][20];
    ele[21][5] != ele[21][21];
    ele[21][5] != ele[21][22];
    ele[21][5] != ele[21][23];
    ele[21][5] != ele[21][24];
    ele[21][5] != ele[21][6];
    ele[21][5] != ele[21][7];
    ele[21][5] != ele[21][8];
    ele[21][5] != ele[21][9];
    ele[21][5] != ele[22][5];
    ele[21][5] != ele[22][6];
    ele[21][5] != ele[22][7];
    ele[21][5] != ele[22][8];
    ele[21][5] != ele[22][9];
    ele[21][5] != ele[23][5];
    ele[21][5] != ele[23][6];
    ele[21][5] != ele[23][7];
    ele[21][5] != ele[23][8];
    ele[21][5] != ele[23][9];
    ele[21][5] != ele[24][5];
    ele[21][5] != ele[24][6];
    ele[21][5] != ele[24][7];
    ele[21][5] != ele[24][8];
    ele[21][5] != ele[24][9];
    ele[21][6] != ele[21][10];
    ele[21][6] != ele[21][11];
    ele[21][6] != ele[21][12];
    ele[21][6] != ele[21][13];
    ele[21][6] != ele[21][14];
    ele[21][6] != ele[21][15];
    ele[21][6] != ele[21][16];
    ele[21][6] != ele[21][17];
    ele[21][6] != ele[21][18];
    ele[21][6] != ele[21][19];
    ele[21][6] != ele[21][20];
    ele[21][6] != ele[21][21];
    ele[21][6] != ele[21][22];
    ele[21][6] != ele[21][23];
    ele[21][6] != ele[21][24];
    ele[21][6] != ele[21][7];
    ele[21][6] != ele[21][8];
    ele[21][6] != ele[21][9];
    ele[21][6] != ele[22][5];
    ele[21][6] != ele[22][6];
    ele[21][6] != ele[22][7];
    ele[21][6] != ele[22][8];
    ele[21][6] != ele[22][9];
    ele[21][6] != ele[23][5];
    ele[21][6] != ele[23][6];
    ele[21][6] != ele[23][7];
    ele[21][6] != ele[23][8];
    ele[21][6] != ele[23][9];
    ele[21][6] != ele[24][5];
    ele[21][6] != ele[24][6];
    ele[21][6] != ele[24][7];
    ele[21][6] != ele[24][8];
    ele[21][6] != ele[24][9];
    ele[21][7] != ele[21][10];
    ele[21][7] != ele[21][11];
    ele[21][7] != ele[21][12];
    ele[21][7] != ele[21][13];
    ele[21][7] != ele[21][14];
    ele[21][7] != ele[21][15];
    ele[21][7] != ele[21][16];
    ele[21][7] != ele[21][17];
    ele[21][7] != ele[21][18];
    ele[21][7] != ele[21][19];
    ele[21][7] != ele[21][20];
    ele[21][7] != ele[21][21];
    ele[21][7] != ele[21][22];
    ele[21][7] != ele[21][23];
    ele[21][7] != ele[21][24];
    ele[21][7] != ele[21][8];
    ele[21][7] != ele[21][9];
    ele[21][7] != ele[22][5];
    ele[21][7] != ele[22][6];
    ele[21][7] != ele[22][7];
    ele[21][7] != ele[22][8];
    ele[21][7] != ele[22][9];
    ele[21][7] != ele[23][5];
    ele[21][7] != ele[23][6];
    ele[21][7] != ele[23][7];
    ele[21][7] != ele[23][8];
    ele[21][7] != ele[23][9];
    ele[21][7] != ele[24][5];
    ele[21][7] != ele[24][6];
    ele[21][7] != ele[24][7];
    ele[21][7] != ele[24][8];
    ele[21][7] != ele[24][9];
    ele[21][8] != ele[21][10];
    ele[21][8] != ele[21][11];
    ele[21][8] != ele[21][12];
    ele[21][8] != ele[21][13];
    ele[21][8] != ele[21][14];
    ele[21][8] != ele[21][15];
    ele[21][8] != ele[21][16];
    ele[21][8] != ele[21][17];
    ele[21][8] != ele[21][18];
    ele[21][8] != ele[21][19];
    ele[21][8] != ele[21][20];
    ele[21][8] != ele[21][21];
    ele[21][8] != ele[21][22];
    ele[21][8] != ele[21][23];
    ele[21][8] != ele[21][24];
    ele[21][8] != ele[21][9];
    ele[21][8] != ele[22][5];
    ele[21][8] != ele[22][6];
    ele[21][8] != ele[22][7];
    ele[21][8] != ele[22][8];
    ele[21][8] != ele[22][9];
    ele[21][8] != ele[23][5];
    ele[21][8] != ele[23][6];
    ele[21][8] != ele[23][7];
    ele[21][8] != ele[23][8];
    ele[21][8] != ele[23][9];
    ele[21][8] != ele[24][5];
    ele[21][8] != ele[24][6];
    ele[21][8] != ele[24][7];
    ele[21][8] != ele[24][8];
    ele[21][8] != ele[24][9];
    ele[21][9] != ele[21][10];
    ele[21][9] != ele[21][11];
    ele[21][9] != ele[21][12];
    ele[21][9] != ele[21][13];
    ele[21][9] != ele[21][14];
    ele[21][9] != ele[21][15];
    ele[21][9] != ele[21][16];
    ele[21][9] != ele[21][17];
    ele[21][9] != ele[21][18];
    ele[21][9] != ele[21][19];
    ele[21][9] != ele[21][20];
    ele[21][9] != ele[21][21];
    ele[21][9] != ele[21][22];
    ele[21][9] != ele[21][23];
    ele[21][9] != ele[21][24];
    ele[21][9] != ele[22][5];
    ele[21][9] != ele[22][6];
    ele[21][9] != ele[22][7];
    ele[21][9] != ele[22][8];
    ele[21][9] != ele[22][9];
    ele[21][9] != ele[23][5];
    ele[21][9] != ele[23][6];
    ele[21][9] != ele[23][7];
    ele[21][9] != ele[23][8];
    ele[21][9] != ele[23][9];
    ele[21][9] != ele[24][5];
    ele[21][9] != ele[24][6];
    ele[21][9] != ele[24][7];
    ele[21][9] != ele[24][8];
    ele[21][9] != ele[24][9];
    ele[22][0] != ele[22][1];
    ele[22][0] != ele[22][10];
    ele[22][0] != ele[22][11];
    ele[22][0] != ele[22][12];
    ele[22][0] != ele[22][13];
    ele[22][0] != ele[22][14];
    ele[22][0] != ele[22][15];
    ele[22][0] != ele[22][16];
    ele[22][0] != ele[22][17];
    ele[22][0] != ele[22][18];
    ele[22][0] != ele[22][19];
    ele[22][0] != ele[22][2];
    ele[22][0] != ele[22][20];
    ele[22][0] != ele[22][21];
    ele[22][0] != ele[22][22];
    ele[22][0] != ele[22][23];
    ele[22][0] != ele[22][24];
    ele[22][0] != ele[22][3];
    ele[22][0] != ele[22][4];
    ele[22][0] != ele[22][5];
    ele[22][0] != ele[22][6];
    ele[22][0] != ele[22][7];
    ele[22][0] != ele[22][8];
    ele[22][0] != ele[22][9];
    ele[22][0] != ele[23][0];
    ele[22][0] != ele[23][1];
    ele[22][0] != ele[23][2];
    ele[22][0] != ele[23][3];
    ele[22][0] != ele[23][4];
    ele[22][0] != ele[24][0];
    ele[22][0] != ele[24][1];
    ele[22][0] != ele[24][2];
    ele[22][0] != ele[24][3];
    ele[22][0] != ele[24][4];
    ele[22][1] != ele[22][10];
    ele[22][1] != ele[22][11];
    ele[22][1] != ele[22][12];
    ele[22][1] != ele[22][13];
    ele[22][1] != ele[22][14];
    ele[22][1] != ele[22][15];
    ele[22][1] != ele[22][16];
    ele[22][1] != ele[22][17];
    ele[22][1] != ele[22][18];
    ele[22][1] != ele[22][19];
    ele[22][1] != ele[22][2];
    ele[22][1] != ele[22][20];
    ele[22][1] != ele[22][21];
    ele[22][1] != ele[22][22];
    ele[22][1] != ele[22][23];
    ele[22][1] != ele[22][24];
    ele[22][1] != ele[22][3];
    ele[22][1] != ele[22][4];
    ele[22][1] != ele[22][5];
    ele[22][1] != ele[22][6];
    ele[22][1] != ele[22][7];
    ele[22][1] != ele[22][8];
    ele[22][1] != ele[22][9];
    ele[22][1] != ele[23][0];
    ele[22][1] != ele[23][1];
    ele[22][1] != ele[23][2];
    ele[22][1] != ele[23][3];
    ele[22][1] != ele[23][4];
    ele[22][1] != ele[24][0];
    ele[22][1] != ele[24][1];
    ele[22][1] != ele[24][2];
    ele[22][1] != ele[24][3];
    ele[22][1] != ele[24][4];
    ele[22][10] != ele[22][11];
    ele[22][10] != ele[22][12];
    ele[22][10] != ele[22][13];
    ele[22][10] != ele[22][14];
    ele[22][10] != ele[22][15];
    ele[22][10] != ele[22][16];
    ele[22][10] != ele[22][17];
    ele[22][10] != ele[22][18];
    ele[22][10] != ele[22][19];
    ele[22][10] != ele[22][20];
    ele[22][10] != ele[22][21];
    ele[22][10] != ele[22][22];
    ele[22][10] != ele[22][23];
    ele[22][10] != ele[22][24];
    ele[22][10] != ele[23][10];
    ele[22][10] != ele[23][11];
    ele[22][10] != ele[23][12];
    ele[22][10] != ele[23][13];
    ele[22][10] != ele[23][14];
    ele[22][10] != ele[24][10];
    ele[22][10] != ele[24][11];
    ele[22][10] != ele[24][12];
    ele[22][10] != ele[24][13];
    ele[22][10] != ele[24][14];
    ele[22][11] != ele[22][12];
    ele[22][11] != ele[22][13];
    ele[22][11] != ele[22][14];
    ele[22][11] != ele[22][15];
    ele[22][11] != ele[22][16];
    ele[22][11] != ele[22][17];
    ele[22][11] != ele[22][18];
    ele[22][11] != ele[22][19];
    ele[22][11] != ele[22][20];
    ele[22][11] != ele[22][21];
    ele[22][11] != ele[22][22];
    ele[22][11] != ele[22][23];
    ele[22][11] != ele[22][24];
    ele[22][11] != ele[23][10];
    ele[22][11] != ele[23][11];
    ele[22][11] != ele[23][12];
    ele[22][11] != ele[23][13];
    ele[22][11] != ele[23][14];
    ele[22][11] != ele[24][10];
    ele[22][11] != ele[24][11];
    ele[22][11] != ele[24][12];
    ele[22][11] != ele[24][13];
    ele[22][11] != ele[24][14];
    ele[22][12] != ele[22][13];
    ele[22][12] != ele[22][14];
    ele[22][12] != ele[22][15];
    ele[22][12] != ele[22][16];
    ele[22][12] != ele[22][17];
    ele[22][12] != ele[22][18];
    ele[22][12] != ele[22][19];
    ele[22][12] != ele[22][20];
    ele[22][12] != ele[22][21];
    ele[22][12] != ele[22][22];
    ele[22][12] != ele[22][23];
    ele[22][12] != ele[22][24];
    ele[22][12] != ele[23][10];
    ele[22][12] != ele[23][11];
    ele[22][12] != ele[23][12];
    ele[22][12] != ele[23][13];
    ele[22][12] != ele[23][14];
    ele[22][12] != ele[24][10];
    ele[22][12] != ele[24][11];
    ele[22][12] != ele[24][12];
    ele[22][12] != ele[24][13];
    ele[22][12] != ele[24][14];
    ele[22][13] != ele[22][14];
    ele[22][13] != ele[22][15];
    ele[22][13] != ele[22][16];
    ele[22][13] != ele[22][17];
    ele[22][13] != ele[22][18];
    ele[22][13] != ele[22][19];
    ele[22][13] != ele[22][20];
    ele[22][13] != ele[22][21];
    ele[22][13] != ele[22][22];
    ele[22][13] != ele[22][23];
    ele[22][13] != ele[22][24];
    ele[22][13] != ele[23][10];
    ele[22][13] != ele[23][11];
    ele[22][13] != ele[23][12];
    ele[22][13] != ele[23][13];
    ele[22][13] != ele[23][14];
    ele[22][13] != ele[24][10];
    ele[22][13] != ele[24][11];
    ele[22][13] != ele[24][12];
    ele[22][13] != ele[24][13];
    ele[22][13] != ele[24][14];
    ele[22][14] != ele[22][15];
    ele[22][14] != ele[22][16];
    ele[22][14] != ele[22][17];
    ele[22][14] != ele[22][18];
    ele[22][14] != ele[22][19];
    ele[22][14] != ele[22][20];
    ele[22][14] != ele[22][21];
    ele[22][14] != ele[22][22];
    ele[22][14] != ele[22][23];
    ele[22][14] != ele[22][24];
    ele[22][14] != ele[23][10];
    ele[22][14] != ele[23][11];
    ele[22][14] != ele[23][12];
    ele[22][14] != ele[23][13];
    ele[22][14] != ele[23][14];
    ele[22][14] != ele[24][10];
    ele[22][14] != ele[24][11];
    ele[22][14] != ele[24][12];
    ele[22][14] != ele[24][13];
    ele[22][14] != ele[24][14];
    ele[22][15] != ele[22][16];
    ele[22][15] != ele[22][17];
    ele[22][15] != ele[22][18];
    ele[22][15] != ele[22][19];
    ele[22][15] != ele[22][20];
    ele[22][15] != ele[22][21];
    ele[22][15] != ele[22][22];
    ele[22][15] != ele[22][23];
    ele[22][15] != ele[22][24];
    ele[22][15] != ele[23][15];
    ele[22][15] != ele[23][16];
    ele[22][15] != ele[23][17];
    ele[22][15] != ele[23][18];
    ele[22][15] != ele[23][19];
    ele[22][15] != ele[24][15];
    ele[22][15] != ele[24][16];
    ele[22][15] != ele[24][17];
    ele[22][15] != ele[24][18];
    ele[22][15] != ele[24][19];
    ele[22][16] != ele[22][17];
    ele[22][16] != ele[22][18];
    ele[22][16] != ele[22][19];
    ele[22][16] != ele[22][20];
    ele[22][16] != ele[22][21];
    ele[22][16] != ele[22][22];
    ele[22][16] != ele[22][23];
    ele[22][16] != ele[22][24];
    ele[22][16] != ele[23][15];
    ele[22][16] != ele[23][16];
    ele[22][16] != ele[23][17];
    ele[22][16] != ele[23][18];
    ele[22][16] != ele[23][19];
    ele[22][16] != ele[24][15];
    ele[22][16] != ele[24][16];
    ele[22][16] != ele[24][17];
    ele[22][16] != ele[24][18];
    ele[22][16] != ele[24][19];
    ele[22][17] != ele[22][18];
    ele[22][17] != ele[22][19];
    ele[22][17] != ele[22][20];
    ele[22][17] != ele[22][21];
    ele[22][17] != ele[22][22];
    ele[22][17] != ele[22][23];
    ele[22][17] != ele[22][24];
    ele[22][17] != ele[23][15];
    ele[22][17] != ele[23][16];
    ele[22][17] != ele[23][17];
    ele[22][17] != ele[23][18];
    ele[22][17] != ele[23][19];
    ele[22][17] != ele[24][15];
    ele[22][17] != ele[24][16];
    ele[22][17] != ele[24][17];
    ele[22][17] != ele[24][18];
    ele[22][17] != ele[24][19];
    ele[22][18] != ele[22][19];
    ele[22][18] != ele[22][20];
    ele[22][18] != ele[22][21];
    ele[22][18] != ele[22][22];
    ele[22][18] != ele[22][23];
    ele[22][18] != ele[22][24];
    ele[22][18] != ele[23][15];
    ele[22][18] != ele[23][16];
    ele[22][18] != ele[23][17];
    ele[22][18] != ele[23][18];
    ele[22][18] != ele[23][19];
    ele[22][18] != ele[24][15];
    ele[22][18] != ele[24][16];
    ele[22][18] != ele[24][17];
    ele[22][18] != ele[24][18];
    ele[22][18] != ele[24][19];
    ele[22][19] != ele[22][20];
    ele[22][19] != ele[22][21];
    ele[22][19] != ele[22][22];
    ele[22][19] != ele[22][23];
    ele[22][19] != ele[22][24];
    ele[22][19] != ele[23][15];
    ele[22][19] != ele[23][16];
    ele[22][19] != ele[23][17];
    ele[22][19] != ele[23][18];
    ele[22][19] != ele[23][19];
    ele[22][19] != ele[24][15];
    ele[22][19] != ele[24][16];
    ele[22][19] != ele[24][17];
    ele[22][19] != ele[24][18];
    ele[22][19] != ele[24][19];
    ele[22][2] != ele[22][10];
    ele[22][2] != ele[22][11];
    ele[22][2] != ele[22][12];
    ele[22][2] != ele[22][13];
    ele[22][2] != ele[22][14];
    ele[22][2] != ele[22][15];
    ele[22][2] != ele[22][16];
    ele[22][2] != ele[22][17];
    ele[22][2] != ele[22][18];
    ele[22][2] != ele[22][19];
    ele[22][2] != ele[22][20];
    ele[22][2] != ele[22][21];
    ele[22][2] != ele[22][22];
    ele[22][2] != ele[22][23];
    ele[22][2] != ele[22][24];
    ele[22][2] != ele[22][3];
    ele[22][2] != ele[22][4];
    ele[22][2] != ele[22][5];
    ele[22][2] != ele[22][6];
    ele[22][2] != ele[22][7];
    ele[22][2] != ele[22][8];
    ele[22][2] != ele[22][9];
    ele[22][2] != ele[23][0];
    ele[22][2] != ele[23][1];
    ele[22][2] != ele[23][2];
    ele[22][2] != ele[23][3];
    ele[22][2] != ele[23][4];
    ele[22][2] != ele[24][0];
    ele[22][2] != ele[24][1];
    ele[22][2] != ele[24][2];
    ele[22][2] != ele[24][3];
    ele[22][2] != ele[24][4];
    ele[22][20] != ele[22][21];
    ele[22][20] != ele[22][22];
    ele[22][20] != ele[22][23];
    ele[22][20] != ele[22][24];
    ele[22][20] != ele[23][20];
    ele[22][20] != ele[23][21];
    ele[22][20] != ele[23][22];
    ele[22][20] != ele[23][23];
    ele[22][20] != ele[23][24];
    ele[22][20] != ele[24][20];
    ele[22][20] != ele[24][21];
    ele[22][20] != ele[24][22];
    ele[22][20] != ele[24][23];
    ele[22][20] != ele[24][24];
    ele[22][21] != ele[22][22];
    ele[22][21] != ele[22][23];
    ele[22][21] != ele[22][24];
    ele[22][21] != ele[23][20];
    ele[22][21] != ele[23][21];
    ele[22][21] != ele[23][22];
    ele[22][21] != ele[23][23];
    ele[22][21] != ele[23][24];
    ele[22][21] != ele[24][20];
    ele[22][21] != ele[24][21];
    ele[22][21] != ele[24][22];
    ele[22][21] != ele[24][23];
    ele[22][21] != ele[24][24];
    ele[22][22] != ele[22][23];
    ele[22][22] != ele[22][24];
    ele[22][22] != ele[23][20];
    ele[22][22] != ele[23][21];
    ele[22][22] != ele[23][22];
    ele[22][22] != ele[23][23];
    ele[22][22] != ele[23][24];
    ele[22][22] != ele[24][20];
    ele[22][22] != ele[24][21];
    ele[22][22] != ele[24][22];
    ele[22][22] != ele[24][23];
    ele[22][22] != ele[24][24];
    ele[22][23] != ele[22][24];
    ele[22][23] != ele[23][20];
    ele[22][23] != ele[23][21];
    ele[22][23] != ele[23][22];
    ele[22][23] != ele[23][23];
    ele[22][23] != ele[23][24];
    ele[22][23] != ele[24][20];
    ele[22][23] != ele[24][21];
    ele[22][23] != ele[24][22];
    ele[22][23] != ele[24][23];
    ele[22][23] != ele[24][24];
    ele[22][24] != ele[23][20];
    ele[22][24] != ele[23][21];
    ele[22][24] != ele[23][22];
    ele[22][24] != ele[23][23];
    ele[22][24] != ele[23][24];
    ele[22][24] != ele[24][20];
    ele[22][24] != ele[24][21];
    ele[22][24] != ele[24][22];
    ele[22][24] != ele[24][23];
    ele[22][24] != ele[24][24];
    ele[22][3] != ele[22][10];
    ele[22][3] != ele[22][11];
    ele[22][3] != ele[22][12];
    ele[22][3] != ele[22][13];
    ele[22][3] != ele[22][14];
    ele[22][3] != ele[22][15];
    ele[22][3] != ele[22][16];
    ele[22][3] != ele[22][17];
    ele[22][3] != ele[22][18];
    ele[22][3] != ele[22][19];
    ele[22][3] != ele[22][20];
    ele[22][3] != ele[22][21];
    ele[22][3] != ele[22][22];
    ele[22][3] != ele[22][23];
    ele[22][3] != ele[22][24];
    ele[22][3] != ele[22][4];
    ele[22][3] != ele[22][5];
    ele[22][3] != ele[22][6];
    ele[22][3] != ele[22][7];
    ele[22][3] != ele[22][8];
    ele[22][3] != ele[22][9];
    ele[22][3] != ele[23][0];
    ele[22][3] != ele[23][1];
    ele[22][3] != ele[23][2];
    ele[22][3] != ele[23][3];
    ele[22][3] != ele[23][4];
    ele[22][3] != ele[24][0];
    ele[22][3] != ele[24][1];
    ele[22][3] != ele[24][2];
    ele[22][3] != ele[24][3];
    ele[22][3] != ele[24][4];
    ele[22][4] != ele[22][10];
    ele[22][4] != ele[22][11];
    ele[22][4] != ele[22][12];
    ele[22][4] != ele[22][13];
    ele[22][4] != ele[22][14];
    ele[22][4] != ele[22][15];
    ele[22][4] != ele[22][16];
    ele[22][4] != ele[22][17];
    ele[22][4] != ele[22][18];
    ele[22][4] != ele[22][19];
    ele[22][4] != ele[22][20];
    ele[22][4] != ele[22][21];
    ele[22][4] != ele[22][22];
    ele[22][4] != ele[22][23];
    ele[22][4] != ele[22][24];
    ele[22][4] != ele[22][5];
    ele[22][4] != ele[22][6];
    ele[22][4] != ele[22][7];
    ele[22][4] != ele[22][8];
    ele[22][4] != ele[22][9];
    ele[22][4] != ele[23][0];
    ele[22][4] != ele[23][1];
    ele[22][4] != ele[23][2];
    ele[22][4] != ele[23][3];
    ele[22][4] != ele[23][4];
    ele[22][4] != ele[24][0];
    ele[22][4] != ele[24][1];
    ele[22][4] != ele[24][2];
    ele[22][4] != ele[24][3];
    ele[22][4] != ele[24][4];
    ele[22][5] != ele[22][10];
    ele[22][5] != ele[22][11];
    ele[22][5] != ele[22][12];
    ele[22][5] != ele[22][13];
    ele[22][5] != ele[22][14];
    ele[22][5] != ele[22][15];
    ele[22][5] != ele[22][16];
    ele[22][5] != ele[22][17];
    ele[22][5] != ele[22][18];
    ele[22][5] != ele[22][19];
    ele[22][5] != ele[22][20];
    ele[22][5] != ele[22][21];
    ele[22][5] != ele[22][22];
    ele[22][5] != ele[22][23];
    ele[22][5] != ele[22][24];
    ele[22][5] != ele[22][6];
    ele[22][5] != ele[22][7];
    ele[22][5] != ele[22][8];
    ele[22][5] != ele[22][9];
    ele[22][5] != ele[23][5];
    ele[22][5] != ele[23][6];
    ele[22][5] != ele[23][7];
    ele[22][5] != ele[23][8];
    ele[22][5] != ele[23][9];
    ele[22][5] != ele[24][5];
    ele[22][5] != ele[24][6];
    ele[22][5] != ele[24][7];
    ele[22][5] != ele[24][8];
    ele[22][5] != ele[24][9];
    ele[22][6] != ele[22][10];
    ele[22][6] != ele[22][11];
    ele[22][6] != ele[22][12];
    ele[22][6] != ele[22][13];
    ele[22][6] != ele[22][14];
    ele[22][6] != ele[22][15];
    ele[22][6] != ele[22][16];
    ele[22][6] != ele[22][17];
    ele[22][6] != ele[22][18];
    ele[22][6] != ele[22][19];
    ele[22][6] != ele[22][20];
    ele[22][6] != ele[22][21];
    ele[22][6] != ele[22][22];
    ele[22][6] != ele[22][23];
    ele[22][6] != ele[22][24];
    ele[22][6] != ele[22][7];
    ele[22][6] != ele[22][8];
    ele[22][6] != ele[22][9];
    ele[22][6] != ele[23][5];
    ele[22][6] != ele[23][6];
    ele[22][6] != ele[23][7];
    ele[22][6] != ele[23][8];
    ele[22][6] != ele[23][9];
    ele[22][6] != ele[24][5];
    ele[22][6] != ele[24][6];
    ele[22][6] != ele[24][7];
    ele[22][6] != ele[24][8];
    ele[22][6] != ele[24][9];
    ele[22][7] != ele[22][10];
    ele[22][7] != ele[22][11];
    ele[22][7] != ele[22][12];
    ele[22][7] != ele[22][13];
    ele[22][7] != ele[22][14];
    ele[22][7] != ele[22][15];
    ele[22][7] != ele[22][16];
    ele[22][7] != ele[22][17];
    ele[22][7] != ele[22][18];
    ele[22][7] != ele[22][19];
    ele[22][7] != ele[22][20];
    ele[22][7] != ele[22][21];
    ele[22][7] != ele[22][22];
    ele[22][7] != ele[22][23];
    ele[22][7] != ele[22][24];
    ele[22][7] != ele[22][8];
    ele[22][7] != ele[22][9];
    ele[22][7] != ele[23][5];
    ele[22][7] != ele[23][6];
    ele[22][7] != ele[23][7];
    ele[22][7] != ele[23][8];
    ele[22][7] != ele[23][9];
    ele[22][7] != ele[24][5];
    ele[22][7] != ele[24][6];
    ele[22][7] != ele[24][7];
    ele[22][7] != ele[24][8];
    ele[22][7] != ele[24][9];
    ele[22][8] != ele[22][10];
    ele[22][8] != ele[22][11];
    ele[22][8] != ele[22][12];
    ele[22][8] != ele[22][13];
    ele[22][8] != ele[22][14];
    ele[22][8] != ele[22][15];
    ele[22][8] != ele[22][16];
    ele[22][8] != ele[22][17];
    ele[22][8] != ele[22][18];
    ele[22][8] != ele[22][19];
    ele[22][8] != ele[22][20];
    ele[22][8] != ele[22][21];
    ele[22][8] != ele[22][22];
    ele[22][8] != ele[22][23];
    ele[22][8] != ele[22][24];
    ele[22][8] != ele[22][9];
    ele[22][8] != ele[23][5];
    ele[22][8] != ele[23][6];
    ele[22][8] != ele[23][7];
    ele[22][8] != ele[23][8];
    ele[22][8] != ele[23][9];
    ele[22][8] != ele[24][5];
    ele[22][8] != ele[24][6];
    ele[22][8] != ele[24][7];
    ele[22][8] != ele[24][8];
    ele[22][8] != ele[24][9];
    ele[22][9] != ele[22][10];
    ele[22][9] != ele[22][11];
    ele[22][9] != ele[22][12];
    ele[22][9] != ele[22][13];
    ele[22][9] != ele[22][14];
    ele[22][9] != ele[22][15];
    ele[22][9] != ele[22][16];
    ele[22][9] != ele[22][17];
    ele[22][9] != ele[22][18];
    ele[22][9] != ele[22][19];
    ele[22][9] != ele[22][20];
    ele[22][9] != ele[22][21];
    ele[22][9] != ele[22][22];
    ele[22][9] != ele[22][23];
    ele[22][9] != ele[22][24];
    ele[22][9] != ele[23][5];
    ele[22][9] != ele[23][6];
    ele[22][9] != ele[23][7];
    ele[22][9] != ele[23][8];
    ele[22][9] != ele[23][9];
    ele[22][9] != ele[24][5];
    ele[22][9] != ele[24][6];
    ele[22][9] != ele[24][7];
    ele[22][9] != ele[24][8];
    ele[22][9] != ele[24][9];
    ele[23][0] != ele[23][1];
    ele[23][0] != ele[23][10];
    ele[23][0] != ele[23][11];
    ele[23][0] != ele[23][12];
    ele[23][0] != ele[23][13];
    ele[23][0] != ele[23][14];
    ele[23][0] != ele[23][15];
    ele[23][0] != ele[23][16];
    ele[23][0] != ele[23][17];
    ele[23][0] != ele[23][18];
    ele[23][0] != ele[23][19];
    ele[23][0] != ele[23][2];
    ele[23][0] != ele[23][20];
    ele[23][0] != ele[23][21];
    ele[23][0] != ele[23][22];
    ele[23][0] != ele[23][23];
    ele[23][0] != ele[23][24];
    ele[23][0] != ele[23][3];
    ele[23][0] != ele[23][4];
    ele[23][0] != ele[23][5];
    ele[23][0] != ele[23][6];
    ele[23][0] != ele[23][7];
    ele[23][0] != ele[23][8];
    ele[23][0] != ele[23][9];
    ele[23][0] != ele[24][0];
    ele[23][0] != ele[24][1];
    ele[23][0] != ele[24][2];
    ele[23][0] != ele[24][3];
    ele[23][0] != ele[24][4];
    ele[23][1] != ele[23][10];
    ele[23][1] != ele[23][11];
    ele[23][1] != ele[23][12];
    ele[23][1] != ele[23][13];
    ele[23][1] != ele[23][14];
    ele[23][1] != ele[23][15];
    ele[23][1] != ele[23][16];
    ele[23][1] != ele[23][17];
    ele[23][1] != ele[23][18];
    ele[23][1] != ele[23][19];
    ele[23][1] != ele[23][2];
    ele[23][1] != ele[23][20];
    ele[23][1] != ele[23][21];
    ele[23][1] != ele[23][22];
    ele[23][1] != ele[23][23];
    ele[23][1] != ele[23][24];
    ele[23][1] != ele[23][3];
    ele[23][1] != ele[23][4];
    ele[23][1] != ele[23][5];
    ele[23][1] != ele[23][6];
    ele[23][1] != ele[23][7];
    ele[23][1] != ele[23][8];
    ele[23][1] != ele[23][9];
    ele[23][1] != ele[24][0];
    ele[23][1] != ele[24][1];
    ele[23][1] != ele[24][2];
    ele[23][1] != ele[24][3];
    ele[23][1] != ele[24][4];
    ele[23][10] != ele[23][11];
    ele[23][10] != ele[23][12];
    ele[23][10] != ele[23][13];
    ele[23][10] != ele[23][14];
    ele[23][10] != ele[23][15];
    ele[23][10] != ele[23][16];
    ele[23][10] != ele[23][17];
    ele[23][10] != ele[23][18];
    ele[23][10] != ele[23][19];
    ele[23][10] != ele[23][20];
    ele[23][10] != ele[23][21];
    ele[23][10] != ele[23][22];
    ele[23][10] != ele[23][23];
    ele[23][10] != ele[23][24];
    ele[23][10] != ele[24][10];
    ele[23][10] != ele[24][11];
    ele[23][10] != ele[24][12];
    ele[23][10] != ele[24][13];
    ele[23][10] != ele[24][14];
    ele[23][11] != ele[23][12];
    ele[23][11] != ele[23][13];
    ele[23][11] != ele[23][14];
    ele[23][11] != ele[23][15];
    ele[23][11] != ele[23][16];
    ele[23][11] != ele[23][17];
    ele[23][11] != ele[23][18];
    ele[23][11] != ele[23][19];
    ele[23][11] != ele[23][20];
    ele[23][11] != ele[23][21];
    ele[23][11] != ele[23][22];
    ele[23][11] != ele[23][23];
    ele[23][11] != ele[23][24];
    ele[23][11] != ele[24][10];
    ele[23][11] != ele[24][11];
    ele[23][11] != ele[24][12];
    ele[23][11] != ele[24][13];
    ele[23][11] != ele[24][14];
    ele[23][12] != ele[23][13];
    ele[23][12] != ele[23][14];
    ele[23][12] != ele[23][15];
    ele[23][12] != ele[23][16];
    ele[23][12] != ele[23][17];
    ele[23][12] != ele[23][18];
    ele[23][12] != ele[23][19];
    ele[23][12] != ele[23][20];
    ele[23][12] != ele[23][21];
    ele[23][12] != ele[23][22];
    ele[23][12] != ele[23][23];
    ele[23][12] != ele[23][24];
    ele[23][12] != ele[24][10];
    ele[23][12] != ele[24][11];
    ele[23][12] != ele[24][12];
    ele[23][12] != ele[24][13];
    ele[23][12] != ele[24][14];
    ele[23][13] != ele[23][14];
    ele[23][13] != ele[23][15];
    ele[23][13] != ele[23][16];
    ele[23][13] != ele[23][17];
    ele[23][13] != ele[23][18];
    ele[23][13] != ele[23][19];
    ele[23][13] != ele[23][20];
    ele[23][13] != ele[23][21];
    ele[23][13] != ele[23][22];
    ele[23][13] != ele[23][23];
    ele[23][13] != ele[23][24];
    ele[23][13] != ele[24][10];
    ele[23][13] != ele[24][11];
    ele[23][13] != ele[24][12];
    ele[23][13] != ele[24][13];
    ele[23][13] != ele[24][14];
    ele[23][14] != ele[23][15];
    ele[23][14] != ele[23][16];
    ele[23][14] != ele[23][17];
    ele[23][14] != ele[23][18];
    ele[23][14] != ele[23][19];
    ele[23][14] != ele[23][20];
    ele[23][14] != ele[23][21];
    ele[23][14] != ele[23][22];
    ele[23][14] != ele[23][23];
    ele[23][14] != ele[23][24];
    ele[23][14] != ele[24][10];
    ele[23][14] != ele[24][11];
    ele[23][14] != ele[24][12];
    ele[23][14] != ele[24][13];
    ele[23][14] != ele[24][14];
    ele[23][15] != ele[23][16];
    ele[23][15] != ele[23][17];
    ele[23][15] != ele[23][18];
    ele[23][15] != ele[23][19];
    ele[23][15] != ele[23][20];
    ele[23][15] != ele[23][21];
    ele[23][15] != ele[23][22];
    ele[23][15] != ele[23][23];
    ele[23][15] != ele[23][24];
    ele[23][15] != ele[24][15];
    ele[23][15] != ele[24][16];
    ele[23][15] != ele[24][17];
    ele[23][15] != ele[24][18];
    ele[23][15] != ele[24][19];
    ele[23][16] != ele[23][17];
    ele[23][16] != ele[23][18];
    ele[23][16] != ele[23][19];
    ele[23][16] != ele[23][20];
    ele[23][16] != ele[23][21];
    ele[23][16] != ele[23][22];
    ele[23][16] != ele[23][23];
    ele[23][16] != ele[23][24];
    ele[23][16] != ele[24][15];
    ele[23][16] != ele[24][16];
    ele[23][16] != ele[24][17];
    ele[23][16] != ele[24][18];
    ele[23][16] != ele[24][19];
    ele[23][17] != ele[23][18];
    ele[23][17] != ele[23][19];
    ele[23][17] != ele[23][20];
    ele[23][17] != ele[23][21];
    ele[23][17] != ele[23][22];
    ele[23][17] != ele[23][23];
    ele[23][17] != ele[23][24];
    ele[23][17] != ele[24][15];
    ele[23][17] != ele[24][16];
    ele[23][17] != ele[24][17];
    ele[23][17] != ele[24][18];
    ele[23][17] != ele[24][19];
    ele[23][18] != ele[23][19];
    ele[23][18] != ele[23][20];
    ele[23][18] != ele[23][21];
    ele[23][18] != ele[23][22];
    ele[23][18] != ele[23][23];
    ele[23][18] != ele[23][24];
    ele[23][18] != ele[24][15];
    ele[23][18] != ele[24][16];
    ele[23][18] != ele[24][17];
    ele[23][18] != ele[24][18];
    ele[23][18] != ele[24][19];
    ele[23][19] != ele[23][20];
    ele[23][19] != ele[23][21];
    ele[23][19] != ele[23][22];
    ele[23][19] != ele[23][23];
    ele[23][19] != ele[23][24];
    ele[23][19] != ele[24][15];
    ele[23][19] != ele[24][16];
    ele[23][19] != ele[24][17];
    ele[23][19] != ele[24][18];
    ele[23][19] != ele[24][19];
    ele[23][2] != ele[23][10];
    ele[23][2] != ele[23][11];
    ele[23][2] != ele[23][12];
    ele[23][2] != ele[23][13];
    ele[23][2] != ele[23][14];
    ele[23][2] != ele[23][15];
    ele[23][2] != ele[23][16];
    ele[23][2] != ele[23][17];
    ele[23][2] != ele[23][18];
    ele[23][2] != ele[23][19];
    ele[23][2] != ele[23][20];
    ele[23][2] != ele[23][21];
    ele[23][2] != ele[23][22];
    ele[23][2] != ele[23][23];
    ele[23][2] != ele[23][24];
    ele[23][2] != ele[23][3];
    ele[23][2] != ele[23][4];
    ele[23][2] != ele[23][5];
    ele[23][2] != ele[23][6];
    ele[23][2] != ele[23][7];
    ele[23][2] != ele[23][8];
    ele[23][2] != ele[23][9];
    ele[23][2] != ele[24][0];
    ele[23][2] != ele[24][1];
    ele[23][2] != ele[24][2];
    ele[23][2] != ele[24][3];
    ele[23][2] != ele[24][4];
    ele[23][20] != ele[23][21];
    ele[23][20] != ele[23][22];
    ele[23][20] != ele[23][23];
    ele[23][20] != ele[23][24];
    ele[23][20] != ele[24][20];
    ele[23][20] != ele[24][21];
    ele[23][20] != ele[24][22];
    ele[23][20] != ele[24][23];
    ele[23][20] != ele[24][24];
    ele[23][21] != ele[23][22];
    ele[23][21] != ele[23][23];
    ele[23][21] != ele[23][24];
    ele[23][21] != ele[24][20];
    ele[23][21] != ele[24][21];
    ele[23][21] != ele[24][22];
    ele[23][21] != ele[24][23];
    ele[23][21] != ele[24][24];
    ele[23][22] != ele[23][23];
    ele[23][22] != ele[23][24];
    ele[23][22] != ele[24][20];
    ele[23][22] != ele[24][21];
    ele[23][22] != ele[24][22];
    ele[23][22] != ele[24][23];
    ele[23][22] != ele[24][24];
    ele[23][23] != ele[23][24];
    ele[23][23] != ele[24][20];
    ele[23][23] != ele[24][21];
    ele[23][23] != ele[24][22];
    ele[23][23] != ele[24][23];
    ele[23][23] != ele[24][24];
    ele[23][24] != ele[24][20];
    ele[23][24] != ele[24][21];
    ele[23][24] != ele[24][22];
    ele[23][24] != ele[24][23];
    ele[23][24] != ele[24][24];
    ele[23][3] != ele[23][10];
    ele[23][3] != ele[23][11];
    ele[23][3] != ele[23][12];
    ele[23][3] != ele[23][13];
    ele[23][3] != ele[23][14];
    ele[23][3] != ele[23][15];
    ele[23][3] != ele[23][16];
    ele[23][3] != ele[23][17];
    ele[23][3] != ele[23][18];
    ele[23][3] != ele[23][19];
    ele[23][3] != ele[23][20];
    ele[23][3] != ele[23][21];
    ele[23][3] != ele[23][22];
    ele[23][3] != ele[23][23];
    ele[23][3] != ele[23][24];
    ele[23][3] != ele[23][4];
    ele[23][3] != ele[23][5];
    ele[23][3] != ele[23][6];
    ele[23][3] != ele[23][7];
    ele[23][3] != ele[23][8];
    ele[23][3] != ele[23][9];
    ele[23][3] != ele[24][0];
    ele[23][3] != ele[24][1];
    ele[23][3] != ele[24][2];
    ele[23][3] != ele[24][3];
    ele[23][3] != ele[24][4];
    ele[23][4] != ele[23][10];
    ele[23][4] != ele[23][11];
    ele[23][4] != ele[23][12];
    ele[23][4] != ele[23][13];
    ele[23][4] != ele[23][14];
    ele[23][4] != ele[23][15];
    ele[23][4] != ele[23][16];
    ele[23][4] != ele[23][17];
    ele[23][4] != ele[23][18];
    ele[23][4] != ele[23][19];
    ele[23][4] != ele[23][20];
    ele[23][4] != ele[23][21];
    ele[23][4] != ele[23][22];
    ele[23][4] != ele[23][23];
    ele[23][4] != ele[23][24];
    ele[23][4] != ele[23][5];
    ele[23][4] != ele[23][6];
    ele[23][4] != ele[23][7];
    ele[23][4] != ele[23][8];
    ele[23][4] != ele[23][9];
    ele[23][4] != ele[24][0];
    ele[23][4] != ele[24][1];
    ele[23][4] != ele[24][2];
    ele[23][4] != ele[24][3];
    ele[23][4] != ele[24][4];
    ele[23][5] != ele[23][10];
    ele[23][5] != ele[23][11];
    ele[23][5] != ele[23][12];
    ele[23][5] != ele[23][13];
    ele[23][5] != ele[23][14];
    ele[23][5] != ele[23][15];
    ele[23][5] != ele[23][16];
    ele[23][5] != ele[23][17];
    ele[23][5] != ele[23][18];
    ele[23][5] != ele[23][19];
    ele[23][5] != ele[23][20];
    ele[23][5] != ele[23][21];
    ele[23][5] != ele[23][22];
    ele[23][5] != ele[23][23];
    ele[23][5] != ele[23][24];
    ele[23][5] != ele[23][6];
    ele[23][5] != ele[23][7];
    ele[23][5] != ele[23][8];
    ele[23][5] != ele[23][9];
    ele[23][5] != ele[24][5];
    ele[23][5] != ele[24][6];
    ele[23][5] != ele[24][7];
    ele[23][5] != ele[24][8];
    ele[23][5] != ele[24][9];
    ele[23][6] != ele[23][10];
    ele[23][6] != ele[23][11];
    ele[23][6] != ele[23][12];
    ele[23][6] != ele[23][13];
    ele[23][6] != ele[23][14];
    ele[23][6] != ele[23][15];
    ele[23][6] != ele[23][16];
    ele[23][6] != ele[23][17];
    ele[23][6] != ele[23][18];
    ele[23][6] != ele[23][19];
    ele[23][6] != ele[23][20];
    ele[23][6] != ele[23][21];
    ele[23][6] != ele[23][22];
    ele[23][6] != ele[23][23];
    ele[23][6] != ele[23][24];
    ele[23][6] != ele[23][7];
    ele[23][6] != ele[23][8];
    ele[23][6] != ele[23][9];
    ele[23][6] != ele[24][5];
    ele[23][6] != ele[24][6];
    ele[23][6] != ele[24][7];
    ele[23][6] != ele[24][8];
    ele[23][6] != ele[24][9];
    ele[23][7] != ele[23][10];
    ele[23][7] != ele[23][11];
    ele[23][7] != ele[23][12];
    ele[23][7] != ele[23][13];
    ele[23][7] != ele[23][14];
    ele[23][7] != ele[23][15];
    ele[23][7] != ele[23][16];
    ele[23][7] != ele[23][17];
    ele[23][7] != ele[23][18];
    ele[23][7] != ele[23][19];
    ele[23][7] != ele[23][20];
    ele[23][7] != ele[23][21];
    ele[23][7] != ele[23][22];
    ele[23][7] != ele[23][23];
    ele[23][7] != ele[23][24];
    ele[23][7] != ele[23][8];
    ele[23][7] != ele[23][9];
    ele[23][7] != ele[24][5];
    ele[23][7] != ele[24][6];
    ele[23][7] != ele[24][7];
    ele[23][7] != ele[24][8];
    ele[23][7] != ele[24][9];
    ele[23][8] != ele[23][10];
    ele[23][8] != ele[23][11];
    ele[23][8] != ele[23][12];
    ele[23][8] != ele[23][13];
    ele[23][8] != ele[23][14];
    ele[23][8] != ele[23][15];
    ele[23][8] != ele[23][16];
    ele[23][8] != ele[23][17];
    ele[23][8] != ele[23][18];
    ele[23][8] != ele[23][19];
    ele[23][8] != ele[23][20];
    ele[23][8] != ele[23][21];
    ele[23][8] != ele[23][22];
    ele[23][8] != ele[23][23];
    ele[23][8] != ele[23][24];
    ele[23][8] != ele[23][9];
    ele[23][8] != ele[24][5];
    ele[23][8] != ele[24][6];
    ele[23][8] != ele[24][7];
    ele[23][8] != ele[24][8];
    ele[23][8] != ele[24][9];
    ele[23][9] != ele[23][10];
    ele[23][9] != ele[23][11];
    ele[23][9] != ele[23][12];
    ele[23][9] != ele[23][13];
    ele[23][9] != ele[23][14];
    ele[23][9] != ele[23][15];
    ele[23][9] != ele[23][16];
    ele[23][9] != ele[23][17];
    ele[23][9] != ele[23][18];
    ele[23][9] != ele[23][19];
    ele[23][9] != ele[23][20];
    ele[23][9] != ele[23][21];
    ele[23][9] != ele[23][22];
    ele[23][9] != ele[23][23];
    ele[23][9] != ele[23][24];
    ele[23][9] != ele[24][5];
    ele[23][9] != ele[24][6];
    ele[23][9] != ele[24][7];
    ele[23][9] != ele[24][8];
    ele[23][9] != ele[24][9];
    ele[24][0] != ele[24][1];
    ele[24][0] != ele[24][10];
    ele[24][0] != ele[24][11];
    ele[24][0] != ele[24][12];
    ele[24][0] != ele[24][13];
    ele[24][0] != ele[24][14];
    ele[24][0] != ele[24][15];
    ele[24][0] != ele[24][16];
    ele[24][0] != ele[24][17];
    ele[24][0] != ele[24][18];
    ele[24][0] != ele[24][19];
    ele[24][0] != ele[24][2];
    ele[24][0] != ele[24][20];
    ele[24][0] != ele[24][21];
    ele[24][0] != ele[24][22];
    ele[24][0] != ele[24][23];
    ele[24][0] != ele[24][24];
    ele[24][0] != ele[24][3];
    ele[24][0] != ele[24][4];
    ele[24][0] != ele[24][5];
    ele[24][0] != ele[24][6];
    ele[24][0] != ele[24][7];
    ele[24][0] != ele[24][8];
    ele[24][0] != ele[24][9];
    ele[24][1] != ele[24][10];
    ele[24][1] != ele[24][11];
    ele[24][1] != ele[24][12];
    ele[24][1] != ele[24][13];
    ele[24][1] != ele[24][14];
    ele[24][1] != ele[24][15];
    ele[24][1] != ele[24][16];
    ele[24][1] != ele[24][17];
    ele[24][1] != ele[24][18];
    ele[24][1] != ele[24][19];
    ele[24][1] != ele[24][2];
    ele[24][1] != ele[24][20];
    ele[24][1] != ele[24][21];
    ele[24][1] != ele[24][22];
    ele[24][1] != ele[24][23];
    ele[24][1] != ele[24][24];
    ele[24][1] != ele[24][3];
    ele[24][1] != ele[24][4];
    ele[24][1] != ele[24][5];
    ele[24][1] != ele[24][6];
    ele[24][1] != ele[24][7];
    ele[24][1] != ele[24][8];
    ele[24][1] != ele[24][9];
    ele[24][10] != ele[24][11];
    ele[24][10] != ele[24][12];
    ele[24][10] != ele[24][13];
    ele[24][10] != ele[24][14];
    ele[24][10] != ele[24][15];
    ele[24][10] != ele[24][16];
    ele[24][10] != ele[24][17];
    ele[24][10] != ele[24][18];
    ele[24][10] != ele[24][19];
    ele[24][10] != ele[24][20];
    ele[24][10] != ele[24][21];
    ele[24][10] != ele[24][22];
    ele[24][10] != ele[24][23];
    ele[24][10] != ele[24][24];
    ele[24][11] != ele[24][12];
    ele[24][11] != ele[24][13];
    ele[24][11] != ele[24][14];
    ele[24][11] != ele[24][15];
    ele[24][11] != ele[24][16];
    ele[24][11] != ele[24][17];
    ele[24][11] != ele[24][18];
    ele[24][11] != ele[24][19];
    ele[24][11] != ele[24][20];
    ele[24][11] != ele[24][21];
    ele[24][11] != ele[24][22];
    ele[24][11] != ele[24][23];
    ele[24][11] != ele[24][24];
    ele[24][12] != ele[24][13];
    ele[24][12] != ele[24][14];
    ele[24][12] != ele[24][15];
    ele[24][12] != ele[24][16];
    ele[24][12] != ele[24][17];
    ele[24][12] != ele[24][18];
    ele[24][12] != ele[24][19];
    ele[24][12] != ele[24][20];
    ele[24][12] != ele[24][21];
    ele[24][12] != ele[24][22];
    ele[24][12] != ele[24][23];
    ele[24][12] != ele[24][24];
    ele[24][13] != ele[24][14];
    ele[24][13] != ele[24][15];
    ele[24][13] != ele[24][16];
    ele[24][13] != ele[24][17];
    ele[24][13] != ele[24][18];
    ele[24][13] != ele[24][19];
    ele[24][13] != ele[24][20];
    ele[24][13] != ele[24][21];
    ele[24][13] != ele[24][22];
    ele[24][13] != ele[24][23];
    ele[24][13] != ele[24][24];
    ele[24][14] != ele[24][15];
    ele[24][14] != ele[24][16];
    ele[24][14] != ele[24][17];
    ele[24][14] != ele[24][18];
    ele[24][14] != ele[24][19];
    ele[24][14] != ele[24][20];
    ele[24][14] != ele[24][21];
    ele[24][14] != ele[24][22];
    ele[24][14] != ele[24][23];
    ele[24][14] != ele[24][24];
    ele[24][15] != ele[24][16];
    ele[24][15] != ele[24][17];
    ele[24][15] != ele[24][18];
    ele[24][15] != ele[24][19];
    ele[24][15] != ele[24][20];
    ele[24][15] != ele[24][21];
    ele[24][15] != ele[24][22];
    ele[24][15] != ele[24][23];
    ele[24][15] != ele[24][24];
    ele[24][16] != ele[24][17];
    ele[24][16] != ele[24][18];
    ele[24][16] != ele[24][19];
    ele[24][16] != ele[24][20];
    ele[24][16] != ele[24][21];
    ele[24][16] != ele[24][22];
    ele[24][16] != ele[24][23];
    ele[24][16] != ele[24][24];
    ele[24][17] != ele[24][18];
    ele[24][17] != ele[24][19];
    ele[24][17] != ele[24][20];
    ele[24][17] != ele[24][21];
    ele[24][17] != ele[24][22];
    ele[24][17] != ele[24][23];
    ele[24][17] != ele[24][24];
    ele[24][18] != ele[24][19];
    ele[24][18] != ele[24][20];
    ele[24][18] != ele[24][21];
    ele[24][18] != ele[24][22];
    ele[24][18] != ele[24][23];
    ele[24][18] != ele[24][24];
    ele[24][19] != ele[24][20];
    ele[24][19] != ele[24][21];
    ele[24][19] != ele[24][22];
    ele[24][19] != ele[24][23];
    ele[24][19] != ele[24][24];
    ele[24][2] != ele[24][10];
    ele[24][2] != ele[24][11];
    ele[24][2] != ele[24][12];
    ele[24][2] != ele[24][13];
    ele[24][2] != ele[24][14];
    ele[24][2] != ele[24][15];
    ele[24][2] != ele[24][16];
    ele[24][2] != ele[24][17];
    ele[24][2] != ele[24][18];
    ele[24][2] != ele[24][19];
    ele[24][2] != ele[24][20];
    ele[24][2] != ele[24][21];
    ele[24][2] != ele[24][22];
    ele[24][2] != ele[24][23];
    ele[24][2] != ele[24][24];
    ele[24][2] != ele[24][3];
    ele[24][2] != ele[24][4];
    ele[24][2] != ele[24][5];
    ele[24][2] != ele[24][6];
    ele[24][2] != ele[24][7];
    ele[24][2] != ele[24][8];
    ele[24][2] != ele[24][9];
    ele[24][20] != ele[24][21];
    ele[24][20] != ele[24][22];
    ele[24][20] != ele[24][23];
    ele[24][20] != ele[24][24];
    ele[24][21] != ele[24][22];
    ele[24][21] != ele[24][23];
    ele[24][21] != ele[24][24];
    ele[24][22] != ele[24][23];
    ele[24][22] != ele[24][24];
    ele[24][23] != ele[24][24];
    ele[24][3] != ele[24][10];
    ele[24][3] != ele[24][11];
    ele[24][3] != ele[24][12];
    ele[24][3] != ele[24][13];
    ele[24][3] != ele[24][14];
    ele[24][3] != ele[24][15];
    ele[24][3] != ele[24][16];
    ele[24][3] != ele[24][17];
    ele[24][3] != ele[24][18];
    ele[24][3] != ele[24][19];
    ele[24][3] != ele[24][20];
    ele[24][3] != ele[24][21];
    ele[24][3] != ele[24][22];
    ele[24][3] != ele[24][23];
    ele[24][3] != ele[24][24];
    ele[24][3] != ele[24][4];
    ele[24][3] != ele[24][5];
    ele[24][3] != ele[24][6];
    ele[24][3] != ele[24][7];
    ele[24][3] != ele[24][8];
    ele[24][3] != ele[24][9];
    ele[24][4] != ele[24][10];
    ele[24][4] != ele[24][11];
    ele[24][4] != ele[24][12];
    ele[24][4] != ele[24][13];
    ele[24][4] != ele[24][14];
    ele[24][4] != ele[24][15];
    ele[24][4] != ele[24][16];
    ele[24][4] != ele[24][17];
    ele[24][4] != ele[24][18];
    ele[24][4] != ele[24][19];
    ele[24][4] != ele[24][20];
    ele[24][4] != ele[24][21];
    ele[24][4] != ele[24][22];
    ele[24][4] != ele[24][23];
    ele[24][4] != ele[24][24];
    ele[24][4] != ele[24][5];
    ele[24][4] != ele[24][6];
    ele[24][4] != ele[24][7];
    ele[24][4] != ele[24][8];
    ele[24][4] != ele[24][9];
    ele[24][5] != ele[24][10];
    ele[24][5] != ele[24][11];
    ele[24][5] != ele[24][12];
    ele[24][5] != ele[24][13];
    ele[24][5] != ele[24][14];
    ele[24][5] != ele[24][15];
    ele[24][5] != ele[24][16];
    ele[24][5] != ele[24][17];
    ele[24][5] != ele[24][18];
    ele[24][5] != ele[24][19];
    ele[24][5] != ele[24][20];
    ele[24][5] != ele[24][21];
    ele[24][5] != ele[24][22];
    ele[24][5] != ele[24][23];
    ele[24][5] != ele[24][24];
    ele[24][5] != ele[24][6];
    ele[24][5] != ele[24][7];
    ele[24][5] != ele[24][8];
    ele[24][5] != ele[24][9];
    ele[24][6] != ele[24][10];
    ele[24][6] != ele[24][11];
    ele[24][6] != ele[24][12];
    ele[24][6] != ele[24][13];
    ele[24][6] != ele[24][14];
    ele[24][6] != ele[24][15];
    ele[24][6] != ele[24][16];
    ele[24][6] != ele[24][17];
    ele[24][6] != ele[24][18];
    ele[24][6] != ele[24][19];
    ele[24][6] != ele[24][20];
    ele[24][6] != ele[24][21];
    ele[24][6] != ele[24][22];
    ele[24][6] != ele[24][23];
    ele[24][6] != ele[24][24];
    ele[24][6] != ele[24][7];
    ele[24][6] != ele[24][8];
    ele[24][6] != ele[24][9];
    ele[24][7] != ele[24][10];
    ele[24][7] != ele[24][11];
    ele[24][7] != ele[24][12];
    ele[24][7] != ele[24][13];
    ele[24][7] != ele[24][14];
    ele[24][7] != ele[24][15];
    ele[24][7] != ele[24][16];
    ele[24][7] != ele[24][17];
    ele[24][7] != ele[24][18];
    ele[24][7] != ele[24][19];
    ele[24][7] != ele[24][20];
    ele[24][7] != ele[24][21];
    ele[24][7] != ele[24][22];
    ele[24][7] != ele[24][23];
    ele[24][7] != ele[24][24];
    ele[24][7] != ele[24][8];
    ele[24][7] != ele[24][9];
    ele[24][8] != ele[24][10];
    ele[24][8] != ele[24][11];
    ele[24][8] != ele[24][12];
    ele[24][8] != ele[24][13];
    ele[24][8] != ele[24][14];
    ele[24][8] != ele[24][15];
    ele[24][8] != ele[24][16];
    ele[24][8] != ele[24][17];
    ele[24][8] != ele[24][18];
    ele[24][8] != ele[24][19];
    ele[24][8] != ele[24][20];
    ele[24][8] != ele[24][21];
    ele[24][8] != ele[24][22];
    ele[24][8] != ele[24][23];
    ele[24][8] != ele[24][24];
    ele[24][8] != ele[24][9];
    ele[24][9] != ele[24][10];
    ele[24][9] != ele[24][11];
    ele[24][9] != ele[24][12];
    ele[24][9] != ele[24][13];
    ele[24][9] != ele[24][14];
    ele[24][9] != ele[24][15];
    ele[24][9] != ele[24][16];
    ele[24][9] != ele[24][17];
    ele[24][9] != ele[24][18];
    ele[24][9] != ele[24][19];
    ele[24][9] != ele[24][20];
    ele[24][9] != ele[24][21];
    ele[24][9] != ele[24][22];
    ele[24][9] != ele[24][23];
    ele[24][9] != ele[24][24];
    ele[3][0] != ele[10][0];
    ele[3][0] != ele[11][0];
    ele[3][0] != ele[12][0];
    ele[3][0] != ele[13][0];
    ele[3][0] != ele[14][0];
    ele[3][0] != ele[15][0];
    ele[3][0] != ele[16][0];
    ele[3][0] != ele[17][0];
    ele[3][0] != ele[18][0];
    ele[3][0] != ele[19][0];
    ele[3][0] != ele[20][0];
    ele[3][0] != ele[21][0];
    ele[3][0] != ele[22][0];
    ele[3][0] != ele[23][0];
    ele[3][0] != ele[24][0];
    ele[3][0] != ele[3][1];
    ele[3][0] != ele[3][10];
    ele[3][0] != ele[3][11];
    ele[3][0] != ele[3][12];
    ele[3][0] != ele[3][13];
    ele[3][0] != ele[3][14];
    ele[3][0] != ele[3][15];
    ele[3][0] != ele[3][16];
    ele[3][0] != ele[3][17];
    ele[3][0] != ele[3][18];
    ele[3][0] != ele[3][19];
    ele[3][0] != ele[3][2];
    ele[3][0] != ele[3][20];
    ele[3][0] != ele[3][21];
    ele[3][0] != ele[3][22];
    ele[3][0] != ele[3][23];
    ele[3][0] != ele[3][24];
    ele[3][0] != ele[3][3];
    ele[3][0] != ele[3][4];
    ele[3][0] != ele[3][5];
    ele[3][0] != ele[3][6];
    ele[3][0] != ele[3][7];
    ele[3][0] != ele[3][8];
    ele[3][0] != ele[3][9];
    ele[3][0] != ele[4][0];
    ele[3][0] != ele[4][1];
    ele[3][0] != ele[4][2];
    ele[3][0] != ele[4][3];
    ele[3][0] != ele[4][4];
    ele[3][0] != ele[5][0];
    ele[3][0] != ele[6][0];
    ele[3][0] != ele[7][0];
    ele[3][0] != ele[8][0];
    ele[3][0] != ele[9][0];
    ele[3][1] != ele[10][1];
    ele[3][1] != ele[11][1];
    ele[3][1] != ele[12][1];
    ele[3][1] != ele[13][1];
    ele[3][1] != ele[14][1];
    ele[3][1] != ele[15][1];
    ele[3][1] != ele[16][1];
    ele[3][1] != ele[17][1];
    ele[3][1] != ele[18][1];
    ele[3][1] != ele[19][1];
    ele[3][1] != ele[20][1];
    ele[3][1] != ele[21][1];
    ele[3][1] != ele[22][1];
    ele[3][1] != ele[23][1];
    ele[3][1] != ele[24][1];
    ele[3][1] != ele[3][10];
    ele[3][1] != ele[3][11];
    ele[3][1] != ele[3][12];
    ele[3][1] != ele[3][13];
    ele[3][1] != ele[3][14];
    ele[3][1] != ele[3][15];
    ele[3][1] != ele[3][16];
    ele[3][1] != ele[3][17];
    ele[3][1] != ele[3][18];
    ele[3][1] != ele[3][19];
    ele[3][1] != ele[3][2];
    ele[3][1] != ele[3][20];
    ele[3][1] != ele[3][21];
    ele[3][1] != ele[3][22];
    ele[3][1] != ele[3][23];
    ele[3][1] != ele[3][24];
    ele[3][1] != ele[3][3];
    ele[3][1] != ele[3][4];
    ele[3][1] != ele[3][5];
    ele[3][1] != ele[3][6];
    ele[3][1] != ele[3][7];
    ele[3][1] != ele[3][8];
    ele[3][1] != ele[3][9];
    ele[3][1] != ele[4][0];
    ele[3][1] != ele[4][1];
    ele[3][1] != ele[4][2];
    ele[3][1] != ele[4][3];
    ele[3][1] != ele[4][4];
    ele[3][1] != ele[5][1];
    ele[3][1] != ele[6][1];
    ele[3][1] != ele[7][1];
    ele[3][1] != ele[8][1];
    ele[3][1] != ele[9][1];
    ele[3][10] != ele[10][10];
    ele[3][10] != ele[11][10];
    ele[3][10] != ele[12][10];
    ele[3][10] != ele[13][10];
    ele[3][10] != ele[14][10];
    ele[3][10] != ele[15][10];
    ele[3][10] != ele[16][10];
    ele[3][10] != ele[17][10];
    ele[3][10] != ele[18][10];
    ele[3][10] != ele[19][10];
    ele[3][10] != ele[20][10];
    ele[3][10] != ele[21][10];
    ele[3][10] != ele[22][10];
    ele[3][10] != ele[23][10];
    ele[3][10] != ele[24][10];
    ele[3][10] != ele[3][11];
    ele[3][10] != ele[3][12];
    ele[3][10] != ele[3][13];
    ele[3][10] != ele[3][14];
    ele[3][10] != ele[3][15];
    ele[3][10] != ele[3][16];
    ele[3][10] != ele[3][17];
    ele[3][10] != ele[3][18];
    ele[3][10] != ele[3][19];
    ele[3][10] != ele[3][20];
    ele[3][10] != ele[3][21];
    ele[3][10] != ele[3][22];
    ele[3][10] != ele[3][23];
    ele[3][10] != ele[3][24];
    ele[3][10] != ele[4][10];
    ele[3][10] != ele[4][11];
    ele[3][10] != ele[4][12];
    ele[3][10] != ele[4][13];
    ele[3][10] != ele[4][14];
    ele[3][10] != ele[5][10];
    ele[3][10] != ele[6][10];
    ele[3][10] != ele[7][10];
    ele[3][10] != ele[8][10];
    ele[3][10] != ele[9][10];
    ele[3][11] != ele[10][11];
    ele[3][11] != ele[11][11];
    ele[3][11] != ele[12][11];
    ele[3][11] != ele[13][11];
    ele[3][11] != ele[14][11];
    ele[3][11] != ele[15][11];
    ele[3][11] != ele[16][11];
    ele[3][11] != ele[17][11];
    ele[3][11] != ele[18][11];
    ele[3][11] != ele[19][11];
    ele[3][11] != ele[20][11];
    ele[3][11] != ele[21][11];
    ele[3][11] != ele[22][11];
    ele[3][11] != ele[23][11];
    ele[3][11] != ele[24][11];
    ele[3][11] != ele[3][12];
    ele[3][11] != ele[3][13];
    ele[3][11] != ele[3][14];
    ele[3][11] != ele[3][15];
    ele[3][11] != ele[3][16];
    ele[3][11] != ele[3][17];
    ele[3][11] != ele[3][18];
    ele[3][11] != ele[3][19];
    ele[3][11] != ele[3][20];
    ele[3][11] != ele[3][21];
    ele[3][11] != ele[3][22];
    ele[3][11] != ele[3][23];
    ele[3][11] != ele[3][24];
    ele[3][11] != ele[4][10];
    ele[3][11] != ele[4][11];
    ele[3][11] != ele[4][12];
    ele[3][11] != ele[4][13];
    ele[3][11] != ele[4][14];
    ele[3][11] != ele[5][11];
    ele[3][11] != ele[6][11];
    ele[3][11] != ele[7][11];
    ele[3][11] != ele[8][11];
    ele[3][11] != ele[9][11];
    ele[3][12] != ele[10][12];
    ele[3][12] != ele[11][12];
    ele[3][12] != ele[12][12];
    ele[3][12] != ele[13][12];
    ele[3][12] != ele[14][12];
    ele[3][12] != ele[15][12];
    ele[3][12] != ele[16][12];
    ele[3][12] != ele[17][12];
    ele[3][12] != ele[18][12];
    ele[3][12] != ele[19][12];
    ele[3][12] != ele[20][12];
    ele[3][12] != ele[21][12];
    ele[3][12] != ele[22][12];
    ele[3][12] != ele[23][12];
    ele[3][12] != ele[24][12];
    ele[3][12] != ele[3][13];
    ele[3][12] != ele[3][14];
    ele[3][12] != ele[3][15];
    ele[3][12] != ele[3][16];
    ele[3][12] != ele[3][17];
    ele[3][12] != ele[3][18];
    ele[3][12] != ele[3][19];
    ele[3][12] != ele[3][20];
    ele[3][12] != ele[3][21];
    ele[3][12] != ele[3][22];
    ele[3][12] != ele[3][23];
    ele[3][12] != ele[3][24];
    ele[3][12] != ele[4][10];
    ele[3][12] != ele[4][11];
    ele[3][12] != ele[4][12];
    ele[3][12] != ele[4][13];
    ele[3][12] != ele[4][14];
    ele[3][12] != ele[5][12];
    ele[3][12] != ele[6][12];
    ele[3][12] != ele[7][12];
    ele[3][12] != ele[8][12];
    ele[3][12] != ele[9][12];
    ele[3][13] != ele[10][13];
    ele[3][13] != ele[11][13];
    ele[3][13] != ele[12][13];
    ele[3][13] != ele[13][13];
    ele[3][13] != ele[14][13];
    ele[3][13] != ele[15][13];
    ele[3][13] != ele[16][13];
    ele[3][13] != ele[17][13];
    ele[3][13] != ele[18][13];
    ele[3][13] != ele[19][13];
    ele[3][13] != ele[20][13];
    ele[3][13] != ele[21][13];
    ele[3][13] != ele[22][13];
    ele[3][13] != ele[23][13];
    ele[3][13] != ele[24][13];
    ele[3][13] != ele[3][14];
    ele[3][13] != ele[3][15];
    ele[3][13] != ele[3][16];
    ele[3][13] != ele[3][17];
    ele[3][13] != ele[3][18];
    ele[3][13] != ele[3][19];
    ele[3][13] != ele[3][20];
    ele[3][13] != ele[3][21];
    ele[3][13] != ele[3][22];
    ele[3][13] != ele[3][23];
    ele[3][13] != ele[3][24];
    ele[3][13] != ele[4][10];
    ele[3][13] != ele[4][11];
    ele[3][13] != ele[4][12];
    ele[3][13] != ele[4][13];
    ele[3][13] != ele[4][14];
    ele[3][13] != ele[5][13];
    ele[3][13] != ele[6][13];
    ele[3][13] != ele[7][13];
    ele[3][13] != ele[8][13];
    ele[3][13] != ele[9][13];
    ele[3][14] != ele[10][14];
    ele[3][14] != ele[11][14];
    ele[3][14] != ele[12][14];
    ele[3][14] != ele[13][14];
    ele[3][14] != ele[14][14];
    ele[3][14] != ele[15][14];
    ele[3][14] != ele[16][14];
    ele[3][14] != ele[17][14];
    ele[3][14] != ele[18][14];
    ele[3][14] != ele[19][14];
    ele[3][14] != ele[20][14];
    ele[3][14] != ele[21][14];
    ele[3][14] != ele[22][14];
    ele[3][14] != ele[23][14];
    ele[3][14] != ele[24][14];
    ele[3][14] != ele[3][15];
    ele[3][14] != ele[3][16];
    ele[3][14] != ele[3][17];
    ele[3][14] != ele[3][18];
    ele[3][14] != ele[3][19];
    ele[3][14] != ele[3][20];
    ele[3][14] != ele[3][21];
    ele[3][14] != ele[3][22];
    ele[3][14] != ele[3][23];
    ele[3][14] != ele[3][24];
    ele[3][14] != ele[4][10];
    ele[3][14] != ele[4][11];
    ele[3][14] != ele[4][12];
    ele[3][14] != ele[4][13];
    ele[3][14] != ele[4][14];
    ele[3][14] != ele[5][14];
    ele[3][14] != ele[6][14];
    ele[3][14] != ele[7][14];
    ele[3][14] != ele[8][14];
    ele[3][14] != ele[9][14];
    ele[3][15] != ele[10][15];
    ele[3][15] != ele[11][15];
    ele[3][15] != ele[12][15];
    ele[3][15] != ele[13][15];
    ele[3][15] != ele[14][15];
    ele[3][15] != ele[15][15];
    ele[3][15] != ele[16][15];
    ele[3][15] != ele[17][15];
    ele[3][15] != ele[18][15];
    ele[3][15] != ele[19][15];
    ele[3][15] != ele[20][15];
    ele[3][15] != ele[21][15];
    ele[3][15] != ele[22][15];
    ele[3][15] != ele[23][15];
    ele[3][15] != ele[24][15];
    ele[3][15] != ele[3][16];
    ele[3][15] != ele[3][17];
    ele[3][15] != ele[3][18];
    ele[3][15] != ele[3][19];
    ele[3][15] != ele[3][20];
    ele[3][15] != ele[3][21];
    ele[3][15] != ele[3][22];
    ele[3][15] != ele[3][23];
    ele[3][15] != ele[3][24];
    ele[3][15] != ele[4][15];
    ele[3][15] != ele[4][16];
    ele[3][15] != ele[4][17];
    ele[3][15] != ele[4][18];
    ele[3][15] != ele[4][19];
    ele[3][15] != ele[5][15];
    ele[3][15] != ele[6][15];
    ele[3][15] != ele[7][15];
    ele[3][15] != ele[8][15];
    ele[3][15] != ele[9][15];
    ele[3][16] != ele[10][16];
    ele[3][16] != ele[11][16];
    ele[3][16] != ele[12][16];
    ele[3][16] != ele[13][16];
    ele[3][16] != ele[14][16];
    ele[3][16] != ele[15][16];
    ele[3][16] != ele[16][16];
    ele[3][16] != ele[17][16];
    ele[3][16] != ele[18][16];
    ele[3][16] != ele[19][16];
    ele[3][16] != ele[20][16];
    ele[3][16] != ele[21][16];
    ele[3][16] != ele[22][16];
    ele[3][16] != ele[23][16];
    ele[3][16] != ele[24][16];
    ele[3][16] != ele[3][17];
    ele[3][16] != ele[3][18];
    ele[3][16] != ele[3][19];
    ele[3][16] != ele[3][20];
    ele[3][16] != ele[3][21];
    ele[3][16] != ele[3][22];
    ele[3][16] != ele[3][23];
    ele[3][16] != ele[3][24];
    ele[3][16] != ele[4][15];
    ele[3][16] != ele[4][16];
    ele[3][16] != ele[4][17];
    ele[3][16] != ele[4][18];
    ele[3][16] != ele[4][19];
    ele[3][16] != ele[5][16];
    ele[3][16] != ele[6][16];
    ele[3][16] != ele[7][16];
    ele[3][16] != ele[8][16];
    ele[3][16] != ele[9][16];
    ele[3][17] != ele[10][17];
    ele[3][17] != ele[11][17];
    ele[3][17] != ele[12][17];
    ele[3][17] != ele[13][17];
    ele[3][17] != ele[14][17];
    ele[3][17] != ele[15][17];
    ele[3][17] != ele[16][17];
    ele[3][17] != ele[17][17];
    ele[3][17] != ele[18][17];
    ele[3][17] != ele[19][17];
    ele[3][17] != ele[20][17];
    ele[3][17] != ele[21][17];
    ele[3][17] != ele[22][17];
    ele[3][17] != ele[23][17];
    ele[3][17] != ele[24][17];
    ele[3][17] != ele[3][18];
    ele[3][17] != ele[3][19];
    ele[3][17] != ele[3][20];
    ele[3][17] != ele[3][21];
    ele[3][17] != ele[3][22];
    ele[3][17] != ele[3][23];
    ele[3][17] != ele[3][24];
    ele[3][17] != ele[4][15];
    ele[3][17] != ele[4][16];
    ele[3][17] != ele[4][17];
    ele[3][17] != ele[4][18];
    ele[3][17] != ele[4][19];
    ele[3][17] != ele[5][17];
    ele[3][17] != ele[6][17];
    ele[3][17] != ele[7][17];
    ele[3][17] != ele[8][17];
    ele[3][17] != ele[9][17];
    ele[3][18] != ele[10][18];
    ele[3][18] != ele[11][18];
    ele[3][18] != ele[12][18];
    ele[3][18] != ele[13][18];
    ele[3][18] != ele[14][18];
    ele[3][18] != ele[15][18];
    ele[3][18] != ele[16][18];
    ele[3][18] != ele[17][18];
    ele[3][18] != ele[18][18];
    ele[3][18] != ele[19][18];
    ele[3][18] != ele[20][18];
    ele[3][18] != ele[21][18];
    ele[3][18] != ele[22][18];
    ele[3][18] != ele[23][18];
    ele[3][18] != ele[24][18];
    ele[3][18] != ele[3][19];
    ele[3][18] != ele[3][20];
    ele[3][18] != ele[3][21];
    ele[3][18] != ele[3][22];
    ele[3][18] != ele[3][23];
    ele[3][18] != ele[3][24];
    ele[3][18] != ele[4][15];
    ele[3][18] != ele[4][16];
    ele[3][18] != ele[4][17];
    ele[3][18] != ele[4][18];
    ele[3][18] != ele[4][19];
    ele[3][18] != ele[5][18];
    ele[3][18] != ele[6][18];
    ele[3][18] != ele[7][18];
    ele[3][18] != ele[8][18];
    ele[3][18] != ele[9][18];
    ele[3][19] != ele[10][19];
    ele[3][19] != ele[11][19];
    ele[3][19] != ele[12][19];
    ele[3][19] != ele[13][19];
    ele[3][19] != ele[14][19];
    ele[3][19] != ele[15][19];
    ele[3][19] != ele[16][19];
    ele[3][19] != ele[17][19];
    ele[3][19] != ele[18][19];
    ele[3][19] != ele[19][19];
    ele[3][19] != ele[20][19];
    ele[3][19] != ele[21][19];
    ele[3][19] != ele[22][19];
    ele[3][19] != ele[23][19];
    ele[3][19] != ele[24][19];
    ele[3][19] != ele[3][20];
    ele[3][19] != ele[3][21];
    ele[3][19] != ele[3][22];
    ele[3][19] != ele[3][23];
    ele[3][19] != ele[3][24];
    ele[3][19] != ele[4][15];
    ele[3][19] != ele[4][16];
    ele[3][19] != ele[4][17];
    ele[3][19] != ele[4][18];
    ele[3][19] != ele[4][19];
    ele[3][19] != ele[5][19];
    ele[3][19] != ele[6][19];
    ele[3][19] != ele[7][19];
    ele[3][19] != ele[8][19];
    ele[3][19] != ele[9][19];
    ele[3][2] != ele[10][2];
    ele[3][2] != ele[11][2];
    ele[3][2] != ele[12][2];
    ele[3][2] != ele[13][2];
    ele[3][2] != ele[14][2];
    ele[3][2] != ele[15][2];
    ele[3][2] != ele[16][2];
    ele[3][2] != ele[17][2];
    ele[3][2] != ele[18][2];
    ele[3][2] != ele[19][2];
    ele[3][2] != ele[20][2];
    ele[3][2] != ele[21][2];
    ele[3][2] != ele[22][2];
    ele[3][2] != ele[23][2];
    ele[3][2] != ele[24][2];
    ele[3][2] != ele[3][10];
    ele[3][2] != ele[3][11];
    ele[3][2] != ele[3][12];
    ele[3][2] != ele[3][13];
    ele[3][2] != ele[3][14];
    ele[3][2] != ele[3][15];
    ele[3][2] != ele[3][16];
    ele[3][2] != ele[3][17];
    ele[3][2] != ele[3][18];
    ele[3][2] != ele[3][19];
    ele[3][2] != ele[3][20];
    ele[3][2] != ele[3][21];
    ele[3][2] != ele[3][22];
    ele[3][2] != ele[3][23];
    ele[3][2] != ele[3][24];
    ele[3][2] != ele[3][3];
    ele[3][2] != ele[3][4];
    ele[3][2] != ele[3][5];
    ele[3][2] != ele[3][6];
    ele[3][2] != ele[3][7];
    ele[3][2] != ele[3][8];
    ele[3][2] != ele[3][9];
    ele[3][2] != ele[4][0];
    ele[3][2] != ele[4][1];
    ele[3][2] != ele[4][2];
    ele[3][2] != ele[4][3];
    ele[3][2] != ele[4][4];
    ele[3][2] != ele[5][2];
    ele[3][2] != ele[6][2];
    ele[3][2] != ele[7][2];
    ele[3][2] != ele[8][2];
    ele[3][2] != ele[9][2];
    ele[3][20] != ele[10][20];
    ele[3][20] != ele[11][20];
    ele[3][20] != ele[12][20];
    ele[3][20] != ele[13][20];
    ele[3][20] != ele[14][20];
    ele[3][20] != ele[15][20];
    ele[3][20] != ele[16][20];
    ele[3][20] != ele[17][20];
    ele[3][20] != ele[18][20];
    ele[3][20] != ele[19][20];
    ele[3][20] != ele[20][20];
    ele[3][20] != ele[21][20];
    ele[3][20] != ele[22][20];
    ele[3][20] != ele[23][20];
    ele[3][20] != ele[24][20];
    ele[3][20] != ele[3][21];
    ele[3][20] != ele[3][22];
    ele[3][20] != ele[3][23];
    ele[3][20] != ele[3][24];
    ele[3][20] != ele[4][20];
    ele[3][20] != ele[4][21];
    ele[3][20] != ele[4][22];
    ele[3][20] != ele[4][23];
    ele[3][20] != ele[4][24];
    ele[3][20] != ele[5][20];
    ele[3][20] != ele[6][20];
    ele[3][20] != ele[7][20];
    ele[3][20] != ele[8][20];
    ele[3][20] != ele[9][20];
    ele[3][21] != ele[10][21];
    ele[3][21] != ele[11][21];
    ele[3][21] != ele[12][21];
    ele[3][21] != ele[13][21];
    ele[3][21] != ele[14][21];
    ele[3][21] != ele[15][21];
    ele[3][21] != ele[16][21];
    ele[3][21] != ele[17][21];
    ele[3][21] != ele[18][21];
    ele[3][21] != ele[19][21];
    ele[3][21] != ele[20][21];
    ele[3][21] != ele[21][21];
    ele[3][21] != ele[22][21];
    ele[3][21] != ele[23][21];
    ele[3][21] != ele[24][21];
    ele[3][21] != ele[3][22];
    ele[3][21] != ele[3][23];
    ele[3][21] != ele[3][24];
    ele[3][21] != ele[4][20];
    ele[3][21] != ele[4][21];
    ele[3][21] != ele[4][22];
    ele[3][21] != ele[4][23];
    ele[3][21] != ele[4][24];
    ele[3][21] != ele[5][21];
    ele[3][21] != ele[6][21];
    ele[3][21] != ele[7][21];
    ele[3][21] != ele[8][21];
    ele[3][21] != ele[9][21];
    ele[3][22] != ele[10][22];
    ele[3][22] != ele[11][22];
    ele[3][22] != ele[12][22];
    ele[3][22] != ele[13][22];
    ele[3][22] != ele[14][22];
    ele[3][22] != ele[15][22];
    ele[3][22] != ele[16][22];
    ele[3][22] != ele[17][22];
    ele[3][22] != ele[18][22];
    ele[3][22] != ele[19][22];
    ele[3][22] != ele[20][22];
    ele[3][22] != ele[21][22];
    ele[3][22] != ele[22][22];
    ele[3][22] != ele[23][22];
    ele[3][22] != ele[24][22];
    ele[3][22] != ele[3][23];
    ele[3][22] != ele[3][24];
    ele[3][22] != ele[4][20];
    ele[3][22] != ele[4][21];
    ele[3][22] != ele[4][22];
    ele[3][22] != ele[4][23];
    ele[3][22] != ele[4][24];
    ele[3][22] != ele[5][22];
    ele[3][22] != ele[6][22];
    ele[3][22] != ele[7][22];
    ele[3][22] != ele[8][22];
    ele[3][22] != ele[9][22];
    ele[3][23] != ele[10][23];
    ele[3][23] != ele[11][23];
    ele[3][23] != ele[12][23];
    ele[3][23] != ele[13][23];
    ele[3][23] != ele[14][23];
    ele[3][23] != ele[15][23];
    ele[3][23] != ele[16][23];
    ele[3][23] != ele[17][23];
    ele[3][23] != ele[18][23];
    ele[3][23] != ele[19][23];
    ele[3][23] != ele[20][23];
    ele[3][23] != ele[21][23];
    ele[3][23] != ele[22][23];
    ele[3][23] != ele[23][23];
    ele[3][23] != ele[24][23];
    ele[3][23] != ele[3][24];
    ele[3][23] != ele[4][20];
    ele[3][23] != ele[4][21];
    ele[3][23] != ele[4][22];
    ele[3][23] != ele[4][23];
    ele[3][23] != ele[4][24];
    ele[3][23] != ele[5][23];
    ele[3][23] != ele[6][23];
    ele[3][23] != ele[7][23];
    ele[3][23] != ele[8][23];
    ele[3][23] != ele[9][23];
    ele[3][24] != ele[10][24];
    ele[3][24] != ele[11][24];
    ele[3][24] != ele[12][24];
    ele[3][24] != ele[13][24];
    ele[3][24] != ele[14][24];
    ele[3][24] != ele[15][24];
    ele[3][24] != ele[16][24];
    ele[3][24] != ele[17][24];
    ele[3][24] != ele[18][24];
    ele[3][24] != ele[19][24];
    ele[3][24] != ele[20][24];
    ele[3][24] != ele[21][24];
    ele[3][24] != ele[22][24];
    ele[3][24] != ele[23][24];
    ele[3][24] != ele[24][24];
    ele[3][24] != ele[4][20];
    ele[3][24] != ele[4][21];
    ele[3][24] != ele[4][22];
    ele[3][24] != ele[4][23];
    ele[3][24] != ele[4][24];
    ele[3][24] != ele[5][24];
    ele[3][24] != ele[6][24];
    ele[3][24] != ele[7][24];
    ele[3][24] != ele[8][24];
    ele[3][24] != ele[9][24];
    ele[3][3] != ele[10][3];
    ele[3][3] != ele[11][3];
    ele[3][3] != ele[12][3];
    ele[3][3] != ele[13][3];
    ele[3][3] != ele[14][3];
    ele[3][3] != ele[15][3];
    ele[3][3] != ele[16][3];
    ele[3][3] != ele[17][3];
    ele[3][3] != ele[18][3];
    ele[3][3] != ele[19][3];
    ele[3][3] != ele[20][3];
    ele[3][3] != ele[21][3];
    ele[3][3] != ele[22][3];
    ele[3][3] != ele[23][3];
    ele[3][3] != ele[24][3];
    ele[3][3] != ele[3][10];
    ele[3][3] != ele[3][11];
    ele[3][3] != ele[3][12];
    ele[3][3] != ele[3][13];
    ele[3][3] != ele[3][14];
    ele[3][3] != ele[3][15];
    ele[3][3] != ele[3][16];
    ele[3][3] != ele[3][17];
    ele[3][3] != ele[3][18];
    ele[3][3] != ele[3][19];
    ele[3][3] != ele[3][20];
    ele[3][3] != ele[3][21];
    ele[3][3] != ele[3][22];
    ele[3][3] != ele[3][23];
    ele[3][3] != ele[3][24];
    ele[3][3] != ele[3][4];
    ele[3][3] != ele[3][5];
    ele[3][3] != ele[3][6];
    ele[3][3] != ele[3][7];
    ele[3][3] != ele[3][8];
    ele[3][3] != ele[3][9];
    ele[3][3] != ele[4][0];
    ele[3][3] != ele[4][1];
    ele[3][3] != ele[4][2];
    ele[3][3] != ele[4][3];
    ele[3][3] != ele[4][4];
    ele[3][3] != ele[5][3];
    ele[3][3] != ele[6][3];
    ele[3][3] != ele[7][3];
    ele[3][3] != ele[8][3];
    ele[3][3] != ele[9][3];
    ele[3][4] != ele[10][4];
    ele[3][4] != ele[11][4];
    ele[3][4] != ele[12][4];
    ele[3][4] != ele[13][4];
    ele[3][4] != ele[14][4];
    ele[3][4] != ele[15][4];
    ele[3][4] != ele[16][4];
    ele[3][4] != ele[17][4];
    ele[3][4] != ele[18][4];
    ele[3][4] != ele[19][4];
    ele[3][4] != ele[20][4];
    ele[3][4] != ele[21][4];
    ele[3][4] != ele[22][4];
    ele[3][4] != ele[23][4];
    ele[3][4] != ele[24][4];
    ele[3][4] != ele[3][10];
    ele[3][4] != ele[3][11];
    ele[3][4] != ele[3][12];
    ele[3][4] != ele[3][13];
    ele[3][4] != ele[3][14];
    ele[3][4] != ele[3][15];
    ele[3][4] != ele[3][16];
    ele[3][4] != ele[3][17];
    ele[3][4] != ele[3][18];
    ele[3][4] != ele[3][19];
    ele[3][4] != ele[3][20];
    ele[3][4] != ele[3][21];
    ele[3][4] != ele[3][22];
    ele[3][4] != ele[3][23];
    ele[3][4] != ele[3][24];
    ele[3][4] != ele[3][5];
    ele[3][4] != ele[3][6];
    ele[3][4] != ele[3][7];
    ele[3][4] != ele[3][8];
    ele[3][4] != ele[3][9];
    ele[3][4] != ele[4][0];
    ele[3][4] != ele[4][1];
    ele[3][4] != ele[4][2];
    ele[3][4] != ele[4][3];
    ele[3][4] != ele[4][4];
    ele[3][4] != ele[5][4];
    ele[3][4] != ele[6][4];
    ele[3][4] != ele[7][4];
    ele[3][4] != ele[8][4];
    ele[3][4] != ele[9][4];
    ele[3][5] != ele[10][5];
    ele[3][5] != ele[11][5];
    ele[3][5] != ele[12][5];
    ele[3][5] != ele[13][5];
    ele[3][5] != ele[14][5];
    ele[3][5] != ele[15][5];
    ele[3][5] != ele[16][5];
    ele[3][5] != ele[17][5];
    ele[3][5] != ele[18][5];
    ele[3][5] != ele[19][5];
    ele[3][5] != ele[20][5];
    ele[3][5] != ele[21][5];
    ele[3][5] != ele[22][5];
    ele[3][5] != ele[23][5];
    ele[3][5] != ele[24][5];
    ele[3][5] != ele[3][10];
    ele[3][5] != ele[3][11];
    ele[3][5] != ele[3][12];
    ele[3][5] != ele[3][13];
    ele[3][5] != ele[3][14];
    ele[3][5] != ele[3][15];
    ele[3][5] != ele[3][16];
    ele[3][5] != ele[3][17];
    ele[3][5] != ele[3][18];
    ele[3][5] != ele[3][19];
    ele[3][5] != ele[3][20];
    ele[3][5] != ele[3][21];
    ele[3][5] != ele[3][22];
    ele[3][5] != ele[3][23];
    ele[3][5] != ele[3][24];
    ele[3][5] != ele[3][6];
    ele[3][5] != ele[3][7];
    ele[3][5] != ele[3][8];
    ele[3][5] != ele[3][9];
    ele[3][5] != ele[4][5];
    ele[3][5] != ele[4][6];
    ele[3][5] != ele[4][7];
    ele[3][5] != ele[4][8];
    ele[3][5] != ele[4][9];
    ele[3][5] != ele[5][5];
    ele[3][5] != ele[6][5];
    ele[3][5] != ele[7][5];
    ele[3][5] != ele[8][5];
    ele[3][5] != ele[9][5];
    ele[3][6] != ele[10][6];
    ele[3][6] != ele[11][6];
    ele[3][6] != ele[12][6];
    ele[3][6] != ele[13][6];
    ele[3][6] != ele[14][6];
    ele[3][6] != ele[15][6];
    ele[3][6] != ele[16][6];
    ele[3][6] != ele[17][6];
    ele[3][6] != ele[18][6];
    ele[3][6] != ele[19][6];
    ele[3][6] != ele[20][6];
    ele[3][6] != ele[21][6];
    ele[3][6] != ele[22][6];
    ele[3][6] != ele[23][6];
    ele[3][6] != ele[24][6];
    ele[3][6] != ele[3][10];
    ele[3][6] != ele[3][11];
    ele[3][6] != ele[3][12];
    ele[3][6] != ele[3][13];
    ele[3][6] != ele[3][14];
    ele[3][6] != ele[3][15];
    ele[3][6] != ele[3][16];
    ele[3][6] != ele[3][17];
    ele[3][6] != ele[3][18];
    ele[3][6] != ele[3][19];
    ele[3][6] != ele[3][20];
    ele[3][6] != ele[3][21];
    ele[3][6] != ele[3][22];
    ele[3][6] != ele[3][23];
    ele[3][6] != ele[3][24];
    ele[3][6] != ele[3][7];
    ele[3][6] != ele[3][8];
    ele[3][6] != ele[3][9];
    ele[3][6] != ele[4][5];
    ele[3][6] != ele[4][6];
    ele[3][6] != ele[4][7];
    ele[3][6] != ele[4][8];
    ele[3][6] != ele[4][9];
    ele[3][6] != ele[5][6];
    ele[3][6] != ele[6][6];
    ele[3][6] != ele[7][6];
    ele[3][6] != ele[8][6];
    ele[3][6] != ele[9][6];
    ele[3][7] != ele[10][7];
    ele[3][7] != ele[11][7];
    ele[3][7] != ele[12][7];
    ele[3][7] != ele[13][7];
    ele[3][7] != ele[14][7];
    ele[3][7] != ele[15][7];
    ele[3][7] != ele[16][7];
    ele[3][7] != ele[17][7];
    ele[3][7] != ele[18][7];
    ele[3][7] != ele[19][7];
    ele[3][7] != ele[20][7];
    ele[3][7] != ele[21][7];
    ele[3][7] != ele[22][7];
    ele[3][7] != ele[23][7];
    ele[3][7] != ele[24][7];
    ele[3][7] != ele[3][10];
    ele[3][7] != ele[3][11];
    ele[3][7] != ele[3][12];
    ele[3][7] != ele[3][13];
    ele[3][7] != ele[3][14];
    ele[3][7] != ele[3][15];
    ele[3][7] != ele[3][16];
    ele[3][7] != ele[3][17];
    ele[3][7] != ele[3][18];
    ele[3][7] != ele[3][19];
    ele[3][7] != ele[3][20];
    ele[3][7] != ele[3][21];
    ele[3][7] != ele[3][22];
    ele[3][7] != ele[3][23];
    ele[3][7] != ele[3][24];
    ele[3][7] != ele[3][8];
    ele[3][7] != ele[3][9];
    ele[3][7] != ele[4][5];
    ele[3][7] != ele[4][6];
    ele[3][7] != ele[4][7];
    ele[3][7] != ele[4][8];
    ele[3][7] != ele[4][9];
    ele[3][7] != ele[5][7];
    ele[3][7] != ele[6][7];
    ele[3][7] != ele[7][7];
    ele[3][7] != ele[8][7];
    ele[3][7] != ele[9][7];
    ele[3][8] != ele[10][8];
    ele[3][8] != ele[11][8];
    ele[3][8] != ele[12][8];
    ele[3][8] != ele[13][8];
    ele[3][8] != ele[14][8];
    ele[3][8] != ele[15][8];
    ele[3][8] != ele[16][8];
    ele[3][8] != ele[17][8];
    ele[3][8] != ele[18][8];
    ele[3][8] != ele[19][8];
    ele[3][8] != ele[20][8];
    ele[3][8] != ele[21][8];
    ele[3][8] != ele[22][8];
    ele[3][8] != ele[23][8];
    ele[3][8] != ele[24][8];
    ele[3][8] != ele[3][10];
    ele[3][8] != ele[3][11];
    ele[3][8] != ele[3][12];
    ele[3][8] != ele[3][13];
    ele[3][8] != ele[3][14];
    ele[3][8] != ele[3][15];
    ele[3][8] != ele[3][16];
    ele[3][8] != ele[3][17];
    ele[3][8] != ele[3][18];
    ele[3][8] != ele[3][19];
    ele[3][8] != ele[3][20];
    ele[3][8] != ele[3][21];
    ele[3][8] != ele[3][22];
    ele[3][8] != ele[3][23];
    ele[3][8] != ele[3][24];
    ele[3][8] != ele[3][9];
    ele[3][8] != ele[4][5];
    ele[3][8] != ele[4][6];
    ele[3][8] != ele[4][7];
    ele[3][8] != ele[4][8];
    ele[3][8] != ele[4][9];
    ele[3][8] != ele[5][8];
    ele[3][8] != ele[6][8];
    ele[3][8] != ele[7][8];
    ele[3][8] != ele[8][8];
    ele[3][8] != ele[9][8];
    ele[3][9] != ele[10][9];
    ele[3][9] != ele[11][9];
    ele[3][9] != ele[12][9];
    ele[3][9] != ele[13][9];
    ele[3][9] != ele[14][9];
    ele[3][9] != ele[15][9];
    ele[3][9] != ele[16][9];
    ele[3][9] != ele[17][9];
    ele[3][9] != ele[18][9];
    ele[3][9] != ele[19][9];
    ele[3][9] != ele[20][9];
    ele[3][9] != ele[21][9];
    ele[3][9] != ele[22][9];
    ele[3][9] != ele[23][9];
    ele[3][9] != ele[24][9];
    ele[3][9] != ele[3][10];
    ele[3][9] != ele[3][11];
    ele[3][9] != ele[3][12];
    ele[3][9] != ele[3][13];
    ele[3][9] != ele[3][14];
    ele[3][9] != ele[3][15];
    ele[3][9] != ele[3][16];
    ele[3][9] != ele[3][17];
    ele[3][9] != ele[3][18];
    ele[3][9] != ele[3][19];
    ele[3][9] != ele[3][20];
    ele[3][9] != ele[3][21];
    ele[3][9] != ele[3][22];
    ele[3][9] != ele[3][23];
    ele[3][9] != ele[3][24];
    ele[3][9] != ele[4][5];
    ele[3][9] != ele[4][6];
    ele[3][9] != ele[4][7];
    ele[3][9] != ele[4][8];
    ele[3][9] != ele[4][9];
    ele[3][9] != ele[5][9];
    ele[3][9] != ele[6][9];
    ele[3][9] != ele[7][9];
    ele[3][9] != ele[8][9];
    ele[3][9] != ele[9][9];
    ele[4][0] != ele[10][0];
    ele[4][0] != ele[11][0];
    ele[4][0] != ele[12][0];
    ele[4][0] != ele[13][0];
    ele[4][0] != ele[14][0];
    ele[4][0] != ele[15][0];
    ele[4][0] != ele[16][0];
    ele[4][0] != ele[17][0];
    ele[4][0] != ele[18][0];
    ele[4][0] != ele[19][0];
    ele[4][0] != ele[20][0];
    ele[4][0] != ele[21][0];
    ele[4][0] != ele[22][0];
    ele[4][0] != ele[23][0];
    ele[4][0] != ele[24][0];
    ele[4][0] != ele[4][1];
    ele[4][0] != ele[4][10];
    ele[4][0] != ele[4][11];
    ele[4][0] != ele[4][12];
    ele[4][0] != ele[4][13];
    ele[4][0] != ele[4][14];
    ele[4][0] != ele[4][15];
    ele[4][0] != ele[4][16];
    ele[4][0] != ele[4][17];
    ele[4][0] != ele[4][18];
    ele[4][0] != ele[4][19];
    ele[4][0] != ele[4][2];
    ele[4][0] != ele[4][20];
    ele[4][0] != ele[4][21];
    ele[4][0] != ele[4][22];
    ele[4][0] != ele[4][23];
    ele[4][0] != ele[4][24];
    ele[4][0] != ele[4][3];
    ele[4][0] != ele[4][4];
    ele[4][0] != ele[4][5];
    ele[4][0] != ele[4][6];
    ele[4][0] != ele[4][7];
    ele[4][0] != ele[4][8];
    ele[4][0] != ele[4][9];
    ele[4][0] != ele[5][0];
    ele[4][0] != ele[6][0];
    ele[4][0] != ele[7][0];
    ele[4][0] != ele[8][0];
    ele[4][0] != ele[9][0];
    ele[4][1] != ele[10][1];
    ele[4][1] != ele[11][1];
    ele[4][1] != ele[12][1];
    ele[4][1] != ele[13][1];
    ele[4][1] != ele[14][1];
    ele[4][1] != ele[15][1];
    ele[4][1] != ele[16][1];
    ele[4][1] != ele[17][1];
    ele[4][1] != ele[18][1];
    ele[4][1] != ele[19][1];
    ele[4][1] != ele[20][1];
    ele[4][1] != ele[21][1];
    ele[4][1] != ele[22][1];
    ele[4][1] != ele[23][1];
    ele[4][1] != ele[24][1];
    ele[4][1] != ele[4][10];
    ele[4][1] != ele[4][11];
    ele[4][1] != ele[4][12];
    ele[4][1] != ele[4][13];
    ele[4][1] != ele[4][14];
    ele[4][1] != ele[4][15];
    ele[4][1] != ele[4][16];
    ele[4][1] != ele[4][17];
    ele[4][1] != ele[4][18];
    ele[4][1] != ele[4][19];
    ele[4][1] != ele[4][2];
    ele[4][1] != ele[4][20];
    ele[4][1] != ele[4][21];
    ele[4][1] != ele[4][22];
    ele[4][1] != ele[4][23];
    ele[4][1] != ele[4][24];
    ele[4][1] != ele[4][3];
    ele[4][1] != ele[4][4];
    ele[4][1] != ele[4][5];
    ele[4][1] != ele[4][6];
    ele[4][1] != ele[4][7];
    ele[4][1] != ele[4][8];
    ele[4][1] != ele[4][9];
    ele[4][1] != ele[5][1];
    ele[4][1] != ele[6][1];
    ele[4][1] != ele[7][1];
    ele[4][1] != ele[8][1];
    ele[4][1] != ele[9][1];
    ele[4][10] != ele[10][10];
    ele[4][10] != ele[11][10];
    ele[4][10] != ele[12][10];
    ele[4][10] != ele[13][10];
    ele[4][10] != ele[14][10];
    ele[4][10] != ele[15][10];
    ele[4][10] != ele[16][10];
    ele[4][10] != ele[17][10];
    ele[4][10] != ele[18][10];
    ele[4][10] != ele[19][10];
    ele[4][10] != ele[20][10];
    ele[4][10] != ele[21][10];
    ele[4][10] != ele[22][10];
    ele[4][10] != ele[23][10];
    ele[4][10] != ele[24][10];
    ele[4][10] != ele[4][11];
    ele[4][10] != ele[4][12];
    ele[4][10] != ele[4][13];
    ele[4][10] != ele[4][14];
    ele[4][10] != ele[4][15];
    ele[4][10] != ele[4][16];
    ele[4][10] != ele[4][17];
    ele[4][10] != ele[4][18];
    ele[4][10] != ele[4][19];
    ele[4][10] != ele[4][20];
    ele[4][10] != ele[4][21];
    ele[4][10] != ele[4][22];
    ele[4][10] != ele[4][23];
    ele[4][10] != ele[4][24];
    ele[4][10] != ele[5][10];
    ele[4][10] != ele[6][10];
    ele[4][10] != ele[7][10];
    ele[4][10] != ele[8][10];
    ele[4][10] != ele[9][10];
    ele[4][11] != ele[10][11];
    ele[4][11] != ele[11][11];
    ele[4][11] != ele[12][11];
    ele[4][11] != ele[13][11];
    ele[4][11] != ele[14][11];
    ele[4][11] != ele[15][11];
    ele[4][11] != ele[16][11];
    ele[4][11] != ele[17][11];
    ele[4][11] != ele[18][11];
    ele[4][11] != ele[19][11];
    ele[4][11] != ele[20][11];
    ele[4][11] != ele[21][11];
    ele[4][11] != ele[22][11];
    ele[4][11] != ele[23][11];
    ele[4][11] != ele[24][11];
    ele[4][11] != ele[4][12];
    ele[4][11] != ele[4][13];
    ele[4][11] != ele[4][14];
    ele[4][11] != ele[4][15];
    ele[4][11] != ele[4][16];
    ele[4][11] != ele[4][17];
    ele[4][11] != ele[4][18];
    ele[4][11] != ele[4][19];
    ele[4][11] != ele[4][20];
    ele[4][11] != ele[4][21];
    ele[4][11] != ele[4][22];
    ele[4][11] != ele[4][23];
    ele[4][11] != ele[4][24];
    ele[4][11] != ele[5][11];
    ele[4][11] != ele[6][11];
    ele[4][11] != ele[7][11];
    ele[4][11] != ele[8][11];
    ele[4][11] != ele[9][11];
    ele[4][12] != ele[10][12];
    ele[4][12] != ele[11][12];
    ele[4][12] != ele[12][12];
    ele[4][12] != ele[13][12];
    ele[4][12] != ele[14][12];
    ele[4][12] != ele[15][12];
    ele[4][12] != ele[16][12];
    ele[4][12] != ele[17][12];
    ele[4][12] != ele[18][12];
    ele[4][12] != ele[19][12];
    ele[4][12] != ele[20][12];
    ele[4][12] != ele[21][12];
    ele[4][12] != ele[22][12];
    ele[4][12] != ele[23][12];
    ele[4][12] != ele[24][12];
    ele[4][12] != ele[4][13];
    ele[4][12] != ele[4][14];
    ele[4][12] != ele[4][15];
    ele[4][12] != ele[4][16];
    ele[4][12] != ele[4][17];
    ele[4][12] != ele[4][18];
    ele[4][12] != ele[4][19];
    ele[4][12] != ele[4][20];
    ele[4][12] != ele[4][21];
    ele[4][12] != ele[4][22];
    ele[4][12] != ele[4][23];
    ele[4][12] != ele[4][24];
    ele[4][12] != ele[5][12];
    ele[4][12] != ele[6][12];
    ele[4][12] != ele[7][12];
    ele[4][12] != ele[8][12];
    ele[4][12] != ele[9][12];
    ele[4][13] != ele[10][13];
    ele[4][13] != ele[11][13];
    ele[4][13] != ele[12][13];
    ele[4][13] != ele[13][13];
    ele[4][13] != ele[14][13];
    ele[4][13] != ele[15][13];
    ele[4][13] != ele[16][13];
    ele[4][13] != ele[17][13];
    ele[4][13] != ele[18][13];
    ele[4][13] != ele[19][13];
    ele[4][13] != ele[20][13];
    ele[4][13] != ele[21][13];
    ele[4][13] != ele[22][13];
    ele[4][13] != ele[23][13];
    ele[4][13] != ele[24][13];
    ele[4][13] != ele[4][14];
    ele[4][13] != ele[4][15];
    ele[4][13] != ele[4][16];
    ele[4][13] != ele[4][17];
    ele[4][13] != ele[4][18];
    ele[4][13] != ele[4][19];
    ele[4][13] != ele[4][20];
    ele[4][13] != ele[4][21];
    ele[4][13] != ele[4][22];
    ele[4][13] != ele[4][23];
    ele[4][13] != ele[4][24];
    ele[4][13] != ele[5][13];
    ele[4][13] != ele[6][13];
    ele[4][13] != ele[7][13];
    ele[4][13] != ele[8][13];
    ele[4][13] != ele[9][13];
    ele[4][14] != ele[10][14];
    ele[4][14] != ele[11][14];
    ele[4][14] != ele[12][14];
    ele[4][14] != ele[13][14];
    ele[4][14] != ele[14][14];
    ele[4][14] != ele[15][14];
    ele[4][14] != ele[16][14];
    ele[4][14] != ele[17][14];
    ele[4][14] != ele[18][14];
    ele[4][14] != ele[19][14];
    ele[4][14] != ele[20][14];
    ele[4][14] != ele[21][14];
    ele[4][14] != ele[22][14];
    ele[4][14] != ele[23][14];
    ele[4][14] != ele[24][14];
    ele[4][14] != ele[4][15];
    ele[4][14] != ele[4][16];
    ele[4][14] != ele[4][17];
    ele[4][14] != ele[4][18];
    ele[4][14] != ele[4][19];
    ele[4][14] != ele[4][20];
    ele[4][14] != ele[4][21];
    ele[4][14] != ele[4][22];
    ele[4][14] != ele[4][23];
    ele[4][14] != ele[4][24];
    ele[4][14] != ele[5][14];
    ele[4][14] != ele[6][14];
    ele[4][14] != ele[7][14];
    ele[4][14] != ele[8][14];
    ele[4][14] != ele[9][14];
    ele[4][15] != ele[10][15];
    ele[4][15] != ele[11][15];
    ele[4][15] != ele[12][15];
    ele[4][15] != ele[13][15];
    ele[4][15] != ele[14][15];
    ele[4][15] != ele[15][15];
    ele[4][15] != ele[16][15];
    ele[4][15] != ele[17][15];
    ele[4][15] != ele[18][15];
    ele[4][15] != ele[19][15];
    ele[4][15] != ele[20][15];
    ele[4][15] != ele[21][15];
    ele[4][15] != ele[22][15];
    ele[4][15] != ele[23][15];
    ele[4][15] != ele[24][15];
    ele[4][15] != ele[4][16];
    ele[4][15] != ele[4][17];
    ele[4][15] != ele[4][18];
    ele[4][15] != ele[4][19];
    ele[4][15] != ele[4][20];
    ele[4][15] != ele[4][21];
    ele[4][15] != ele[4][22];
    ele[4][15] != ele[4][23];
    ele[4][15] != ele[4][24];
    ele[4][15] != ele[5][15];
    ele[4][15] != ele[6][15];
    ele[4][15] != ele[7][15];
    ele[4][15] != ele[8][15];
    ele[4][15] != ele[9][15];
    ele[4][16] != ele[10][16];
    ele[4][16] != ele[11][16];
    ele[4][16] != ele[12][16];
    ele[4][16] != ele[13][16];
    ele[4][16] != ele[14][16];
    ele[4][16] != ele[15][16];
    ele[4][16] != ele[16][16];
    ele[4][16] != ele[17][16];
    ele[4][16] != ele[18][16];
    ele[4][16] != ele[19][16];
    ele[4][16] != ele[20][16];
    ele[4][16] != ele[21][16];
    ele[4][16] != ele[22][16];
    ele[4][16] != ele[23][16];
    ele[4][16] != ele[24][16];
    ele[4][16] != ele[4][17];
    ele[4][16] != ele[4][18];
    ele[4][16] != ele[4][19];
    ele[4][16] != ele[4][20];
    ele[4][16] != ele[4][21];
    ele[4][16] != ele[4][22];
    ele[4][16] != ele[4][23];
    ele[4][16] != ele[4][24];
    ele[4][16] != ele[5][16];
    ele[4][16] != ele[6][16];
    ele[4][16] != ele[7][16];
    ele[4][16] != ele[8][16];
    ele[4][16] != ele[9][16];
    ele[4][17] != ele[10][17];
    ele[4][17] != ele[11][17];
    ele[4][17] != ele[12][17];
    ele[4][17] != ele[13][17];
    ele[4][17] != ele[14][17];
    ele[4][17] != ele[15][17];
    ele[4][17] != ele[16][17];
    ele[4][17] != ele[17][17];
    ele[4][17] != ele[18][17];
    ele[4][17] != ele[19][17];
    ele[4][17] != ele[20][17];
    ele[4][17] != ele[21][17];
    ele[4][17] != ele[22][17];
    ele[4][17] != ele[23][17];
    ele[4][17] != ele[24][17];
    ele[4][17] != ele[4][18];
    ele[4][17] != ele[4][19];
    ele[4][17] != ele[4][20];
    ele[4][17] != ele[4][21];
    ele[4][17] != ele[4][22];
    ele[4][17] != ele[4][23];
    ele[4][17] != ele[4][24];
    ele[4][17] != ele[5][17];
    ele[4][17] != ele[6][17];
    ele[4][17] != ele[7][17];
    ele[4][17] != ele[8][17];
    ele[4][17] != ele[9][17];
    ele[4][18] != ele[10][18];
    ele[4][18] != ele[11][18];
    ele[4][18] != ele[12][18];
    ele[4][18] != ele[13][18];
    ele[4][18] != ele[14][18];
    ele[4][18] != ele[15][18];
    ele[4][18] != ele[16][18];
    ele[4][18] != ele[17][18];
    ele[4][18] != ele[18][18];
    ele[4][18] != ele[19][18];
    ele[4][18] != ele[20][18];
    ele[4][18] != ele[21][18];
    ele[4][18] != ele[22][18];
    ele[4][18] != ele[23][18];
    ele[4][18] != ele[24][18];
    ele[4][18] != ele[4][19];
    ele[4][18] != ele[4][20];
    ele[4][18] != ele[4][21];
    ele[4][18] != ele[4][22];
    ele[4][18] != ele[4][23];
    ele[4][18] != ele[4][24];
    ele[4][18] != ele[5][18];
    ele[4][18] != ele[6][18];
    ele[4][18] != ele[7][18];
    ele[4][18] != ele[8][18];
    ele[4][18] != ele[9][18];
    ele[4][19] != ele[10][19];
    ele[4][19] != ele[11][19];
    ele[4][19] != ele[12][19];
    ele[4][19] != ele[13][19];
    ele[4][19] != ele[14][19];
    ele[4][19] != ele[15][19];
    ele[4][19] != ele[16][19];
    ele[4][19] != ele[17][19];
    ele[4][19] != ele[18][19];
    ele[4][19] != ele[19][19];
    ele[4][19] != ele[20][19];
    ele[4][19] != ele[21][19];
    ele[4][19] != ele[22][19];
    ele[4][19] != ele[23][19];
    ele[4][19] != ele[24][19];
    ele[4][19] != ele[4][20];
    ele[4][19] != ele[4][21];
    ele[4][19] != ele[4][22];
    ele[4][19] != ele[4][23];
    ele[4][19] != ele[4][24];
    ele[4][19] != ele[5][19];
    ele[4][19] != ele[6][19];
    ele[4][19] != ele[7][19];
    ele[4][19] != ele[8][19];
    ele[4][19] != ele[9][19];
    ele[4][2] != ele[10][2];
    ele[4][2] != ele[11][2];
    ele[4][2] != ele[12][2];
    ele[4][2] != ele[13][2];
    ele[4][2] != ele[14][2];
    ele[4][2] != ele[15][2];
    ele[4][2] != ele[16][2];
    ele[4][2] != ele[17][2];
    ele[4][2] != ele[18][2];
    ele[4][2] != ele[19][2];
    ele[4][2] != ele[20][2];
    ele[4][2] != ele[21][2];
    ele[4][2] != ele[22][2];
    ele[4][2] != ele[23][2];
    ele[4][2] != ele[24][2];
    ele[4][2] != ele[4][10];
    ele[4][2] != ele[4][11];
    ele[4][2] != ele[4][12];
    ele[4][2] != ele[4][13];
    ele[4][2] != ele[4][14];
    ele[4][2] != ele[4][15];
    ele[4][2] != ele[4][16];
    ele[4][2] != ele[4][17];
    ele[4][2] != ele[4][18];
    ele[4][2] != ele[4][19];
    ele[4][2] != ele[4][20];
    ele[4][2] != ele[4][21];
    ele[4][2] != ele[4][22];
    ele[4][2] != ele[4][23];
    ele[4][2] != ele[4][24];
    ele[4][2] != ele[4][3];
    ele[4][2] != ele[4][4];
    ele[4][2] != ele[4][5];
    ele[4][2] != ele[4][6];
    ele[4][2] != ele[4][7];
    ele[4][2] != ele[4][8];
    ele[4][2] != ele[4][9];
    ele[4][2] != ele[5][2];
    ele[4][2] != ele[6][2];
    ele[4][2] != ele[7][2];
    ele[4][2] != ele[8][2];
    ele[4][2] != ele[9][2];
    ele[4][20] != ele[10][20];
    ele[4][20] != ele[11][20];
    ele[4][20] != ele[12][20];
    ele[4][20] != ele[13][20];
    ele[4][20] != ele[14][20];
    ele[4][20] != ele[15][20];
    ele[4][20] != ele[16][20];
    ele[4][20] != ele[17][20];
    ele[4][20] != ele[18][20];
    ele[4][20] != ele[19][20];
    ele[4][20] != ele[20][20];
    ele[4][20] != ele[21][20];
    ele[4][20] != ele[22][20];
    ele[4][20] != ele[23][20];
    ele[4][20] != ele[24][20];
    ele[4][20] != ele[4][21];
    ele[4][20] != ele[4][22];
    ele[4][20] != ele[4][23];
    ele[4][20] != ele[4][24];
    ele[4][20] != ele[5][20];
    ele[4][20] != ele[6][20];
    ele[4][20] != ele[7][20];
    ele[4][20] != ele[8][20];
    ele[4][20] != ele[9][20];
    ele[4][21] != ele[10][21];
    ele[4][21] != ele[11][21];
    ele[4][21] != ele[12][21];
    ele[4][21] != ele[13][21];
    ele[4][21] != ele[14][21];
    ele[4][21] != ele[15][21];
    ele[4][21] != ele[16][21];
    ele[4][21] != ele[17][21];
    ele[4][21] != ele[18][21];
    ele[4][21] != ele[19][21];
    ele[4][21] != ele[20][21];
    ele[4][21] != ele[21][21];
    ele[4][21] != ele[22][21];
    ele[4][21] != ele[23][21];
    ele[4][21] != ele[24][21];
    ele[4][21] != ele[4][22];
    ele[4][21] != ele[4][23];
    ele[4][21] != ele[4][24];
    ele[4][21] != ele[5][21];
    ele[4][21] != ele[6][21];
    ele[4][21] != ele[7][21];
    ele[4][21] != ele[8][21];
    ele[4][21] != ele[9][21];
    ele[4][22] != ele[10][22];
    ele[4][22] != ele[11][22];
    ele[4][22] != ele[12][22];
    ele[4][22] != ele[13][22];
    ele[4][22] != ele[14][22];
    ele[4][22] != ele[15][22];
    ele[4][22] != ele[16][22];
    ele[4][22] != ele[17][22];
    ele[4][22] != ele[18][22];
    ele[4][22] != ele[19][22];
    ele[4][22] != ele[20][22];
    ele[4][22] != ele[21][22];
    ele[4][22] != ele[22][22];
    ele[4][22] != ele[23][22];
    ele[4][22] != ele[24][22];
    ele[4][22] != ele[4][23];
    ele[4][22] != ele[4][24];
    ele[4][22] != ele[5][22];
    ele[4][22] != ele[6][22];
    ele[4][22] != ele[7][22];
    ele[4][22] != ele[8][22];
    ele[4][22] != ele[9][22];
    ele[4][23] != ele[10][23];
    ele[4][23] != ele[11][23];
    ele[4][23] != ele[12][23];
    ele[4][23] != ele[13][23];
    ele[4][23] != ele[14][23];
    ele[4][23] != ele[15][23];
    ele[4][23] != ele[16][23];
    ele[4][23] != ele[17][23];
    ele[4][23] != ele[18][23];
    ele[4][23] != ele[19][23];
    ele[4][23] != ele[20][23];
    ele[4][23] != ele[21][23];
    ele[4][23] != ele[22][23];
    ele[4][23] != ele[23][23];
    ele[4][23] != ele[24][23];
    ele[4][23] != ele[4][24];
    ele[4][23] != ele[5][23];
    ele[4][23] != ele[6][23];
    ele[4][23] != ele[7][23];
    ele[4][23] != ele[8][23];
    ele[4][23] != ele[9][23];
    ele[4][24] != ele[10][24];
    ele[4][24] != ele[11][24];
    ele[4][24] != ele[12][24];
    ele[4][24] != ele[13][24];
    ele[4][24] != ele[14][24];
    ele[4][24] != ele[15][24];
    ele[4][24] != ele[16][24];
    ele[4][24] != ele[17][24];
    ele[4][24] != ele[18][24];
    ele[4][24] != ele[19][24];
    ele[4][24] != ele[20][24];
    ele[4][24] != ele[21][24];
    ele[4][24] != ele[22][24];
    ele[4][24] != ele[23][24];
    ele[4][24] != ele[24][24];
    ele[4][24] != ele[5][24];
    ele[4][24] != ele[6][24];
    ele[4][24] != ele[7][24];
    ele[4][24] != ele[8][24];
    ele[4][24] != ele[9][24];
    ele[4][3] != ele[10][3];
    ele[4][3] != ele[11][3];
    ele[4][3] != ele[12][3];
    ele[4][3] != ele[13][3];
    ele[4][3] != ele[14][3];
    ele[4][3] != ele[15][3];
    ele[4][3] != ele[16][3];
    ele[4][3] != ele[17][3];
    ele[4][3] != ele[18][3];
    ele[4][3] != ele[19][3];
    ele[4][3] != ele[20][3];
    ele[4][3] != ele[21][3];
    ele[4][3] != ele[22][3];
    ele[4][3] != ele[23][3];
    ele[4][3] != ele[24][3];
    ele[4][3] != ele[4][10];
    ele[4][3] != ele[4][11];
    ele[4][3] != ele[4][12];
    ele[4][3] != ele[4][13];
    ele[4][3] != ele[4][14];
    ele[4][3] != ele[4][15];
    ele[4][3] != ele[4][16];
    ele[4][3] != ele[4][17];
    ele[4][3] != ele[4][18];
    ele[4][3] != ele[4][19];
    ele[4][3] != ele[4][20];
    ele[4][3] != ele[4][21];
    ele[4][3] != ele[4][22];
    ele[4][3] != ele[4][23];
    ele[4][3] != ele[4][24];
    ele[4][3] != ele[4][4];
    ele[4][3] != ele[4][5];
    ele[4][3] != ele[4][6];
    ele[4][3] != ele[4][7];
    ele[4][3] != ele[4][8];
    ele[4][3] != ele[4][9];
    ele[4][3] != ele[5][3];
    ele[4][3] != ele[6][3];
    ele[4][3] != ele[7][3];
    ele[4][3] != ele[8][3];
    ele[4][3] != ele[9][3];
    ele[4][4] != ele[10][4];
    ele[4][4] != ele[11][4];
    ele[4][4] != ele[12][4];
    ele[4][4] != ele[13][4];
    ele[4][4] != ele[14][4];
    ele[4][4] != ele[15][4];
    ele[4][4] != ele[16][4];
    ele[4][4] != ele[17][4];
    ele[4][4] != ele[18][4];
    ele[4][4] != ele[19][4];
    ele[4][4] != ele[20][4];
    ele[4][4] != ele[21][4];
    ele[4][4] != ele[22][4];
    ele[4][4] != ele[23][4];
    ele[4][4] != ele[24][4];
    ele[4][4] != ele[4][10];
    ele[4][4] != ele[4][11];
    ele[4][4] != ele[4][12];
    ele[4][4] != ele[4][13];
    ele[4][4] != ele[4][14];
    ele[4][4] != ele[4][15];
    ele[4][4] != ele[4][16];
    ele[4][4] != ele[4][17];
    ele[4][4] != ele[4][18];
    ele[4][4] != ele[4][19];
    ele[4][4] != ele[4][20];
    ele[4][4] != ele[4][21];
    ele[4][4] != ele[4][22];
    ele[4][4] != ele[4][23];
    ele[4][4] != ele[4][24];
    ele[4][4] != ele[4][5];
    ele[4][4] != ele[4][6];
    ele[4][4] != ele[4][7];
    ele[4][4] != ele[4][8];
    ele[4][4] != ele[4][9];
    ele[4][4] != ele[5][4];
    ele[4][4] != ele[6][4];
    ele[4][4] != ele[7][4];
    ele[4][4] != ele[8][4];
    ele[4][4] != ele[9][4];
    ele[4][5] != ele[10][5];
    ele[4][5] != ele[11][5];
    ele[4][5] != ele[12][5];
    ele[4][5] != ele[13][5];
    ele[4][5] != ele[14][5];
    ele[4][5] != ele[15][5];
    ele[4][5] != ele[16][5];
    ele[4][5] != ele[17][5];
    ele[4][5] != ele[18][5];
    ele[4][5] != ele[19][5];
    ele[4][5] != ele[20][5];
    ele[4][5] != ele[21][5];
    ele[4][5] != ele[22][5];
    ele[4][5] != ele[23][5];
    ele[4][5] != ele[24][5];
    ele[4][5] != ele[4][10];
    ele[4][5] != ele[4][11];
    ele[4][5] != ele[4][12];
    ele[4][5] != ele[4][13];
    ele[4][5] != ele[4][14];
    ele[4][5] != ele[4][15];
    ele[4][5] != ele[4][16];
    ele[4][5] != ele[4][17];
    ele[4][5] != ele[4][18];
    ele[4][5] != ele[4][19];
    ele[4][5] != ele[4][20];
    ele[4][5] != ele[4][21];
    ele[4][5] != ele[4][22];
    ele[4][5] != ele[4][23];
    ele[4][5] != ele[4][24];
    ele[4][5] != ele[4][6];
    ele[4][5] != ele[4][7];
    ele[4][5] != ele[4][8];
    ele[4][5] != ele[4][9];
    ele[4][5] != ele[5][5];
    ele[4][5] != ele[6][5];
    ele[4][5] != ele[7][5];
    ele[4][5] != ele[8][5];
    ele[4][5] != ele[9][5];
    ele[4][6] != ele[10][6];
    ele[4][6] != ele[11][6];
    ele[4][6] != ele[12][6];
    ele[4][6] != ele[13][6];
    ele[4][6] != ele[14][6];
    ele[4][6] != ele[15][6];
    ele[4][6] != ele[16][6];
    ele[4][6] != ele[17][6];
    ele[4][6] != ele[18][6];
    ele[4][6] != ele[19][6];
    ele[4][6] != ele[20][6];
    ele[4][6] != ele[21][6];
    ele[4][6] != ele[22][6];
    ele[4][6] != ele[23][6];
    ele[4][6] != ele[24][6];
    ele[4][6] != ele[4][10];
    ele[4][6] != ele[4][11];
    ele[4][6] != ele[4][12];
    ele[4][6] != ele[4][13];
    ele[4][6] != ele[4][14];
    ele[4][6] != ele[4][15];
    ele[4][6] != ele[4][16];
    ele[4][6] != ele[4][17];
    ele[4][6] != ele[4][18];
    ele[4][6] != ele[4][19];
    ele[4][6] != ele[4][20];
    ele[4][6] != ele[4][21];
    ele[4][6] != ele[4][22];
    ele[4][6] != ele[4][23];
    ele[4][6] != ele[4][24];
    ele[4][6] != ele[4][7];
    ele[4][6] != ele[4][8];
    ele[4][6] != ele[4][9];
    ele[4][6] != ele[5][6];
    ele[4][6] != ele[6][6];
    ele[4][6] != ele[7][6];
    ele[4][6] != ele[8][6];
    ele[4][6] != ele[9][6];
    ele[4][7] != ele[10][7];
    ele[4][7] != ele[11][7];
    ele[4][7] != ele[12][7];
    ele[4][7] != ele[13][7];
    ele[4][7] != ele[14][7];
    ele[4][7] != ele[15][7];
    ele[4][7] != ele[16][7];
    ele[4][7] != ele[17][7];
    ele[4][7] != ele[18][7];
    ele[4][7] != ele[19][7];
    ele[4][7] != ele[20][7];
    ele[4][7] != ele[21][7];
    ele[4][7] != ele[22][7];
    ele[4][7] != ele[23][7];
    ele[4][7] != ele[24][7];
    ele[4][7] != ele[4][10];
    ele[4][7] != ele[4][11];
    ele[4][7] != ele[4][12];
    ele[4][7] != ele[4][13];
    ele[4][7] != ele[4][14];
    ele[4][7] != ele[4][15];
    ele[4][7] != ele[4][16];
    ele[4][7] != ele[4][17];
    ele[4][7] != ele[4][18];
    ele[4][7] != ele[4][19];
    ele[4][7] != ele[4][20];
    ele[4][7] != ele[4][21];
    ele[4][7] != ele[4][22];
    ele[4][7] != ele[4][23];
    ele[4][7] != ele[4][24];
    ele[4][7] != ele[4][8];
    ele[4][7] != ele[4][9];
    ele[4][7] != ele[5][7];
    ele[4][7] != ele[6][7];
    ele[4][7] != ele[7][7];
    ele[4][7] != ele[8][7];
    ele[4][7] != ele[9][7];
    ele[4][8] != ele[10][8];
    ele[4][8] != ele[11][8];
    ele[4][8] != ele[12][8];
    ele[4][8] != ele[13][8];
    ele[4][8] != ele[14][8];
    ele[4][8] != ele[15][8];
    ele[4][8] != ele[16][8];
    ele[4][8] != ele[17][8];
    ele[4][8] != ele[18][8];
    ele[4][8] != ele[19][8];
    ele[4][8] != ele[20][8];
    ele[4][8] != ele[21][8];
    ele[4][8] != ele[22][8];
    ele[4][8] != ele[23][8];
    ele[4][8] != ele[24][8];
    ele[4][8] != ele[4][10];
    ele[4][8] != ele[4][11];
    ele[4][8] != ele[4][12];
    ele[4][8] != ele[4][13];
    ele[4][8] != ele[4][14];
    ele[4][8] != ele[4][15];
    ele[4][8] != ele[4][16];
    ele[4][8] != ele[4][17];
    ele[4][8] != ele[4][18];
    ele[4][8] != ele[4][19];
    ele[4][8] != ele[4][20];
    ele[4][8] != ele[4][21];
    ele[4][8] != ele[4][22];
    ele[4][8] != ele[4][23];
    ele[4][8] != ele[4][24];
    ele[4][8] != ele[4][9];
    ele[4][8] != ele[5][8];
    ele[4][8] != ele[6][8];
    ele[4][8] != ele[7][8];
    ele[4][8] != ele[8][8];
    ele[4][8] != ele[9][8];
    ele[4][9] != ele[10][9];
    ele[4][9] != ele[11][9];
    ele[4][9] != ele[12][9];
    ele[4][9] != ele[13][9];
    ele[4][9] != ele[14][9];
    ele[4][9] != ele[15][9];
    ele[4][9] != ele[16][9];
    ele[4][9] != ele[17][9];
    ele[4][9] != ele[18][9];
    ele[4][9] != ele[19][9];
    ele[4][9] != ele[20][9];
    ele[4][9] != ele[21][9];
    ele[4][9] != ele[22][9];
    ele[4][9] != ele[23][9];
    ele[4][9] != ele[24][9];
    ele[4][9] != ele[4][10];
    ele[4][9] != ele[4][11];
    ele[4][9] != ele[4][12];
    ele[4][9] != ele[4][13];
    ele[4][9] != ele[4][14];
    ele[4][9] != ele[4][15];
    ele[4][9] != ele[4][16];
    ele[4][9] != ele[4][17];
    ele[4][9] != ele[4][18];
    ele[4][9] != ele[4][19];
    ele[4][9] != ele[4][20];
    ele[4][9] != ele[4][21];
    ele[4][9] != ele[4][22];
    ele[4][9] != ele[4][23];
    ele[4][9] != ele[4][24];
    ele[4][9] != ele[5][9];
    ele[4][9] != ele[6][9];
    ele[4][9] != ele[7][9];
    ele[4][9] != ele[8][9];
    ele[4][9] != ele[9][9];
    ele[5][0] != ele[10][0];
    ele[5][0] != ele[11][0];
    ele[5][0] != ele[12][0];
    ele[5][0] != ele[13][0];
    ele[5][0] != ele[14][0];
    ele[5][0] != ele[15][0];
    ele[5][0] != ele[16][0];
    ele[5][0] != ele[17][0];
    ele[5][0] != ele[18][0];
    ele[5][0] != ele[19][0];
    ele[5][0] != ele[20][0];
    ele[5][0] != ele[21][0];
    ele[5][0] != ele[22][0];
    ele[5][0] != ele[23][0];
    ele[5][0] != ele[24][0];
    ele[5][0] != ele[5][1];
    ele[5][0] != ele[5][10];
    ele[5][0] != ele[5][11];
    ele[5][0] != ele[5][12];
    ele[5][0] != ele[5][13];
    ele[5][0] != ele[5][14];
    ele[5][0] != ele[5][15];
    ele[5][0] != ele[5][16];
    ele[5][0] != ele[5][17];
    ele[5][0] != ele[5][18];
    ele[5][0] != ele[5][19];
    ele[5][0] != ele[5][2];
    ele[5][0] != ele[5][20];
    ele[5][0] != ele[5][21];
    ele[5][0] != ele[5][22];
    ele[5][0] != ele[5][23];
    ele[5][0] != ele[5][24];
    ele[5][0] != ele[5][3];
    ele[5][0] != ele[5][4];
    ele[5][0] != ele[5][5];
    ele[5][0] != ele[5][6];
    ele[5][0] != ele[5][7];
    ele[5][0] != ele[5][8];
    ele[5][0] != ele[5][9];
    ele[5][0] != ele[6][0];
    ele[5][0] != ele[6][1];
    ele[5][0] != ele[6][2];
    ele[5][0] != ele[6][3];
    ele[5][0] != ele[6][4];
    ele[5][0] != ele[7][0];
    ele[5][0] != ele[7][1];
    ele[5][0] != ele[7][2];
    ele[5][0] != ele[7][3];
    ele[5][0] != ele[7][4];
    ele[5][0] != ele[8][0];
    ele[5][0] != ele[8][1];
    ele[5][0] != ele[8][2];
    ele[5][0] != ele[8][3];
    ele[5][0] != ele[8][4];
    ele[5][0] != ele[9][0];
    ele[5][0] != ele[9][1];
    ele[5][0] != ele[9][2];
    ele[5][0] != ele[9][3];
    ele[5][0] != ele[9][4];
    ele[5][1] != ele[10][1];
    ele[5][1] != ele[11][1];
    ele[5][1] != ele[12][1];
    ele[5][1] != ele[13][1];
    ele[5][1] != ele[14][1];
    ele[5][1] != ele[15][1];
    ele[5][1] != ele[16][1];
    ele[5][1] != ele[17][1];
    ele[5][1] != ele[18][1];
    ele[5][1] != ele[19][1];
    ele[5][1] != ele[20][1];
    ele[5][1] != ele[21][1];
    ele[5][1] != ele[22][1];
    ele[5][1] != ele[23][1];
    ele[5][1] != ele[24][1];
    ele[5][1] != ele[5][10];
    ele[5][1] != ele[5][11];
    ele[5][1] != ele[5][12];
    ele[5][1] != ele[5][13];
    ele[5][1] != ele[5][14];
    ele[5][1] != ele[5][15];
    ele[5][1] != ele[5][16];
    ele[5][1] != ele[5][17];
    ele[5][1] != ele[5][18];
    ele[5][1] != ele[5][19];
    ele[5][1] != ele[5][2];
    ele[5][1] != ele[5][20];
    ele[5][1] != ele[5][21];
    ele[5][1] != ele[5][22];
    ele[5][1] != ele[5][23];
    ele[5][1] != ele[5][24];
    ele[5][1] != ele[5][3];
    ele[5][1] != ele[5][4];
    ele[5][1] != ele[5][5];
    ele[5][1] != ele[5][6];
    ele[5][1] != ele[5][7];
    ele[5][1] != ele[5][8];
    ele[5][1] != ele[5][9];
    ele[5][1] != ele[6][0];
    ele[5][1] != ele[6][1];
    ele[5][1] != ele[6][2];
    ele[5][1] != ele[6][3];
    ele[5][1] != ele[6][4];
    ele[5][1] != ele[7][0];
    ele[5][1] != ele[7][1];
    ele[5][1] != ele[7][2];
    ele[5][1] != ele[7][3];
    ele[5][1] != ele[7][4];
    ele[5][1] != ele[8][0];
    ele[5][1] != ele[8][1];
    ele[5][1] != ele[8][2];
    ele[5][1] != ele[8][3];
    ele[5][1] != ele[8][4];
    ele[5][1] != ele[9][0];
    ele[5][1] != ele[9][1];
    ele[5][1] != ele[9][2];
    ele[5][1] != ele[9][3];
    ele[5][1] != ele[9][4];
    ele[5][10] != ele[10][10];
    ele[5][10] != ele[11][10];
    ele[5][10] != ele[12][10];
    ele[5][10] != ele[13][10];
    ele[5][10] != ele[14][10];
    ele[5][10] != ele[15][10];
    ele[5][10] != ele[16][10];
    ele[5][10] != ele[17][10];
    ele[5][10] != ele[18][10];
    ele[5][10] != ele[19][10];
    ele[5][10] != ele[20][10];
    ele[5][10] != ele[21][10];
    ele[5][10] != ele[22][10];
    ele[5][10] != ele[23][10];
    ele[5][10] != ele[24][10];
    ele[5][10] != ele[5][11];
    ele[5][10] != ele[5][12];
    ele[5][10] != ele[5][13];
    ele[5][10] != ele[5][14];
    ele[5][10] != ele[5][15];
    ele[5][10] != ele[5][16];
    ele[5][10] != ele[5][17];
    ele[5][10] != ele[5][18];
    ele[5][10] != ele[5][19];
    ele[5][10] != ele[5][20];
    ele[5][10] != ele[5][21];
    ele[5][10] != ele[5][22];
    ele[5][10] != ele[5][23];
    ele[5][10] != ele[5][24];
    ele[5][10] != ele[6][10];
    ele[5][10] != ele[6][11];
    ele[5][10] != ele[6][12];
    ele[5][10] != ele[6][13];
    ele[5][10] != ele[6][14];
    ele[5][10] != ele[7][10];
    ele[5][10] != ele[7][11];
    ele[5][10] != ele[7][12];
    ele[5][10] != ele[7][13];
    ele[5][10] != ele[7][14];
    ele[5][10] != ele[8][10];
    ele[5][10] != ele[8][11];
    ele[5][10] != ele[8][12];
    ele[5][10] != ele[8][13];
    ele[5][10] != ele[8][14];
    ele[5][10] != ele[9][10];
    ele[5][10] != ele[9][11];
    ele[5][10] != ele[9][12];
    ele[5][10] != ele[9][13];
    ele[5][10] != ele[9][14];
    ele[5][11] != ele[10][11];
    ele[5][11] != ele[11][11];
    ele[5][11] != ele[12][11];
    ele[5][11] != ele[13][11];
    ele[5][11] != ele[14][11];
    ele[5][11] != ele[15][11];
    ele[5][11] != ele[16][11];
    ele[5][11] != ele[17][11];
    ele[5][11] != ele[18][11];
    ele[5][11] != ele[19][11];
    ele[5][11] != ele[20][11];
    ele[5][11] != ele[21][11];
    ele[5][11] != ele[22][11];
    ele[5][11] != ele[23][11];
    ele[5][11] != ele[24][11];
    ele[5][11] != ele[5][12];
    ele[5][11] != ele[5][13];
    ele[5][11] != ele[5][14];
    ele[5][11] != ele[5][15];
    ele[5][11] != ele[5][16];
    ele[5][11] != ele[5][17];
    ele[5][11] != ele[5][18];
    ele[5][11] != ele[5][19];
    ele[5][11] != ele[5][20];
    ele[5][11] != ele[5][21];
    ele[5][11] != ele[5][22];
    ele[5][11] != ele[5][23];
    ele[5][11] != ele[5][24];
    ele[5][11] != ele[6][10];
    ele[5][11] != ele[6][11];
    ele[5][11] != ele[6][12];
    ele[5][11] != ele[6][13];
    ele[5][11] != ele[6][14];
    ele[5][11] != ele[7][10];
    ele[5][11] != ele[7][11];
    ele[5][11] != ele[7][12];
    ele[5][11] != ele[7][13];
    ele[5][11] != ele[7][14];
    ele[5][11] != ele[8][10];
    ele[5][11] != ele[8][11];
    ele[5][11] != ele[8][12];
    ele[5][11] != ele[8][13];
    ele[5][11] != ele[8][14];
    ele[5][11] != ele[9][10];
    ele[5][11] != ele[9][11];
    ele[5][11] != ele[9][12];
    ele[5][11] != ele[9][13];
    ele[5][11] != ele[9][14];
    ele[5][12] != ele[10][12];
    ele[5][12] != ele[11][12];
    ele[5][12] != ele[12][12];
    ele[5][12] != ele[13][12];
    ele[5][12] != ele[14][12];
    ele[5][12] != ele[15][12];
    ele[5][12] != ele[16][12];
    ele[5][12] != ele[17][12];
    ele[5][12] != ele[18][12];
    ele[5][12] != ele[19][12];
    ele[5][12] != ele[20][12];
    ele[5][12] != ele[21][12];
    ele[5][12] != ele[22][12];
    ele[5][12] != ele[23][12];
    ele[5][12] != ele[24][12];
    ele[5][12] != ele[5][13];
    ele[5][12] != ele[5][14];
    ele[5][12] != ele[5][15];
    ele[5][12] != ele[5][16];
    ele[5][12] != ele[5][17];
    ele[5][12] != ele[5][18];
    ele[5][12] != ele[5][19];
    ele[5][12] != ele[5][20];
    ele[5][12] != ele[5][21];
    ele[5][12] != ele[5][22];
    ele[5][12] != ele[5][23];
    ele[5][12] != ele[5][24];
    ele[5][12] != ele[6][10];
    ele[5][12] != ele[6][11];
    ele[5][12] != ele[6][12];
    ele[5][12] != ele[6][13];
    ele[5][12] != ele[6][14];
    ele[5][12] != ele[7][10];
    ele[5][12] != ele[7][11];
    ele[5][12] != ele[7][12];
    ele[5][12] != ele[7][13];
    ele[5][12] != ele[7][14];
    ele[5][12] != ele[8][10];
    ele[5][12] != ele[8][11];
    ele[5][12] != ele[8][12];
    ele[5][12] != ele[8][13];
    ele[5][12] != ele[8][14];
    ele[5][12] != ele[9][10];
    ele[5][12] != ele[9][11];
    ele[5][12] != ele[9][12];
    ele[5][12] != ele[9][13];
    ele[5][12] != ele[9][14];
    ele[5][13] != ele[10][13];
    ele[5][13] != ele[11][13];
    ele[5][13] != ele[12][13];
    ele[5][13] != ele[13][13];
    ele[5][13] != ele[14][13];
    ele[5][13] != ele[15][13];
    ele[5][13] != ele[16][13];
    ele[5][13] != ele[17][13];
    ele[5][13] != ele[18][13];
    ele[5][13] != ele[19][13];
    ele[5][13] != ele[20][13];
    ele[5][13] != ele[21][13];
    ele[5][13] != ele[22][13];
    ele[5][13] != ele[23][13];
    ele[5][13] != ele[24][13];
    ele[5][13] != ele[5][14];
    ele[5][13] != ele[5][15];
    ele[5][13] != ele[5][16];
    ele[5][13] != ele[5][17];
    ele[5][13] != ele[5][18];
    ele[5][13] != ele[5][19];
    ele[5][13] != ele[5][20];
    ele[5][13] != ele[5][21];
    ele[5][13] != ele[5][22];
    ele[5][13] != ele[5][23];
    ele[5][13] != ele[5][24];
    ele[5][13] != ele[6][10];
    ele[5][13] != ele[6][11];
    ele[5][13] != ele[6][12];
    ele[5][13] != ele[6][13];
    ele[5][13] != ele[6][14];
    ele[5][13] != ele[7][10];
    ele[5][13] != ele[7][11];
    ele[5][13] != ele[7][12];
    ele[5][13] != ele[7][13];
    ele[5][13] != ele[7][14];
    ele[5][13] != ele[8][10];
    ele[5][13] != ele[8][11];
    ele[5][13] != ele[8][12];
    ele[5][13] != ele[8][13];
    ele[5][13] != ele[8][14];
    ele[5][13] != ele[9][10];
    ele[5][13] != ele[9][11];
    ele[5][13] != ele[9][12];
    ele[5][13] != ele[9][13];
    ele[5][13] != ele[9][14];
    ele[5][14] != ele[10][14];
    ele[5][14] != ele[11][14];
    ele[5][14] != ele[12][14];
    ele[5][14] != ele[13][14];
    ele[5][14] != ele[14][14];
    ele[5][14] != ele[15][14];
    ele[5][14] != ele[16][14];
    ele[5][14] != ele[17][14];
    ele[5][14] != ele[18][14];
    ele[5][14] != ele[19][14];
    ele[5][14] != ele[20][14];
    ele[5][14] != ele[21][14];
    ele[5][14] != ele[22][14];
    ele[5][14] != ele[23][14];
    ele[5][14] != ele[24][14];
    ele[5][14] != ele[5][15];
    ele[5][14] != ele[5][16];
    ele[5][14] != ele[5][17];
    ele[5][14] != ele[5][18];
    ele[5][14] != ele[5][19];
    ele[5][14] != ele[5][20];
    ele[5][14] != ele[5][21];
    ele[5][14] != ele[5][22];
    ele[5][14] != ele[5][23];
    ele[5][14] != ele[5][24];
    ele[5][14] != ele[6][10];
    ele[5][14] != ele[6][11];
    ele[5][14] != ele[6][12];
    ele[5][14] != ele[6][13];
    ele[5][14] != ele[6][14];
    ele[5][14] != ele[7][10];
    ele[5][14] != ele[7][11];
    ele[5][14] != ele[7][12];
    ele[5][14] != ele[7][13];
    ele[5][14] != ele[7][14];
    ele[5][14] != ele[8][10];
    ele[5][14] != ele[8][11];
    ele[5][14] != ele[8][12];
    ele[5][14] != ele[8][13];
    ele[5][14] != ele[8][14];
    ele[5][14] != ele[9][10];
    ele[5][14] != ele[9][11];
    ele[5][14] != ele[9][12];
    ele[5][14] != ele[9][13];
    ele[5][14] != ele[9][14];
    ele[5][15] != ele[10][15];
    ele[5][15] != ele[11][15];
    ele[5][15] != ele[12][15];
    ele[5][15] != ele[13][15];
    ele[5][15] != ele[14][15];
    ele[5][15] != ele[15][15];
    ele[5][15] != ele[16][15];
    ele[5][15] != ele[17][15];
    ele[5][15] != ele[18][15];
    ele[5][15] != ele[19][15];
    ele[5][15] != ele[20][15];
    ele[5][15] != ele[21][15];
    ele[5][15] != ele[22][15];
    ele[5][15] != ele[23][15];
    ele[5][15] != ele[24][15];
    ele[5][15] != ele[5][16];
    ele[5][15] != ele[5][17];
    ele[5][15] != ele[5][18];
    ele[5][15] != ele[5][19];
    ele[5][15] != ele[5][20];
    ele[5][15] != ele[5][21];
    ele[5][15] != ele[5][22];
    ele[5][15] != ele[5][23];
    ele[5][15] != ele[5][24];
    ele[5][15] != ele[6][15];
    ele[5][15] != ele[6][16];
    ele[5][15] != ele[6][17];
    ele[5][15] != ele[6][18];
    ele[5][15] != ele[6][19];
    ele[5][15] != ele[7][15];
    ele[5][15] != ele[7][16];
    ele[5][15] != ele[7][17];
    ele[5][15] != ele[7][18];
    ele[5][15] != ele[7][19];
    ele[5][15] != ele[8][15];
    ele[5][15] != ele[8][16];
    ele[5][15] != ele[8][17];
    ele[5][15] != ele[8][18];
    ele[5][15] != ele[8][19];
    ele[5][15] != ele[9][15];
    ele[5][15] != ele[9][16];
    ele[5][15] != ele[9][17];
    ele[5][15] != ele[9][18];
    ele[5][15] != ele[9][19];
    ele[5][16] != ele[10][16];
    ele[5][16] != ele[11][16];
    ele[5][16] != ele[12][16];
    ele[5][16] != ele[13][16];
    ele[5][16] != ele[14][16];
    ele[5][16] != ele[15][16];
    ele[5][16] != ele[16][16];
    ele[5][16] != ele[17][16];
    ele[5][16] != ele[18][16];
    ele[5][16] != ele[19][16];
    ele[5][16] != ele[20][16];
    ele[5][16] != ele[21][16];
    ele[5][16] != ele[22][16];
    ele[5][16] != ele[23][16];
    ele[5][16] != ele[24][16];
    ele[5][16] != ele[5][17];
    ele[5][16] != ele[5][18];
    ele[5][16] != ele[5][19];
    ele[5][16] != ele[5][20];
    ele[5][16] != ele[5][21];
    ele[5][16] != ele[5][22];
    ele[5][16] != ele[5][23];
    ele[5][16] != ele[5][24];
    ele[5][16] != ele[6][15];
    ele[5][16] != ele[6][16];
    ele[5][16] != ele[6][17];
    ele[5][16] != ele[6][18];
    ele[5][16] != ele[6][19];
    ele[5][16] != ele[7][15];
    ele[5][16] != ele[7][16];
    ele[5][16] != ele[7][17];
    ele[5][16] != ele[7][18];
    ele[5][16] != ele[7][19];
    ele[5][16] != ele[8][15];
    ele[5][16] != ele[8][16];
    ele[5][16] != ele[8][17];
    ele[5][16] != ele[8][18];
    ele[5][16] != ele[8][19];
    ele[5][16] != ele[9][15];
    ele[5][16] != ele[9][16];
    ele[5][16] != ele[9][17];
    ele[5][16] != ele[9][18];
    ele[5][16] != ele[9][19];
    ele[5][17] != ele[10][17];
    ele[5][17] != ele[11][17];
    ele[5][17] != ele[12][17];
    ele[5][17] != ele[13][17];
    ele[5][17] != ele[14][17];
    ele[5][17] != ele[15][17];
    ele[5][17] != ele[16][17];
    ele[5][17] != ele[17][17];
    ele[5][17] != ele[18][17];
    ele[5][17] != ele[19][17];
    ele[5][17] != ele[20][17];
    ele[5][17] != ele[21][17];
    ele[5][17] != ele[22][17];
    ele[5][17] != ele[23][17];
    ele[5][17] != ele[24][17];
    ele[5][17] != ele[5][18];
    ele[5][17] != ele[5][19];
    ele[5][17] != ele[5][20];
    ele[5][17] != ele[5][21];
    ele[5][17] != ele[5][22];
    ele[5][17] != ele[5][23];
    ele[5][17] != ele[5][24];
    ele[5][17] != ele[6][15];
    ele[5][17] != ele[6][16];
    ele[5][17] != ele[6][17];
    ele[5][17] != ele[6][18];
    ele[5][17] != ele[6][19];
    ele[5][17] != ele[7][15];
    ele[5][17] != ele[7][16];
    ele[5][17] != ele[7][17];
    ele[5][17] != ele[7][18];
    ele[5][17] != ele[7][19];
    ele[5][17] != ele[8][15];
    ele[5][17] != ele[8][16];
    ele[5][17] != ele[8][17];
    ele[5][17] != ele[8][18];
    ele[5][17] != ele[8][19];
    ele[5][17] != ele[9][15];
    ele[5][17] != ele[9][16];
    ele[5][17] != ele[9][17];
    ele[5][17] != ele[9][18];
    ele[5][17] != ele[9][19];
    ele[5][18] != ele[10][18];
    ele[5][18] != ele[11][18];
    ele[5][18] != ele[12][18];
    ele[5][18] != ele[13][18];
    ele[5][18] != ele[14][18];
    ele[5][18] != ele[15][18];
    ele[5][18] != ele[16][18];
    ele[5][18] != ele[17][18];
    ele[5][18] != ele[18][18];
    ele[5][18] != ele[19][18];
    ele[5][18] != ele[20][18];
    ele[5][18] != ele[21][18];
    ele[5][18] != ele[22][18];
    ele[5][18] != ele[23][18];
    ele[5][18] != ele[24][18];
    ele[5][18] != ele[5][19];
    ele[5][18] != ele[5][20];
    ele[5][18] != ele[5][21];
    ele[5][18] != ele[5][22];
    ele[5][18] != ele[5][23];
    ele[5][18] != ele[5][24];
    ele[5][18] != ele[6][15];
    ele[5][18] != ele[6][16];
    ele[5][18] != ele[6][17];
    ele[5][18] != ele[6][18];
    ele[5][18] != ele[6][19];
    ele[5][18] != ele[7][15];
    ele[5][18] != ele[7][16];
    ele[5][18] != ele[7][17];
    ele[5][18] != ele[7][18];
    ele[5][18] != ele[7][19];
    ele[5][18] != ele[8][15];
    ele[5][18] != ele[8][16];
    ele[5][18] != ele[8][17];
    ele[5][18] != ele[8][18];
    ele[5][18] != ele[8][19];
    ele[5][18] != ele[9][15];
    ele[5][18] != ele[9][16];
    ele[5][18] != ele[9][17];
    ele[5][18] != ele[9][18];
    ele[5][18] != ele[9][19];
    ele[5][19] != ele[10][19];
    ele[5][19] != ele[11][19];
    ele[5][19] != ele[12][19];
    ele[5][19] != ele[13][19];
    ele[5][19] != ele[14][19];
    ele[5][19] != ele[15][19];
    ele[5][19] != ele[16][19];
    ele[5][19] != ele[17][19];
    ele[5][19] != ele[18][19];
    ele[5][19] != ele[19][19];
    ele[5][19] != ele[20][19];
    ele[5][19] != ele[21][19];
    ele[5][19] != ele[22][19];
    ele[5][19] != ele[23][19];
    ele[5][19] != ele[24][19];
    ele[5][19] != ele[5][20];
    ele[5][19] != ele[5][21];
    ele[5][19] != ele[5][22];
    ele[5][19] != ele[5][23];
    ele[5][19] != ele[5][24];
    ele[5][19] != ele[6][15];
    ele[5][19] != ele[6][16];
    ele[5][19] != ele[6][17];
    ele[5][19] != ele[6][18];
    ele[5][19] != ele[6][19];
    ele[5][19] != ele[7][15];
    ele[5][19] != ele[7][16];
    ele[5][19] != ele[7][17];
    ele[5][19] != ele[7][18];
    ele[5][19] != ele[7][19];
    ele[5][19] != ele[8][15];
    ele[5][19] != ele[8][16];
    ele[5][19] != ele[8][17];
    ele[5][19] != ele[8][18];
    ele[5][19] != ele[8][19];
    ele[5][19] != ele[9][15];
    ele[5][19] != ele[9][16];
    ele[5][19] != ele[9][17];
    ele[5][19] != ele[9][18];
    ele[5][19] != ele[9][19];
    ele[5][2] != ele[10][2];
    ele[5][2] != ele[11][2];
    ele[5][2] != ele[12][2];
    ele[5][2] != ele[13][2];
    ele[5][2] != ele[14][2];
    ele[5][2] != ele[15][2];
    ele[5][2] != ele[16][2];
    ele[5][2] != ele[17][2];
    ele[5][2] != ele[18][2];
    ele[5][2] != ele[19][2];
    ele[5][2] != ele[20][2];
    ele[5][2] != ele[21][2];
    ele[5][2] != ele[22][2];
    ele[5][2] != ele[23][2];
    ele[5][2] != ele[24][2];
    ele[5][2] != ele[5][10];
    ele[5][2] != ele[5][11];
    ele[5][2] != ele[5][12];
    ele[5][2] != ele[5][13];
    ele[5][2] != ele[5][14];
    ele[5][2] != ele[5][15];
    ele[5][2] != ele[5][16];
    ele[5][2] != ele[5][17];
    ele[5][2] != ele[5][18];
    ele[5][2] != ele[5][19];
    ele[5][2] != ele[5][20];
    ele[5][2] != ele[5][21];
    ele[5][2] != ele[5][22];
    ele[5][2] != ele[5][23];
    ele[5][2] != ele[5][24];
    ele[5][2] != ele[5][3];
    ele[5][2] != ele[5][4];
    ele[5][2] != ele[5][5];
    ele[5][2] != ele[5][6];
    ele[5][2] != ele[5][7];
    ele[5][2] != ele[5][8];
    ele[5][2] != ele[5][9];
    ele[5][2] != ele[6][0];
    ele[5][2] != ele[6][1];
    ele[5][2] != ele[6][2];
    ele[5][2] != ele[6][3];
    ele[5][2] != ele[6][4];
    ele[5][2] != ele[7][0];
    ele[5][2] != ele[7][1];
    ele[5][2] != ele[7][2];
    ele[5][2] != ele[7][3];
    ele[5][2] != ele[7][4];
    ele[5][2] != ele[8][0];
    ele[5][2] != ele[8][1];
    ele[5][2] != ele[8][2];
    ele[5][2] != ele[8][3];
    ele[5][2] != ele[8][4];
    ele[5][2] != ele[9][0];
    ele[5][2] != ele[9][1];
    ele[5][2] != ele[9][2];
    ele[5][2] != ele[9][3];
    ele[5][2] != ele[9][4];
    ele[5][20] != ele[10][20];
    ele[5][20] != ele[11][20];
    ele[5][20] != ele[12][20];
    ele[5][20] != ele[13][20];
    ele[5][20] != ele[14][20];
    ele[5][20] != ele[15][20];
    ele[5][20] != ele[16][20];
    ele[5][20] != ele[17][20];
    ele[5][20] != ele[18][20];
    ele[5][20] != ele[19][20];
    ele[5][20] != ele[20][20];
    ele[5][20] != ele[21][20];
    ele[5][20] != ele[22][20];
    ele[5][20] != ele[23][20];
    ele[5][20] != ele[24][20];
    ele[5][20] != ele[5][21];
    ele[5][20] != ele[5][22];
    ele[5][20] != ele[5][23];
    ele[5][20] != ele[5][24];
    ele[5][20] != ele[6][20];
    ele[5][20] != ele[6][21];
    ele[5][20] != ele[6][22];
    ele[5][20] != ele[6][23];
    ele[5][20] != ele[6][24];
    ele[5][20] != ele[7][20];
    ele[5][20] != ele[7][21];
    ele[5][20] != ele[7][22];
    ele[5][20] != ele[7][23];
    ele[5][20] != ele[7][24];
    ele[5][20] != ele[8][20];
    ele[5][20] != ele[8][21];
    ele[5][20] != ele[8][22];
    ele[5][20] != ele[8][23];
    ele[5][20] != ele[8][24];
    ele[5][20] != ele[9][20];
    ele[5][20] != ele[9][21];
    ele[5][20] != ele[9][22];
    ele[5][20] != ele[9][23];
    ele[5][20] != ele[9][24];
    ele[5][21] != ele[10][21];
    ele[5][21] != ele[11][21];
    ele[5][21] != ele[12][21];
    ele[5][21] != ele[13][21];
    ele[5][21] != ele[14][21];
    ele[5][21] != ele[15][21];
    ele[5][21] != ele[16][21];
    ele[5][21] != ele[17][21];
    ele[5][21] != ele[18][21];
    ele[5][21] != ele[19][21];
    ele[5][21] != ele[20][21];
    ele[5][21] != ele[21][21];
    ele[5][21] != ele[22][21];
    ele[5][21] != ele[23][21];
    ele[5][21] != ele[24][21];
    ele[5][21] != ele[5][22];
    ele[5][21] != ele[5][23];
    ele[5][21] != ele[5][24];
    ele[5][21] != ele[6][20];
    ele[5][21] != ele[6][21];
    ele[5][21] != ele[6][22];
    ele[5][21] != ele[6][23];
    ele[5][21] != ele[6][24];
    ele[5][21] != ele[7][20];
    ele[5][21] != ele[7][21];
    ele[5][21] != ele[7][22];
    ele[5][21] != ele[7][23];
    ele[5][21] != ele[7][24];
    ele[5][21] != ele[8][20];
    ele[5][21] != ele[8][21];
    ele[5][21] != ele[8][22];
    ele[5][21] != ele[8][23];
    ele[5][21] != ele[8][24];
    ele[5][21] != ele[9][20];
    ele[5][21] != ele[9][21];
    ele[5][21] != ele[9][22];
    ele[5][21] != ele[9][23];
    ele[5][21] != ele[9][24];
    ele[5][22] != ele[10][22];
    ele[5][22] != ele[11][22];
    ele[5][22] != ele[12][22];
    ele[5][22] != ele[13][22];
    ele[5][22] != ele[14][22];
    ele[5][22] != ele[15][22];
    ele[5][22] != ele[16][22];
    ele[5][22] != ele[17][22];
    ele[5][22] != ele[18][22];
    ele[5][22] != ele[19][22];
    ele[5][22] != ele[20][22];
    ele[5][22] != ele[21][22];
    ele[5][22] != ele[22][22];
    ele[5][22] != ele[23][22];
    ele[5][22] != ele[24][22];
    ele[5][22] != ele[5][23];
    ele[5][22] != ele[5][24];
    ele[5][22] != ele[6][20];
    ele[5][22] != ele[6][21];
    ele[5][22] != ele[6][22];
    ele[5][22] != ele[6][23];
    ele[5][22] != ele[6][24];
    ele[5][22] != ele[7][20];
    ele[5][22] != ele[7][21];
    ele[5][22] != ele[7][22];
    ele[5][22] != ele[7][23];
    ele[5][22] != ele[7][24];
    ele[5][22] != ele[8][20];
    ele[5][22] != ele[8][21];
    ele[5][22] != ele[8][22];
    ele[5][22] != ele[8][23];
    ele[5][22] != ele[8][24];
    ele[5][22] != ele[9][20];
    ele[5][22] != ele[9][21];
    ele[5][22] != ele[9][22];
    ele[5][22] != ele[9][23];
    ele[5][22] != ele[9][24];
    ele[5][23] != ele[10][23];
    ele[5][23] != ele[11][23];
    ele[5][23] != ele[12][23];
    ele[5][23] != ele[13][23];
    ele[5][23] != ele[14][23];
    ele[5][23] != ele[15][23];
    ele[5][23] != ele[16][23];
    ele[5][23] != ele[17][23];
    ele[5][23] != ele[18][23];
    ele[5][23] != ele[19][23];
    ele[5][23] != ele[20][23];
    ele[5][23] != ele[21][23];
    ele[5][23] != ele[22][23];
    ele[5][23] != ele[23][23];
    ele[5][23] != ele[24][23];
    ele[5][23] != ele[5][24];
    ele[5][23] != ele[6][20];
    ele[5][23] != ele[6][21];
    ele[5][23] != ele[6][22];
    ele[5][23] != ele[6][23];
    ele[5][23] != ele[6][24];
    ele[5][23] != ele[7][20];
    ele[5][23] != ele[7][21];
    ele[5][23] != ele[7][22];
    ele[5][23] != ele[7][23];
    ele[5][23] != ele[7][24];
    ele[5][23] != ele[8][20];
    ele[5][23] != ele[8][21];
    ele[5][23] != ele[8][22];
    ele[5][23] != ele[8][23];
    ele[5][23] != ele[8][24];
    ele[5][23] != ele[9][20];
    ele[5][23] != ele[9][21];
    ele[5][23] != ele[9][22];
    ele[5][23] != ele[9][23];
    ele[5][23] != ele[9][24];
    ele[5][24] != ele[10][24];
    ele[5][24] != ele[11][24];
    ele[5][24] != ele[12][24];
    ele[5][24] != ele[13][24];
    ele[5][24] != ele[14][24];
    ele[5][24] != ele[15][24];
    ele[5][24] != ele[16][24];
    ele[5][24] != ele[17][24];
    ele[5][24] != ele[18][24];
    ele[5][24] != ele[19][24];
    ele[5][24] != ele[20][24];
    ele[5][24] != ele[21][24];
    ele[5][24] != ele[22][24];
    ele[5][24] != ele[23][24];
    ele[5][24] != ele[24][24];
    ele[5][24] != ele[6][20];
    ele[5][24] != ele[6][21];
    ele[5][24] != ele[6][22];
    ele[5][24] != ele[6][23];
    ele[5][24] != ele[6][24];
    ele[5][24] != ele[7][20];
    ele[5][24] != ele[7][21];
    ele[5][24] != ele[7][22];
    ele[5][24] != ele[7][23];
    ele[5][24] != ele[7][24];
    ele[5][24] != ele[8][20];
    ele[5][24] != ele[8][21];
    ele[5][24] != ele[8][22];
    ele[5][24] != ele[8][23];
    ele[5][24] != ele[8][24];
    ele[5][24] != ele[9][20];
    ele[5][24] != ele[9][21];
    ele[5][24] != ele[9][22];
    ele[5][24] != ele[9][23];
    ele[5][24] != ele[9][24];
    ele[5][3] != ele[10][3];
    ele[5][3] != ele[11][3];
    ele[5][3] != ele[12][3];
    ele[5][3] != ele[13][3];
    ele[5][3] != ele[14][3];
    ele[5][3] != ele[15][3];
    ele[5][3] != ele[16][3];
    ele[5][3] != ele[17][3];
    ele[5][3] != ele[18][3];
    ele[5][3] != ele[19][3];
    ele[5][3] != ele[20][3];
    ele[5][3] != ele[21][3];
    ele[5][3] != ele[22][3];
    ele[5][3] != ele[23][3];
    ele[5][3] != ele[24][3];
    ele[5][3] != ele[5][10];
    ele[5][3] != ele[5][11];
    ele[5][3] != ele[5][12];
    ele[5][3] != ele[5][13];
    ele[5][3] != ele[5][14];
    ele[5][3] != ele[5][15];
    ele[5][3] != ele[5][16];
    ele[5][3] != ele[5][17];
    ele[5][3] != ele[5][18];
    ele[5][3] != ele[5][19];
    ele[5][3] != ele[5][20];
    ele[5][3] != ele[5][21];
    ele[5][3] != ele[5][22];
    ele[5][3] != ele[5][23];
    ele[5][3] != ele[5][24];
    ele[5][3] != ele[5][4];
    ele[5][3] != ele[5][5];
    ele[5][3] != ele[5][6];
    ele[5][3] != ele[5][7];
    ele[5][3] != ele[5][8];
    ele[5][3] != ele[5][9];
    ele[5][3] != ele[6][0];
    ele[5][3] != ele[6][1];
    ele[5][3] != ele[6][2];
    ele[5][3] != ele[6][3];
    ele[5][3] != ele[6][4];
    ele[5][3] != ele[7][0];
    ele[5][3] != ele[7][1];
    ele[5][3] != ele[7][2];
    ele[5][3] != ele[7][3];
    ele[5][3] != ele[7][4];
    ele[5][3] != ele[8][0];
    ele[5][3] != ele[8][1];
    ele[5][3] != ele[8][2];
    ele[5][3] != ele[8][3];
    ele[5][3] != ele[8][4];
    ele[5][3] != ele[9][0];
    ele[5][3] != ele[9][1];
    ele[5][3] != ele[9][2];
    ele[5][3] != ele[9][3];
    ele[5][3] != ele[9][4];
    ele[5][4] != ele[10][4];
    ele[5][4] != ele[11][4];
    ele[5][4] != ele[12][4];
    ele[5][4] != ele[13][4];
    ele[5][4] != ele[14][4];
    ele[5][4] != ele[15][4];
    ele[5][4] != ele[16][4];
    ele[5][4] != ele[17][4];
    ele[5][4] != ele[18][4];
    ele[5][4] != ele[19][4];
    ele[5][4] != ele[20][4];
    ele[5][4] != ele[21][4];
    ele[5][4] != ele[22][4];
    ele[5][4] != ele[23][4];
    ele[5][4] != ele[24][4];
    ele[5][4] != ele[5][10];
    ele[5][4] != ele[5][11];
    ele[5][4] != ele[5][12];
    ele[5][4] != ele[5][13];
    ele[5][4] != ele[5][14];
    ele[5][4] != ele[5][15];
    ele[5][4] != ele[5][16];
    ele[5][4] != ele[5][17];
    ele[5][4] != ele[5][18];
    ele[5][4] != ele[5][19];
    ele[5][4] != ele[5][20];
    ele[5][4] != ele[5][21];
    ele[5][4] != ele[5][22];
    ele[5][4] != ele[5][23];
    ele[5][4] != ele[5][24];
    ele[5][4] != ele[5][5];
    ele[5][4] != ele[5][6];
    ele[5][4] != ele[5][7];
    ele[5][4] != ele[5][8];
    ele[5][4] != ele[5][9];
    ele[5][4] != ele[6][0];
    ele[5][4] != ele[6][1];
    ele[5][4] != ele[6][2];
    ele[5][4] != ele[6][3];
    ele[5][4] != ele[6][4];
    ele[5][4] != ele[7][0];
    ele[5][4] != ele[7][1];
    ele[5][4] != ele[7][2];
    ele[5][4] != ele[7][3];
    ele[5][4] != ele[7][4];
    ele[5][4] != ele[8][0];
    ele[5][4] != ele[8][1];
    ele[5][4] != ele[8][2];
    ele[5][4] != ele[8][3];
    ele[5][4] != ele[8][4];
    ele[5][4] != ele[9][0];
    ele[5][4] != ele[9][1];
    ele[5][4] != ele[9][2];
    ele[5][4] != ele[9][3];
    ele[5][4] != ele[9][4];
    ele[5][5] != ele[10][5];
    ele[5][5] != ele[11][5];
    ele[5][5] != ele[12][5];
    ele[5][5] != ele[13][5];
    ele[5][5] != ele[14][5];
    ele[5][5] != ele[15][5];
    ele[5][5] != ele[16][5];
    ele[5][5] != ele[17][5];
    ele[5][5] != ele[18][5];
    ele[5][5] != ele[19][5];
    ele[5][5] != ele[20][5];
    ele[5][5] != ele[21][5];
    ele[5][5] != ele[22][5];
    ele[5][5] != ele[23][5];
    ele[5][5] != ele[24][5];
    ele[5][5] != ele[5][10];
    ele[5][5] != ele[5][11];
    ele[5][5] != ele[5][12];
    ele[5][5] != ele[5][13];
    ele[5][5] != ele[5][14];
    ele[5][5] != ele[5][15];
    ele[5][5] != ele[5][16];
    ele[5][5] != ele[5][17];
    ele[5][5] != ele[5][18];
    ele[5][5] != ele[5][19];
    ele[5][5] != ele[5][20];
    ele[5][5] != ele[5][21];
    ele[5][5] != ele[5][22];
    ele[5][5] != ele[5][23];
    ele[5][5] != ele[5][24];
    ele[5][5] != ele[5][6];
    ele[5][5] != ele[5][7];
    ele[5][5] != ele[5][8];
    ele[5][5] != ele[5][9];
    ele[5][5] != ele[6][5];
    ele[5][5] != ele[6][6];
    ele[5][5] != ele[6][7];
    ele[5][5] != ele[6][8];
    ele[5][5] != ele[6][9];
    ele[5][5] != ele[7][5];
    ele[5][5] != ele[7][6];
    ele[5][5] != ele[7][7];
    ele[5][5] != ele[7][8];
    ele[5][5] != ele[7][9];
    ele[5][5] != ele[8][5];
    ele[5][5] != ele[8][6];
    ele[5][5] != ele[8][7];
    ele[5][5] != ele[8][8];
    ele[5][5] != ele[8][9];
    ele[5][5] != ele[9][5];
    ele[5][5] != ele[9][6];
    ele[5][5] != ele[9][7];
    ele[5][5] != ele[9][8];
    ele[5][5] != ele[9][9];
    ele[5][6] != ele[10][6];
    ele[5][6] != ele[11][6];
    ele[5][6] != ele[12][6];
    ele[5][6] != ele[13][6];
    ele[5][6] != ele[14][6];
    ele[5][6] != ele[15][6];
    ele[5][6] != ele[16][6];
    ele[5][6] != ele[17][6];
    ele[5][6] != ele[18][6];
    ele[5][6] != ele[19][6];
    ele[5][6] != ele[20][6];
    ele[5][6] != ele[21][6];
    ele[5][6] != ele[22][6];
    ele[5][6] != ele[23][6];
    ele[5][6] != ele[24][6];
    ele[5][6] != ele[5][10];
    ele[5][6] != ele[5][11];
    ele[5][6] != ele[5][12];
    ele[5][6] != ele[5][13];
    ele[5][6] != ele[5][14];
    ele[5][6] != ele[5][15];
    ele[5][6] != ele[5][16];
    ele[5][6] != ele[5][17];
    ele[5][6] != ele[5][18];
    ele[5][6] != ele[5][19];
    ele[5][6] != ele[5][20];
    ele[5][6] != ele[5][21];
    ele[5][6] != ele[5][22];
    ele[5][6] != ele[5][23];
    ele[5][6] != ele[5][24];
    ele[5][6] != ele[5][7];
    ele[5][6] != ele[5][8];
    ele[5][6] != ele[5][9];
    ele[5][6] != ele[6][5];
    ele[5][6] != ele[6][6];
    ele[5][6] != ele[6][7];
    ele[5][6] != ele[6][8];
    ele[5][6] != ele[6][9];
    ele[5][6] != ele[7][5];
    ele[5][6] != ele[7][6];
    ele[5][6] != ele[7][7];
    ele[5][6] != ele[7][8];
    ele[5][6] != ele[7][9];
    ele[5][6] != ele[8][5];
    ele[5][6] != ele[8][6];
    ele[5][6] != ele[8][7];
    ele[5][6] != ele[8][8];
    ele[5][6] != ele[8][9];
    ele[5][6] != ele[9][5];
    ele[5][6] != ele[9][6];
    ele[5][6] != ele[9][7];
    ele[5][6] != ele[9][8];
    ele[5][6] != ele[9][9];
    ele[5][7] != ele[10][7];
    ele[5][7] != ele[11][7];
    ele[5][7] != ele[12][7];
    ele[5][7] != ele[13][7];
    ele[5][7] != ele[14][7];
    ele[5][7] != ele[15][7];
    ele[5][7] != ele[16][7];
    ele[5][7] != ele[17][7];
    ele[5][7] != ele[18][7];
    ele[5][7] != ele[19][7];
    ele[5][7] != ele[20][7];
    ele[5][7] != ele[21][7];
    ele[5][7] != ele[22][7];
    ele[5][7] != ele[23][7];
    ele[5][7] != ele[24][7];
    ele[5][7] != ele[5][10];
    ele[5][7] != ele[5][11];
    ele[5][7] != ele[5][12];
    ele[5][7] != ele[5][13];
    ele[5][7] != ele[5][14];
    ele[5][7] != ele[5][15];
    ele[5][7] != ele[5][16];
    ele[5][7] != ele[5][17];
    ele[5][7] != ele[5][18];
    ele[5][7] != ele[5][19];
    ele[5][7] != ele[5][20];
    ele[5][7] != ele[5][21];
    ele[5][7] != ele[5][22];
    ele[5][7] != ele[5][23];
    ele[5][7] != ele[5][24];
    ele[5][7] != ele[5][8];
    ele[5][7] != ele[5][9];
    ele[5][7] != ele[6][5];
    ele[5][7] != ele[6][6];
    ele[5][7] != ele[6][7];
    ele[5][7] != ele[6][8];
    ele[5][7] != ele[6][9];
    ele[5][7] != ele[7][5];
    ele[5][7] != ele[7][6];
    ele[5][7] != ele[7][7];
    ele[5][7] != ele[7][8];
    ele[5][7] != ele[7][9];
    ele[5][7] != ele[8][5];
    ele[5][7] != ele[8][6];
    ele[5][7] != ele[8][7];
    ele[5][7] != ele[8][8];
    ele[5][7] != ele[8][9];
    ele[5][7] != ele[9][5];
    ele[5][7] != ele[9][6];
    ele[5][7] != ele[9][7];
    ele[5][7] != ele[9][8];
    ele[5][7] != ele[9][9];
    ele[5][8] != ele[10][8];
    ele[5][8] != ele[11][8];
    ele[5][8] != ele[12][8];
    ele[5][8] != ele[13][8];
    ele[5][8] != ele[14][8];
    ele[5][8] != ele[15][8];
    ele[5][8] != ele[16][8];
    ele[5][8] != ele[17][8];
    ele[5][8] != ele[18][8];
    ele[5][8] != ele[19][8];
    ele[5][8] != ele[20][8];
    ele[5][8] != ele[21][8];
    ele[5][8] != ele[22][8];
    ele[5][8] != ele[23][8];
    ele[5][8] != ele[24][8];
    ele[5][8] != ele[5][10];
    ele[5][8] != ele[5][11];
    ele[5][8] != ele[5][12];
    ele[5][8] != ele[5][13];
    ele[5][8] != ele[5][14];
    ele[5][8] != ele[5][15];
    ele[5][8] != ele[5][16];
    ele[5][8] != ele[5][17];
    ele[5][8] != ele[5][18];
    ele[5][8] != ele[5][19];
    ele[5][8] != ele[5][20];
    ele[5][8] != ele[5][21];
    ele[5][8] != ele[5][22];
    ele[5][8] != ele[5][23];
    ele[5][8] != ele[5][24];
    ele[5][8] != ele[5][9];
    ele[5][8] != ele[6][5];
    ele[5][8] != ele[6][6];
    ele[5][8] != ele[6][7];
    ele[5][8] != ele[6][8];
    ele[5][8] != ele[6][9];
    ele[5][8] != ele[7][5];
    ele[5][8] != ele[7][6];
    ele[5][8] != ele[7][7];
    ele[5][8] != ele[7][8];
    ele[5][8] != ele[7][9];
    ele[5][8] != ele[8][5];
    ele[5][8] != ele[8][6];
    ele[5][8] != ele[8][7];
    ele[5][8] != ele[8][8];
    ele[5][8] != ele[8][9];
    ele[5][8] != ele[9][5];
    ele[5][8] != ele[9][6];
    ele[5][8] != ele[9][7];
    ele[5][8] != ele[9][8];
    ele[5][8] != ele[9][9];
    ele[5][9] != ele[10][9];
    ele[5][9] != ele[11][9];
    ele[5][9] != ele[12][9];
    ele[5][9] != ele[13][9];
    ele[5][9] != ele[14][9];
    ele[5][9] != ele[15][9];
    ele[5][9] != ele[16][9];
    ele[5][9] != ele[17][9];
    ele[5][9] != ele[18][9];
    ele[5][9] != ele[19][9];
    ele[5][9] != ele[20][9];
    ele[5][9] != ele[21][9];
    ele[5][9] != ele[22][9];
    ele[5][9] != ele[23][9];
    ele[5][9] != ele[24][9];
    ele[5][9] != ele[5][10];
    ele[5][9] != ele[5][11];
    ele[5][9] != ele[5][12];
    ele[5][9] != ele[5][13];
    ele[5][9] != ele[5][14];
    ele[5][9] != ele[5][15];
    ele[5][9] != ele[5][16];
    ele[5][9] != ele[5][17];
    ele[5][9] != ele[5][18];
    ele[5][9] != ele[5][19];
    ele[5][9] != ele[5][20];
    ele[5][9] != ele[5][21];
    ele[5][9] != ele[5][22];
    ele[5][9] != ele[5][23];
    ele[5][9] != ele[5][24];
    ele[5][9] != ele[6][5];
    ele[5][9] != ele[6][6];
    ele[5][9] != ele[6][7];
    ele[5][9] != ele[6][8];
    ele[5][9] != ele[6][9];
    ele[5][9] != ele[7][5];
    ele[5][9] != ele[7][6];
    ele[5][9] != ele[7][7];
    ele[5][9] != ele[7][8];
    ele[5][9] != ele[7][9];
    ele[5][9] != ele[8][5];
    ele[5][9] != ele[8][6];
    ele[5][9] != ele[8][7];
    ele[5][9] != ele[8][8];
    ele[5][9] != ele[8][9];
    ele[5][9] != ele[9][5];
    ele[5][9] != ele[9][6];
    ele[5][9] != ele[9][7];
    ele[5][9] != ele[9][8];
    ele[5][9] != ele[9][9];
    ele[6][0] != ele[10][0];
    ele[6][0] != ele[11][0];
    ele[6][0] != ele[12][0];
    ele[6][0] != ele[13][0];
    ele[6][0] != ele[14][0];
    ele[6][0] != ele[15][0];
    ele[6][0] != ele[16][0];
    ele[6][0] != ele[17][0];
    ele[6][0] != ele[18][0];
    ele[6][0] != ele[19][0];
    ele[6][0] != ele[20][0];
    ele[6][0] != ele[21][0];
    ele[6][0] != ele[22][0];
    ele[6][0] != ele[23][0];
    ele[6][0] != ele[24][0];
    ele[6][0] != ele[6][1];
    ele[6][0] != ele[6][10];
    ele[6][0] != ele[6][11];
    ele[6][0] != ele[6][12];
    ele[6][0] != ele[6][13];
    ele[6][0] != ele[6][14];
    ele[6][0] != ele[6][15];
    ele[6][0] != ele[6][16];
    ele[6][0] != ele[6][17];
    ele[6][0] != ele[6][18];
    ele[6][0] != ele[6][19];
    ele[6][0] != ele[6][2];
    ele[6][0] != ele[6][20];
    ele[6][0] != ele[6][21];
    ele[6][0] != ele[6][22];
    ele[6][0] != ele[6][23];
    ele[6][0] != ele[6][24];
    ele[6][0] != ele[6][3];
    ele[6][0] != ele[6][4];
    ele[6][0] != ele[6][5];
    ele[6][0] != ele[6][6];
    ele[6][0] != ele[6][7];
    ele[6][0] != ele[6][8];
    ele[6][0] != ele[6][9];
    ele[6][0] != ele[7][0];
    ele[6][0] != ele[7][1];
    ele[6][0] != ele[7][2];
    ele[6][0] != ele[7][3];
    ele[6][0] != ele[7][4];
    ele[6][0] != ele[8][0];
    ele[6][0] != ele[8][1];
    ele[6][0] != ele[8][2];
    ele[6][0] != ele[8][3];
    ele[6][0] != ele[8][4];
    ele[6][0] != ele[9][0];
    ele[6][0] != ele[9][1];
    ele[6][0] != ele[9][2];
    ele[6][0] != ele[9][3];
    ele[6][0] != ele[9][4];
    ele[6][1] != ele[10][1];
    ele[6][1] != ele[11][1];
    ele[6][1] != ele[12][1];
    ele[6][1] != ele[13][1];
    ele[6][1] != ele[14][1];
    ele[6][1] != ele[15][1];
    ele[6][1] != ele[16][1];
    ele[6][1] != ele[17][1];
    ele[6][1] != ele[18][1];
    ele[6][1] != ele[19][1];
    ele[6][1] != ele[20][1];
    ele[6][1] != ele[21][1];
    ele[6][1] != ele[22][1];
    ele[6][1] != ele[23][1];
    ele[6][1] != ele[24][1];
    ele[6][1] != ele[6][10];
    ele[6][1] != ele[6][11];
    ele[6][1] != ele[6][12];
    ele[6][1] != ele[6][13];
    ele[6][1] != ele[6][14];
    ele[6][1] != ele[6][15];
    ele[6][1] != ele[6][16];
    ele[6][1] != ele[6][17];
    ele[6][1] != ele[6][18];
    ele[6][1] != ele[6][19];
    ele[6][1] != ele[6][2];
    ele[6][1] != ele[6][20];
    ele[6][1] != ele[6][21];
    ele[6][1] != ele[6][22];
    ele[6][1] != ele[6][23];
    ele[6][1] != ele[6][24];
    ele[6][1] != ele[6][3];
    ele[6][1] != ele[6][4];
    ele[6][1] != ele[6][5];
    ele[6][1] != ele[6][6];
    ele[6][1] != ele[6][7];
    ele[6][1] != ele[6][8];
    ele[6][1] != ele[6][9];
    ele[6][1] != ele[7][0];
    ele[6][1] != ele[7][1];
    ele[6][1] != ele[7][2];
    ele[6][1] != ele[7][3];
    ele[6][1] != ele[7][4];
    ele[6][1] != ele[8][0];
    ele[6][1] != ele[8][1];
    ele[6][1] != ele[8][2];
    ele[6][1] != ele[8][3];
    ele[6][1] != ele[8][4];
    ele[6][1] != ele[9][0];
    ele[6][1] != ele[9][1];
    ele[6][1] != ele[9][2];
    ele[6][1] != ele[9][3];
    ele[6][1] != ele[9][4];
    ele[6][10] != ele[10][10];
    ele[6][10] != ele[11][10];
    ele[6][10] != ele[12][10];
    ele[6][10] != ele[13][10];
    ele[6][10] != ele[14][10];
    ele[6][10] != ele[15][10];
    ele[6][10] != ele[16][10];
    ele[6][10] != ele[17][10];
    ele[6][10] != ele[18][10];
    ele[6][10] != ele[19][10];
    ele[6][10] != ele[20][10];
    ele[6][10] != ele[21][10];
    ele[6][10] != ele[22][10];
    ele[6][10] != ele[23][10];
    ele[6][10] != ele[24][10];
    ele[6][10] != ele[6][11];
    ele[6][10] != ele[6][12];
    ele[6][10] != ele[6][13];
    ele[6][10] != ele[6][14];
    ele[6][10] != ele[6][15];
    ele[6][10] != ele[6][16];
    ele[6][10] != ele[6][17];
    ele[6][10] != ele[6][18];
    ele[6][10] != ele[6][19];
    ele[6][10] != ele[6][20];
    ele[6][10] != ele[6][21];
    ele[6][10] != ele[6][22];
    ele[6][10] != ele[6][23];
    ele[6][10] != ele[6][24];
    ele[6][10] != ele[7][10];
    ele[6][10] != ele[7][11];
    ele[6][10] != ele[7][12];
    ele[6][10] != ele[7][13];
    ele[6][10] != ele[7][14];
    ele[6][10] != ele[8][10];
    ele[6][10] != ele[8][11];
    ele[6][10] != ele[8][12];
    ele[6][10] != ele[8][13];
    ele[6][10] != ele[8][14];
    ele[6][10] != ele[9][10];
    ele[6][10] != ele[9][11];
    ele[6][10] != ele[9][12];
    ele[6][10] != ele[9][13];
    ele[6][10] != ele[9][14];
    ele[6][11] != ele[10][11];
    ele[6][11] != ele[11][11];
    ele[6][11] != ele[12][11];
    ele[6][11] != ele[13][11];
    ele[6][11] != ele[14][11];
    ele[6][11] != ele[15][11];
    ele[6][11] != ele[16][11];
    ele[6][11] != ele[17][11];
    ele[6][11] != ele[18][11];
    ele[6][11] != ele[19][11];
    ele[6][11] != ele[20][11];
    ele[6][11] != ele[21][11];
    ele[6][11] != ele[22][11];
    ele[6][11] != ele[23][11];
    ele[6][11] != ele[24][11];
    ele[6][11] != ele[6][12];
    ele[6][11] != ele[6][13];
    ele[6][11] != ele[6][14];
    ele[6][11] != ele[6][15];
    ele[6][11] != ele[6][16];
    ele[6][11] != ele[6][17];
    ele[6][11] != ele[6][18];
    ele[6][11] != ele[6][19];
    ele[6][11] != ele[6][20];
    ele[6][11] != ele[6][21];
    ele[6][11] != ele[6][22];
    ele[6][11] != ele[6][23];
    ele[6][11] != ele[6][24];
    ele[6][11] != ele[7][10];
    ele[6][11] != ele[7][11];
    ele[6][11] != ele[7][12];
    ele[6][11] != ele[7][13];
    ele[6][11] != ele[7][14];
    ele[6][11] != ele[8][10];
    ele[6][11] != ele[8][11];
    ele[6][11] != ele[8][12];
    ele[6][11] != ele[8][13];
    ele[6][11] != ele[8][14];
    ele[6][11] != ele[9][10];
    ele[6][11] != ele[9][11];
    ele[6][11] != ele[9][12];
    ele[6][11] != ele[9][13];
    ele[6][11] != ele[9][14];
    ele[6][12] != ele[10][12];
    ele[6][12] != ele[11][12];
    ele[6][12] != ele[12][12];
    ele[6][12] != ele[13][12];
    ele[6][12] != ele[14][12];
    ele[6][12] != ele[15][12];
    ele[6][12] != ele[16][12];
    ele[6][12] != ele[17][12];
    ele[6][12] != ele[18][12];
    ele[6][12] != ele[19][12];
    ele[6][12] != ele[20][12];
    ele[6][12] != ele[21][12];
    ele[6][12] != ele[22][12];
    ele[6][12] != ele[23][12];
    ele[6][12] != ele[24][12];
    ele[6][12] != ele[6][13];
    ele[6][12] != ele[6][14];
    ele[6][12] != ele[6][15];
    ele[6][12] != ele[6][16];
    ele[6][12] != ele[6][17];
    ele[6][12] != ele[6][18];
    ele[6][12] != ele[6][19];
    ele[6][12] != ele[6][20];
    ele[6][12] != ele[6][21];
    ele[6][12] != ele[6][22];
    ele[6][12] != ele[6][23];
    ele[6][12] != ele[6][24];
    ele[6][12] != ele[7][10];
    ele[6][12] != ele[7][11];
    ele[6][12] != ele[7][12];
    ele[6][12] != ele[7][13];
    ele[6][12] != ele[7][14];
    ele[6][12] != ele[8][10];
    ele[6][12] != ele[8][11];
    ele[6][12] != ele[8][12];
    ele[6][12] != ele[8][13];
    ele[6][12] != ele[8][14];
    ele[6][12] != ele[9][10];
    ele[6][12] != ele[9][11];
    ele[6][12] != ele[9][12];
    ele[6][12] != ele[9][13];
    ele[6][12] != ele[9][14];
    ele[6][13] != ele[10][13];
    ele[6][13] != ele[11][13];
    ele[6][13] != ele[12][13];
    ele[6][13] != ele[13][13];
    ele[6][13] != ele[14][13];
    ele[6][13] != ele[15][13];
    ele[6][13] != ele[16][13];
    ele[6][13] != ele[17][13];
    ele[6][13] != ele[18][13];
    ele[6][13] != ele[19][13];
    ele[6][13] != ele[20][13];
    ele[6][13] != ele[21][13];
    ele[6][13] != ele[22][13];
    ele[6][13] != ele[23][13];
    ele[6][13] != ele[24][13];
    ele[6][13] != ele[6][14];
    ele[6][13] != ele[6][15];
    ele[6][13] != ele[6][16];
    ele[6][13] != ele[6][17];
    ele[6][13] != ele[6][18];
    ele[6][13] != ele[6][19];
    ele[6][13] != ele[6][20];
    ele[6][13] != ele[6][21];
    ele[6][13] != ele[6][22];
    ele[6][13] != ele[6][23];
    ele[6][13] != ele[6][24];
    ele[6][13] != ele[7][10];
    ele[6][13] != ele[7][11];
    ele[6][13] != ele[7][12];
    ele[6][13] != ele[7][13];
    ele[6][13] != ele[7][14];
    ele[6][13] != ele[8][10];
    ele[6][13] != ele[8][11];
    ele[6][13] != ele[8][12];
    ele[6][13] != ele[8][13];
    ele[6][13] != ele[8][14];
    ele[6][13] != ele[9][10];
    ele[6][13] != ele[9][11];
    ele[6][13] != ele[9][12];
    ele[6][13] != ele[9][13];
    ele[6][13] != ele[9][14];
    ele[6][14] != ele[10][14];
    ele[6][14] != ele[11][14];
    ele[6][14] != ele[12][14];
    ele[6][14] != ele[13][14];
    ele[6][14] != ele[14][14];
    ele[6][14] != ele[15][14];
    ele[6][14] != ele[16][14];
    ele[6][14] != ele[17][14];
    ele[6][14] != ele[18][14];
    ele[6][14] != ele[19][14];
    ele[6][14] != ele[20][14];
    ele[6][14] != ele[21][14];
    ele[6][14] != ele[22][14];
    ele[6][14] != ele[23][14];
    ele[6][14] != ele[24][14];
    ele[6][14] != ele[6][15];
    ele[6][14] != ele[6][16];
    ele[6][14] != ele[6][17];
    ele[6][14] != ele[6][18];
    ele[6][14] != ele[6][19];
    ele[6][14] != ele[6][20];
    ele[6][14] != ele[6][21];
    ele[6][14] != ele[6][22];
    ele[6][14] != ele[6][23];
    ele[6][14] != ele[6][24];
    ele[6][14] != ele[7][10];
    ele[6][14] != ele[7][11];
    ele[6][14] != ele[7][12];
    ele[6][14] != ele[7][13];
    ele[6][14] != ele[7][14];
    ele[6][14] != ele[8][10];
    ele[6][14] != ele[8][11];
    ele[6][14] != ele[8][12];
    ele[6][14] != ele[8][13];
    ele[6][14] != ele[8][14];
    ele[6][14] != ele[9][10];
    ele[6][14] != ele[9][11];
    ele[6][14] != ele[9][12];
    ele[6][14] != ele[9][13];
    ele[6][14] != ele[9][14];
    ele[6][15] != ele[10][15];
    ele[6][15] != ele[11][15];
    ele[6][15] != ele[12][15];
    ele[6][15] != ele[13][15];
    ele[6][15] != ele[14][15];
    ele[6][15] != ele[15][15];
    ele[6][15] != ele[16][15];
    ele[6][15] != ele[17][15];
    ele[6][15] != ele[18][15];
    ele[6][15] != ele[19][15];
    ele[6][15] != ele[20][15];
    ele[6][15] != ele[21][15];
    ele[6][15] != ele[22][15];
    ele[6][15] != ele[23][15];
    ele[6][15] != ele[24][15];
    ele[6][15] != ele[6][16];
    ele[6][15] != ele[6][17];
    ele[6][15] != ele[6][18];
    ele[6][15] != ele[6][19];
    ele[6][15] != ele[6][20];
    ele[6][15] != ele[6][21];
    ele[6][15] != ele[6][22];
    ele[6][15] != ele[6][23];
    ele[6][15] != ele[6][24];
    ele[6][15] != ele[7][15];
    ele[6][15] != ele[7][16];
    ele[6][15] != ele[7][17];
    ele[6][15] != ele[7][18];
    ele[6][15] != ele[7][19];
    ele[6][15] != ele[8][15];
    ele[6][15] != ele[8][16];
    ele[6][15] != ele[8][17];
    ele[6][15] != ele[8][18];
    ele[6][15] != ele[8][19];
    ele[6][15] != ele[9][15];
    ele[6][15] != ele[9][16];
    ele[6][15] != ele[9][17];
    ele[6][15] != ele[9][18];
    ele[6][15] != ele[9][19];
    ele[6][16] != ele[10][16];
    ele[6][16] != ele[11][16];
    ele[6][16] != ele[12][16];
    ele[6][16] != ele[13][16];
    ele[6][16] != ele[14][16];
    ele[6][16] != ele[15][16];
    ele[6][16] != ele[16][16];
    ele[6][16] != ele[17][16];
    ele[6][16] != ele[18][16];
    ele[6][16] != ele[19][16];
    ele[6][16] != ele[20][16];
    ele[6][16] != ele[21][16];
    ele[6][16] != ele[22][16];
    ele[6][16] != ele[23][16];
    ele[6][16] != ele[24][16];
    ele[6][16] != ele[6][17];
    ele[6][16] != ele[6][18];
    ele[6][16] != ele[6][19];
    ele[6][16] != ele[6][20];
    ele[6][16] != ele[6][21];
    ele[6][16] != ele[6][22];
    ele[6][16] != ele[6][23];
    ele[6][16] != ele[6][24];
    ele[6][16] != ele[7][15];
    ele[6][16] != ele[7][16];
    ele[6][16] != ele[7][17];
    ele[6][16] != ele[7][18];
    ele[6][16] != ele[7][19];
    ele[6][16] != ele[8][15];
    ele[6][16] != ele[8][16];
    ele[6][16] != ele[8][17];
    ele[6][16] != ele[8][18];
    ele[6][16] != ele[8][19];
    ele[6][16] != ele[9][15];
    ele[6][16] != ele[9][16];
    ele[6][16] != ele[9][17];
    ele[6][16] != ele[9][18];
    ele[6][16] != ele[9][19];
    ele[6][17] != ele[10][17];
    ele[6][17] != ele[11][17];
    ele[6][17] != ele[12][17];
    ele[6][17] != ele[13][17];
    ele[6][17] != ele[14][17];
    ele[6][17] != ele[15][17];
    ele[6][17] != ele[16][17];
    ele[6][17] != ele[17][17];
    ele[6][17] != ele[18][17];
    ele[6][17] != ele[19][17];
    ele[6][17] != ele[20][17];
    ele[6][17] != ele[21][17];
    ele[6][17] != ele[22][17];
    ele[6][17] != ele[23][17];
    ele[6][17] != ele[24][17];
    ele[6][17] != ele[6][18];
    ele[6][17] != ele[6][19];
    ele[6][17] != ele[6][20];
    ele[6][17] != ele[6][21];
    ele[6][17] != ele[6][22];
    ele[6][17] != ele[6][23];
    ele[6][17] != ele[6][24];
    ele[6][17] != ele[7][15];
    ele[6][17] != ele[7][16];
    ele[6][17] != ele[7][17];
    ele[6][17] != ele[7][18];
    ele[6][17] != ele[7][19];
    ele[6][17] != ele[8][15];
    ele[6][17] != ele[8][16];
    ele[6][17] != ele[8][17];
    ele[6][17] != ele[8][18];
    ele[6][17] != ele[8][19];
    ele[6][17] != ele[9][15];
    ele[6][17] != ele[9][16];
    ele[6][17] != ele[9][17];
    ele[6][17] != ele[9][18];
    ele[6][17] != ele[9][19];
    ele[6][18] != ele[10][18];
    ele[6][18] != ele[11][18];
    ele[6][18] != ele[12][18];
    ele[6][18] != ele[13][18];
    ele[6][18] != ele[14][18];
    ele[6][18] != ele[15][18];
    ele[6][18] != ele[16][18];
    ele[6][18] != ele[17][18];
    ele[6][18] != ele[18][18];
    ele[6][18] != ele[19][18];
    ele[6][18] != ele[20][18];
    ele[6][18] != ele[21][18];
    ele[6][18] != ele[22][18];
    ele[6][18] != ele[23][18];
    ele[6][18] != ele[24][18];
    ele[6][18] != ele[6][19];
    ele[6][18] != ele[6][20];
    ele[6][18] != ele[6][21];
    ele[6][18] != ele[6][22];
    ele[6][18] != ele[6][23];
    ele[6][18] != ele[6][24];
    ele[6][18] != ele[7][15];
    ele[6][18] != ele[7][16];
    ele[6][18] != ele[7][17];
    ele[6][18] != ele[7][18];
    ele[6][18] != ele[7][19];
    ele[6][18] != ele[8][15];
    ele[6][18] != ele[8][16];
    ele[6][18] != ele[8][17];
    ele[6][18] != ele[8][18];
    ele[6][18] != ele[8][19];
    ele[6][18] != ele[9][15];
    ele[6][18] != ele[9][16];
    ele[6][18] != ele[9][17];
    ele[6][18] != ele[9][18];
    ele[6][18] != ele[9][19];
    ele[6][19] != ele[10][19];
    ele[6][19] != ele[11][19];
    ele[6][19] != ele[12][19];
    ele[6][19] != ele[13][19];
    ele[6][19] != ele[14][19];
    ele[6][19] != ele[15][19];
    ele[6][19] != ele[16][19];
    ele[6][19] != ele[17][19];
    ele[6][19] != ele[18][19];
    ele[6][19] != ele[19][19];
    ele[6][19] != ele[20][19];
    ele[6][19] != ele[21][19];
    ele[6][19] != ele[22][19];
    ele[6][19] != ele[23][19];
    ele[6][19] != ele[24][19];
    ele[6][19] != ele[6][20];
    ele[6][19] != ele[6][21];
    ele[6][19] != ele[6][22];
    ele[6][19] != ele[6][23];
    ele[6][19] != ele[6][24];
    ele[6][19] != ele[7][15];
    ele[6][19] != ele[7][16];
    ele[6][19] != ele[7][17];
    ele[6][19] != ele[7][18];
    ele[6][19] != ele[7][19];
    ele[6][19] != ele[8][15];
    ele[6][19] != ele[8][16];
    ele[6][19] != ele[8][17];
    ele[6][19] != ele[8][18];
    ele[6][19] != ele[8][19];
    ele[6][19] != ele[9][15];
    ele[6][19] != ele[9][16];
    ele[6][19] != ele[9][17];
    ele[6][19] != ele[9][18];
    ele[6][19] != ele[9][19];
    ele[6][2] != ele[10][2];
    ele[6][2] != ele[11][2];
    ele[6][2] != ele[12][2];
    ele[6][2] != ele[13][2];
    ele[6][2] != ele[14][2];
    ele[6][2] != ele[15][2];
    ele[6][2] != ele[16][2];
    ele[6][2] != ele[17][2];
    ele[6][2] != ele[18][2];
    ele[6][2] != ele[19][2];
    ele[6][2] != ele[20][2];
    ele[6][2] != ele[21][2];
    ele[6][2] != ele[22][2];
    ele[6][2] != ele[23][2];
    ele[6][2] != ele[24][2];
    ele[6][2] != ele[6][10];
    ele[6][2] != ele[6][11];
    ele[6][2] != ele[6][12];
    ele[6][2] != ele[6][13];
    ele[6][2] != ele[6][14];
    ele[6][2] != ele[6][15];
    ele[6][2] != ele[6][16];
    ele[6][2] != ele[6][17];
    ele[6][2] != ele[6][18];
    ele[6][2] != ele[6][19];
    ele[6][2] != ele[6][20];
    ele[6][2] != ele[6][21];
    ele[6][2] != ele[6][22];
    ele[6][2] != ele[6][23];
    ele[6][2] != ele[6][24];
    ele[6][2] != ele[6][3];
    ele[6][2] != ele[6][4];
    ele[6][2] != ele[6][5];
    ele[6][2] != ele[6][6];
    ele[6][2] != ele[6][7];
    ele[6][2] != ele[6][8];
    ele[6][2] != ele[6][9];
    ele[6][2] != ele[7][0];
    ele[6][2] != ele[7][1];
    ele[6][2] != ele[7][2];
    ele[6][2] != ele[7][3];
    ele[6][2] != ele[7][4];
    ele[6][2] != ele[8][0];
    ele[6][2] != ele[8][1];
    ele[6][2] != ele[8][2];
    ele[6][2] != ele[8][3];
    ele[6][2] != ele[8][4];
    ele[6][2] != ele[9][0];
    ele[6][2] != ele[9][1];
    ele[6][2] != ele[9][2];
    ele[6][2] != ele[9][3];
    ele[6][2] != ele[9][4];
    ele[6][20] != ele[10][20];
    ele[6][20] != ele[11][20];
    ele[6][20] != ele[12][20];
    ele[6][20] != ele[13][20];
    ele[6][20] != ele[14][20];
    ele[6][20] != ele[15][20];
    ele[6][20] != ele[16][20];
    ele[6][20] != ele[17][20];
    ele[6][20] != ele[18][20];
    ele[6][20] != ele[19][20];
    ele[6][20] != ele[20][20];
    ele[6][20] != ele[21][20];
    ele[6][20] != ele[22][20];
    ele[6][20] != ele[23][20];
    ele[6][20] != ele[24][20];
    ele[6][20] != ele[6][21];
    ele[6][20] != ele[6][22];
    ele[6][20] != ele[6][23];
    ele[6][20] != ele[6][24];
    ele[6][20] != ele[7][20];
    ele[6][20] != ele[7][21];
    ele[6][20] != ele[7][22];
    ele[6][20] != ele[7][23];
    ele[6][20] != ele[7][24];
    ele[6][20] != ele[8][20];
    ele[6][20] != ele[8][21];
    ele[6][20] != ele[8][22];
    ele[6][20] != ele[8][23];
    ele[6][20] != ele[8][24];
    ele[6][20] != ele[9][20];
    ele[6][20] != ele[9][21];
    ele[6][20] != ele[9][22];
    ele[6][20] != ele[9][23];
    ele[6][20] != ele[9][24];
    ele[6][21] != ele[10][21];
    ele[6][21] != ele[11][21];
    ele[6][21] != ele[12][21];
    ele[6][21] != ele[13][21];
    ele[6][21] != ele[14][21];
    ele[6][21] != ele[15][21];
    ele[6][21] != ele[16][21];
    ele[6][21] != ele[17][21];
    ele[6][21] != ele[18][21];
    ele[6][21] != ele[19][21];
    ele[6][21] != ele[20][21];
    ele[6][21] != ele[21][21];
    ele[6][21] != ele[22][21];
    ele[6][21] != ele[23][21];
    ele[6][21] != ele[24][21];
    ele[6][21] != ele[6][22];
    ele[6][21] != ele[6][23];
    ele[6][21] != ele[6][24];
    ele[6][21] != ele[7][20];
    ele[6][21] != ele[7][21];
    ele[6][21] != ele[7][22];
    ele[6][21] != ele[7][23];
    ele[6][21] != ele[7][24];
    ele[6][21] != ele[8][20];
    ele[6][21] != ele[8][21];
    ele[6][21] != ele[8][22];
    ele[6][21] != ele[8][23];
    ele[6][21] != ele[8][24];
    ele[6][21] != ele[9][20];
    ele[6][21] != ele[9][21];
    ele[6][21] != ele[9][22];
    ele[6][21] != ele[9][23];
    ele[6][21] != ele[9][24];
    ele[6][22] != ele[10][22];
    ele[6][22] != ele[11][22];
    ele[6][22] != ele[12][22];
    ele[6][22] != ele[13][22];
    ele[6][22] != ele[14][22];
    ele[6][22] != ele[15][22];
    ele[6][22] != ele[16][22];
    ele[6][22] != ele[17][22];
    ele[6][22] != ele[18][22];
    ele[6][22] != ele[19][22];
    ele[6][22] != ele[20][22];
    ele[6][22] != ele[21][22];
    ele[6][22] != ele[22][22];
    ele[6][22] != ele[23][22];
    ele[6][22] != ele[24][22];
    ele[6][22] != ele[6][23];
    ele[6][22] != ele[6][24];
    ele[6][22] != ele[7][20];
    ele[6][22] != ele[7][21];
    ele[6][22] != ele[7][22];
    ele[6][22] != ele[7][23];
    ele[6][22] != ele[7][24];
    ele[6][22] != ele[8][20];
    ele[6][22] != ele[8][21];
    ele[6][22] != ele[8][22];
    ele[6][22] != ele[8][23];
    ele[6][22] != ele[8][24];
    ele[6][22] != ele[9][20];
    ele[6][22] != ele[9][21];
    ele[6][22] != ele[9][22];
    ele[6][22] != ele[9][23];
    ele[6][22] != ele[9][24];
    ele[6][23] != ele[10][23];
    ele[6][23] != ele[11][23];
    ele[6][23] != ele[12][23];
    ele[6][23] != ele[13][23];
    ele[6][23] != ele[14][23];
    ele[6][23] != ele[15][23];
    ele[6][23] != ele[16][23];
    ele[6][23] != ele[17][23];
    ele[6][23] != ele[18][23];
    ele[6][23] != ele[19][23];
    ele[6][23] != ele[20][23];
    ele[6][23] != ele[21][23];
    ele[6][23] != ele[22][23];
    ele[6][23] != ele[23][23];
    ele[6][23] != ele[24][23];
    ele[6][23] != ele[6][24];
    ele[6][23] != ele[7][20];
    ele[6][23] != ele[7][21];
    ele[6][23] != ele[7][22];
    ele[6][23] != ele[7][23];
    ele[6][23] != ele[7][24];
    ele[6][23] != ele[8][20];
    ele[6][23] != ele[8][21];
    ele[6][23] != ele[8][22];
    ele[6][23] != ele[8][23];
    ele[6][23] != ele[8][24];
    ele[6][23] != ele[9][20];
    ele[6][23] != ele[9][21];
    ele[6][23] != ele[9][22];
    ele[6][23] != ele[9][23];
    ele[6][23] != ele[9][24];
    ele[6][24] != ele[10][24];
    ele[6][24] != ele[11][24];
    ele[6][24] != ele[12][24];
    ele[6][24] != ele[13][24];
    ele[6][24] != ele[14][24];
    ele[6][24] != ele[15][24];
    ele[6][24] != ele[16][24];
    ele[6][24] != ele[17][24];
    ele[6][24] != ele[18][24];
    ele[6][24] != ele[19][24];
    ele[6][24] != ele[20][24];
    ele[6][24] != ele[21][24];
    ele[6][24] != ele[22][24];
    ele[6][24] != ele[23][24];
    ele[6][24] != ele[24][24];
    ele[6][24] != ele[7][20];
    ele[6][24] != ele[7][21];
    ele[6][24] != ele[7][22];
    ele[6][24] != ele[7][23];
    ele[6][24] != ele[7][24];
    ele[6][24] != ele[8][20];
    ele[6][24] != ele[8][21];
    ele[6][24] != ele[8][22];
    ele[6][24] != ele[8][23];
    ele[6][24] != ele[8][24];
    ele[6][24] != ele[9][20];
    ele[6][24] != ele[9][21];
    ele[6][24] != ele[9][22];
    ele[6][24] != ele[9][23];
    ele[6][24] != ele[9][24];
    ele[6][3] != ele[10][3];
    ele[6][3] != ele[11][3];
    ele[6][3] != ele[12][3];
    ele[6][3] != ele[13][3];
    ele[6][3] != ele[14][3];
    ele[6][3] != ele[15][3];
    ele[6][3] != ele[16][3];
    ele[6][3] != ele[17][3];
    ele[6][3] != ele[18][3];
    ele[6][3] != ele[19][3];
    ele[6][3] != ele[20][3];
    ele[6][3] != ele[21][3];
    ele[6][3] != ele[22][3];
    ele[6][3] != ele[23][3];
    ele[6][3] != ele[24][3];
    ele[6][3] != ele[6][10];
    ele[6][3] != ele[6][11];
    ele[6][3] != ele[6][12];
    ele[6][3] != ele[6][13];
    ele[6][3] != ele[6][14];
    ele[6][3] != ele[6][15];
    ele[6][3] != ele[6][16];
    ele[6][3] != ele[6][17];
    ele[6][3] != ele[6][18];
    ele[6][3] != ele[6][19];
    ele[6][3] != ele[6][20];
    ele[6][3] != ele[6][21];
    ele[6][3] != ele[6][22];
    ele[6][3] != ele[6][23];
    ele[6][3] != ele[6][24];
    ele[6][3] != ele[6][4];
    ele[6][3] != ele[6][5];
    ele[6][3] != ele[6][6];
    ele[6][3] != ele[6][7];
    ele[6][3] != ele[6][8];
    ele[6][3] != ele[6][9];
    ele[6][3] != ele[7][0];
    ele[6][3] != ele[7][1];
    ele[6][3] != ele[7][2];
    ele[6][3] != ele[7][3];
    ele[6][3] != ele[7][4];
    ele[6][3] != ele[8][0];
    ele[6][3] != ele[8][1];
    ele[6][3] != ele[8][2];
    ele[6][3] != ele[8][3];
    ele[6][3] != ele[8][4];
    ele[6][3] != ele[9][0];
    ele[6][3] != ele[9][1];
    ele[6][3] != ele[9][2];
    ele[6][3] != ele[9][3];
    ele[6][3] != ele[9][4];
    ele[6][4] != ele[10][4];
    ele[6][4] != ele[11][4];
    ele[6][4] != ele[12][4];
    ele[6][4] != ele[13][4];
    ele[6][4] != ele[14][4];
    ele[6][4] != ele[15][4];
    ele[6][4] != ele[16][4];
    ele[6][4] != ele[17][4];
    ele[6][4] != ele[18][4];
    ele[6][4] != ele[19][4];
    ele[6][4] != ele[20][4];
    ele[6][4] != ele[21][4];
    ele[6][4] != ele[22][4];
    ele[6][4] != ele[23][4];
    ele[6][4] != ele[24][4];
    ele[6][4] != ele[6][10];
    ele[6][4] != ele[6][11];
    ele[6][4] != ele[6][12];
    ele[6][4] != ele[6][13];
    ele[6][4] != ele[6][14];
    ele[6][4] != ele[6][15];
    ele[6][4] != ele[6][16];
    ele[6][4] != ele[6][17];
    ele[6][4] != ele[6][18];
    ele[6][4] != ele[6][19];
    ele[6][4] != ele[6][20];
    ele[6][4] != ele[6][21];
    ele[6][4] != ele[6][22];
    ele[6][4] != ele[6][23];
    ele[6][4] != ele[6][24];
    ele[6][4] != ele[6][5];
    ele[6][4] != ele[6][6];
    ele[6][4] != ele[6][7];
    ele[6][4] != ele[6][8];
    ele[6][4] != ele[6][9];
    ele[6][4] != ele[7][0];
    ele[6][4] != ele[7][1];
    ele[6][4] != ele[7][2];
    ele[6][4] != ele[7][3];
    ele[6][4] != ele[7][4];
    ele[6][4] != ele[8][0];
    ele[6][4] != ele[8][1];
    ele[6][4] != ele[8][2];
    ele[6][4] != ele[8][3];
    ele[6][4] != ele[8][4];
    ele[6][4] != ele[9][0];
    ele[6][4] != ele[9][1];
    ele[6][4] != ele[9][2];
    ele[6][4] != ele[9][3];
    ele[6][4] != ele[9][4];
    ele[6][5] != ele[10][5];
    ele[6][5] != ele[11][5];
    ele[6][5] != ele[12][5];
    ele[6][5] != ele[13][5];
    ele[6][5] != ele[14][5];
    ele[6][5] != ele[15][5];
    ele[6][5] != ele[16][5];
    ele[6][5] != ele[17][5];
    ele[6][5] != ele[18][5];
    ele[6][5] != ele[19][5];
    ele[6][5] != ele[20][5];
    ele[6][5] != ele[21][5];
    ele[6][5] != ele[22][5];
    ele[6][5] != ele[23][5];
    ele[6][5] != ele[24][5];
    ele[6][5] != ele[6][10];
    ele[6][5] != ele[6][11];
    ele[6][5] != ele[6][12];
    ele[6][5] != ele[6][13];
    ele[6][5] != ele[6][14];
    ele[6][5] != ele[6][15];
    ele[6][5] != ele[6][16];
    ele[6][5] != ele[6][17];
    ele[6][5] != ele[6][18];
    ele[6][5] != ele[6][19];
    ele[6][5] != ele[6][20];
    ele[6][5] != ele[6][21];
    ele[6][5] != ele[6][22];
    ele[6][5] != ele[6][23];
    ele[6][5] != ele[6][24];
    ele[6][5] != ele[6][6];
    ele[6][5] != ele[6][7];
    ele[6][5] != ele[6][8];
    ele[6][5] != ele[6][9];
    ele[6][5] != ele[7][5];
    ele[6][5] != ele[7][6];
    ele[6][5] != ele[7][7];
    ele[6][5] != ele[7][8];
    ele[6][5] != ele[7][9];
    ele[6][5] != ele[8][5];
    ele[6][5] != ele[8][6];
    ele[6][5] != ele[8][7];
    ele[6][5] != ele[8][8];
    ele[6][5] != ele[8][9];
    ele[6][5] != ele[9][5];
    ele[6][5] != ele[9][6];
    ele[6][5] != ele[9][7];
    ele[6][5] != ele[9][8];
    ele[6][5] != ele[9][9];
    ele[6][6] != ele[10][6];
    ele[6][6] != ele[11][6];
    ele[6][6] != ele[12][6];
    ele[6][6] != ele[13][6];
    ele[6][6] != ele[14][6];
    ele[6][6] != ele[15][6];
    ele[6][6] != ele[16][6];
    ele[6][6] != ele[17][6];
    ele[6][6] != ele[18][6];
    ele[6][6] != ele[19][6];
    ele[6][6] != ele[20][6];
    ele[6][6] != ele[21][6];
    ele[6][6] != ele[22][6];
    ele[6][6] != ele[23][6];
    ele[6][6] != ele[24][6];
    ele[6][6] != ele[6][10];
    ele[6][6] != ele[6][11];
    ele[6][6] != ele[6][12];
    ele[6][6] != ele[6][13];
    ele[6][6] != ele[6][14];
    ele[6][6] != ele[6][15];
    ele[6][6] != ele[6][16];
    ele[6][6] != ele[6][17];
    ele[6][6] != ele[6][18];
    ele[6][6] != ele[6][19];
    ele[6][6] != ele[6][20];
    ele[6][6] != ele[6][21];
    ele[6][6] != ele[6][22];
    ele[6][6] != ele[6][23];
    ele[6][6] != ele[6][24];
    ele[6][6] != ele[6][7];
    ele[6][6] != ele[6][8];
    ele[6][6] != ele[6][9];
    ele[6][6] != ele[7][5];
    ele[6][6] != ele[7][6];
    ele[6][6] != ele[7][7];
    ele[6][6] != ele[7][8];
    ele[6][6] != ele[7][9];
    ele[6][6] != ele[8][5];
    ele[6][6] != ele[8][6];
    ele[6][6] != ele[8][7];
    ele[6][6] != ele[8][8];
    ele[6][6] != ele[8][9];
    ele[6][6] != ele[9][5];
    ele[6][6] != ele[9][6];
    ele[6][6] != ele[9][7];
    ele[6][6] != ele[9][8];
    ele[6][6] != ele[9][9];
    ele[6][7] != ele[10][7];
    ele[6][7] != ele[11][7];
    ele[6][7] != ele[12][7];
    ele[6][7] != ele[13][7];
    ele[6][7] != ele[14][7];
    ele[6][7] != ele[15][7];
    ele[6][7] != ele[16][7];
    ele[6][7] != ele[17][7];
    ele[6][7] != ele[18][7];
    ele[6][7] != ele[19][7];
    ele[6][7] != ele[20][7];
    ele[6][7] != ele[21][7];
    ele[6][7] != ele[22][7];
    ele[6][7] != ele[23][7];
    ele[6][7] != ele[24][7];
    ele[6][7] != ele[6][10];
    ele[6][7] != ele[6][11];
    ele[6][7] != ele[6][12];
    ele[6][7] != ele[6][13];
    ele[6][7] != ele[6][14];
    ele[6][7] != ele[6][15];
    ele[6][7] != ele[6][16];
    ele[6][7] != ele[6][17];
    ele[6][7] != ele[6][18];
    ele[6][7] != ele[6][19];
    ele[6][7] != ele[6][20];
    ele[6][7] != ele[6][21];
    ele[6][7] != ele[6][22];
    ele[6][7] != ele[6][23];
    ele[6][7] != ele[6][24];
    ele[6][7] != ele[6][8];
    ele[6][7] != ele[6][9];
    ele[6][7] != ele[7][5];
    ele[6][7] != ele[7][6];
    ele[6][7] != ele[7][7];
    ele[6][7] != ele[7][8];
    ele[6][7] != ele[7][9];
    ele[6][7] != ele[8][5];
    ele[6][7] != ele[8][6];
    ele[6][7] != ele[8][7];
    ele[6][7] != ele[8][8];
    ele[6][7] != ele[8][9];
    ele[6][7] != ele[9][5];
    ele[6][7] != ele[9][6];
    ele[6][7] != ele[9][7];
    ele[6][7] != ele[9][8];
    ele[6][7] != ele[9][9];
    ele[6][8] != ele[10][8];
    ele[6][8] != ele[11][8];
    ele[6][8] != ele[12][8];
    ele[6][8] != ele[13][8];
    ele[6][8] != ele[14][8];
    ele[6][8] != ele[15][8];
    ele[6][8] != ele[16][8];
    ele[6][8] != ele[17][8];
    ele[6][8] != ele[18][8];
    ele[6][8] != ele[19][8];
    ele[6][8] != ele[20][8];
    ele[6][8] != ele[21][8];
    ele[6][8] != ele[22][8];
    ele[6][8] != ele[23][8];
    ele[6][8] != ele[24][8];
    ele[6][8] != ele[6][10];
    ele[6][8] != ele[6][11];
    ele[6][8] != ele[6][12];
    ele[6][8] != ele[6][13];
    ele[6][8] != ele[6][14];
    ele[6][8] != ele[6][15];
    ele[6][8] != ele[6][16];
    ele[6][8] != ele[6][17];
    ele[6][8] != ele[6][18];
    ele[6][8] != ele[6][19];
    ele[6][8] != ele[6][20];
    ele[6][8] != ele[6][21];
    ele[6][8] != ele[6][22];
    ele[6][8] != ele[6][23];
    ele[6][8] != ele[6][24];
    ele[6][8] != ele[6][9];
    ele[6][8] != ele[7][5];
    ele[6][8] != ele[7][6];
    ele[6][8] != ele[7][7];
    ele[6][8] != ele[7][8];
    ele[6][8] != ele[7][9];
    ele[6][8] != ele[8][5];
    ele[6][8] != ele[8][6];
    ele[6][8] != ele[8][7];
    ele[6][8] != ele[8][8];
    ele[6][8] != ele[8][9];
    ele[6][8] != ele[9][5];
    ele[6][8] != ele[9][6];
    ele[6][8] != ele[9][7];
    ele[6][8] != ele[9][8];
    ele[6][8] != ele[9][9];
    ele[6][9] != ele[10][9];
    ele[6][9] != ele[11][9];
    ele[6][9] != ele[12][9];
    ele[6][9] != ele[13][9];
    ele[6][9] != ele[14][9];
    ele[6][9] != ele[15][9];
    ele[6][9] != ele[16][9];
    ele[6][9] != ele[17][9];
    ele[6][9] != ele[18][9];
    ele[6][9] != ele[19][9];
    ele[6][9] != ele[20][9];
    ele[6][9] != ele[21][9];
    ele[6][9] != ele[22][9];
    ele[6][9] != ele[23][9];
    ele[6][9] != ele[24][9];
    ele[6][9] != ele[6][10];
    ele[6][9] != ele[6][11];
    ele[6][9] != ele[6][12];
    ele[6][9] != ele[6][13];
    ele[6][9] != ele[6][14];
    ele[6][9] != ele[6][15];
    ele[6][9] != ele[6][16];
    ele[6][9] != ele[6][17];
    ele[6][9] != ele[6][18];
    ele[6][9] != ele[6][19];
    ele[6][9] != ele[6][20];
    ele[6][9] != ele[6][21];
    ele[6][9] != ele[6][22];
    ele[6][9] != ele[6][23];
    ele[6][9] != ele[6][24];
    ele[6][9] != ele[7][5];
    ele[6][9] != ele[7][6];
    ele[6][9] != ele[7][7];
    ele[6][9] != ele[7][8];
    ele[6][9] != ele[7][9];
    ele[6][9] != ele[8][5];
    ele[6][9] != ele[8][6];
    ele[6][9] != ele[8][7];
    ele[6][9] != ele[8][8];
    ele[6][9] != ele[8][9];
    ele[6][9] != ele[9][5];
    ele[6][9] != ele[9][6];
    ele[6][9] != ele[9][7];
    ele[6][9] != ele[9][8];
    ele[6][9] != ele[9][9];
    ele[7][0] != ele[10][0];
    ele[7][0] != ele[11][0];
    ele[7][0] != ele[12][0];
    ele[7][0] != ele[13][0];
    ele[7][0] != ele[14][0];
    ele[7][0] != ele[15][0];
    ele[7][0] != ele[16][0];
    ele[7][0] != ele[17][0];
    ele[7][0] != ele[18][0];
    ele[7][0] != ele[19][0];
    ele[7][0] != ele[20][0];
    ele[7][0] != ele[21][0];
    ele[7][0] != ele[22][0];
    ele[7][0] != ele[23][0];
    ele[7][0] != ele[24][0];
    ele[7][0] != ele[7][1];
    ele[7][0] != ele[7][10];
    ele[7][0] != ele[7][11];
    ele[7][0] != ele[7][12];
    ele[7][0] != ele[7][13];
    ele[7][0] != ele[7][14];
    ele[7][0] != ele[7][15];
    ele[7][0] != ele[7][16];
    ele[7][0] != ele[7][17];
    ele[7][0] != ele[7][18];
    ele[7][0] != ele[7][19];
    ele[7][0] != ele[7][2];
    ele[7][0] != ele[7][20];
    ele[7][0] != ele[7][21];
    ele[7][0] != ele[7][22];
    ele[7][0] != ele[7][23];
    ele[7][0] != ele[7][24];
    ele[7][0] != ele[7][3];
    ele[7][0] != ele[7][4];
    ele[7][0] != ele[7][5];
    ele[7][0] != ele[7][6];
    ele[7][0] != ele[7][7];
    ele[7][0] != ele[7][8];
    ele[7][0] != ele[7][9];
    ele[7][0] != ele[8][0];
    ele[7][0] != ele[8][1];
    ele[7][0] != ele[8][2];
    ele[7][0] != ele[8][3];
    ele[7][0] != ele[8][4];
    ele[7][0] != ele[9][0];
    ele[7][0] != ele[9][1];
    ele[7][0] != ele[9][2];
    ele[7][0] != ele[9][3];
    ele[7][0] != ele[9][4];
    ele[7][1] != ele[10][1];
    ele[7][1] != ele[11][1];
    ele[7][1] != ele[12][1];
    ele[7][1] != ele[13][1];
    ele[7][1] != ele[14][1];
    ele[7][1] != ele[15][1];
    ele[7][1] != ele[16][1];
    ele[7][1] != ele[17][1];
    ele[7][1] != ele[18][1];
    ele[7][1] != ele[19][1];
    ele[7][1] != ele[20][1];
    ele[7][1] != ele[21][1];
    ele[7][1] != ele[22][1];
    ele[7][1] != ele[23][1];
    ele[7][1] != ele[24][1];
    ele[7][1] != ele[7][10];
    ele[7][1] != ele[7][11];
    ele[7][1] != ele[7][12];
    ele[7][1] != ele[7][13];
    ele[7][1] != ele[7][14];
    ele[7][1] != ele[7][15];
    ele[7][1] != ele[7][16];
    ele[7][1] != ele[7][17];
    ele[7][1] != ele[7][18];
    ele[7][1] != ele[7][19];
    ele[7][1] != ele[7][2];
    ele[7][1] != ele[7][20];
    ele[7][1] != ele[7][21];
    ele[7][1] != ele[7][22];
    ele[7][1] != ele[7][23];
    ele[7][1] != ele[7][24];
    ele[7][1] != ele[7][3];
    ele[7][1] != ele[7][4];
    ele[7][1] != ele[7][5];
    ele[7][1] != ele[7][6];
    ele[7][1] != ele[7][7];
    ele[7][1] != ele[7][8];
    ele[7][1] != ele[7][9];
    ele[7][1] != ele[8][0];
    ele[7][1] != ele[8][1];
    ele[7][1] != ele[8][2];
    ele[7][1] != ele[8][3];
    ele[7][1] != ele[8][4];
    ele[7][1] != ele[9][0];
    ele[7][1] != ele[9][1];
    ele[7][1] != ele[9][2];
    ele[7][1] != ele[9][3];
    ele[7][1] != ele[9][4];
    ele[7][10] != ele[10][10];
    ele[7][10] != ele[11][10];
    ele[7][10] != ele[12][10];
    ele[7][10] != ele[13][10];
    ele[7][10] != ele[14][10];
    ele[7][10] != ele[15][10];
    ele[7][10] != ele[16][10];
    ele[7][10] != ele[17][10];
    ele[7][10] != ele[18][10];
    ele[7][10] != ele[19][10];
    ele[7][10] != ele[20][10];
    ele[7][10] != ele[21][10];
    ele[7][10] != ele[22][10];
    ele[7][10] != ele[23][10];
    ele[7][10] != ele[24][10];
    ele[7][10] != ele[7][11];
    ele[7][10] != ele[7][12];
    ele[7][10] != ele[7][13];
    ele[7][10] != ele[7][14];
    ele[7][10] != ele[7][15];
    ele[7][10] != ele[7][16];
    ele[7][10] != ele[7][17];
    ele[7][10] != ele[7][18];
    ele[7][10] != ele[7][19];
    ele[7][10] != ele[7][20];
    ele[7][10] != ele[7][21];
    ele[7][10] != ele[7][22];
    ele[7][10] != ele[7][23];
    ele[7][10] != ele[7][24];
    ele[7][10] != ele[8][10];
    ele[7][10] != ele[8][11];
    ele[7][10] != ele[8][12];
    ele[7][10] != ele[8][13];
    ele[7][10] != ele[8][14];
    ele[7][10] != ele[9][10];
    ele[7][10] != ele[9][11];
    ele[7][10] != ele[9][12];
    ele[7][10] != ele[9][13];
    ele[7][10] != ele[9][14];
    ele[7][11] != ele[10][11];
    ele[7][11] != ele[11][11];
    ele[7][11] != ele[12][11];
    ele[7][11] != ele[13][11];
    ele[7][11] != ele[14][11];
    ele[7][11] != ele[15][11];
    ele[7][11] != ele[16][11];
    ele[7][11] != ele[17][11];
    ele[7][11] != ele[18][11];
    ele[7][11] != ele[19][11];
    ele[7][11] != ele[20][11];
    ele[7][11] != ele[21][11];
    ele[7][11] != ele[22][11];
    ele[7][11] != ele[23][11];
    ele[7][11] != ele[24][11];
    ele[7][11] != ele[7][12];
    ele[7][11] != ele[7][13];
    ele[7][11] != ele[7][14];
    ele[7][11] != ele[7][15];
    ele[7][11] != ele[7][16];
    ele[7][11] != ele[7][17];
    ele[7][11] != ele[7][18];
    ele[7][11] != ele[7][19];
    ele[7][11] != ele[7][20];
    ele[7][11] != ele[7][21];
    ele[7][11] != ele[7][22];
    ele[7][11] != ele[7][23];
    ele[7][11] != ele[7][24];
    ele[7][11] != ele[8][10];
    ele[7][11] != ele[8][11];
    ele[7][11] != ele[8][12];
    ele[7][11] != ele[8][13];
    ele[7][11] != ele[8][14];
    ele[7][11] != ele[9][10];
    ele[7][11] != ele[9][11];
    ele[7][11] != ele[9][12];
    ele[7][11] != ele[9][13];
    ele[7][11] != ele[9][14];
    ele[7][12] != ele[10][12];
    ele[7][12] != ele[11][12];
    ele[7][12] != ele[12][12];
    ele[7][12] != ele[13][12];
    ele[7][12] != ele[14][12];
    ele[7][12] != ele[15][12];
    ele[7][12] != ele[16][12];
    ele[7][12] != ele[17][12];
    ele[7][12] != ele[18][12];
    ele[7][12] != ele[19][12];
    ele[7][12] != ele[20][12];
    ele[7][12] != ele[21][12];
    ele[7][12] != ele[22][12];
    ele[7][12] != ele[23][12];
    ele[7][12] != ele[24][12];
    ele[7][12] != ele[7][13];
    ele[7][12] != ele[7][14];
    ele[7][12] != ele[7][15];
    ele[7][12] != ele[7][16];
    ele[7][12] != ele[7][17];
    ele[7][12] != ele[7][18];
    ele[7][12] != ele[7][19];
    ele[7][12] != ele[7][20];
    ele[7][12] != ele[7][21];
    ele[7][12] != ele[7][22];
    ele[7][12] != ele[7][23];
    ele[7][12] != ele[7][24];
    ele[7][12] != ele[8][10];
    ele[7][12] != ele[8][11];
    ele[7][12] != ele[8][12];
    ele[7][12] != ele[8][13];
    ele[7][12] != ele[8][14];
    ele[7][12] != ele[9][10];
    ele[7][12] != ele[9][11];
    ele[7][12] != ele[9][12];
    ele[7][12] != ele[9][13];
    ele[7][12] != ele[9][14];
    ele[7][13] != ele[10][13];
    ele[7][13] != ele[11][13];
    ele[7][13] != ele[12][13];
    ele[7][13] != ele[13][13];
    ele[7][13] != ele[14][13];
    ele[7][13] != ele[15][13];
    ele[7][13] != ele[16][13];
    ele[7][13] != ele[17][13];
    ele[7][13] != ele[18][13];
    ele[7][13] != ele[19][13];
    ele[7][13] != ele[20][13];
    ele[7][13] != ele[21][13];
    ele[7][13] != ele[22][13];
    ele[7][13] != ele[23][13];
    ele[7][13] != ele[24][13];
    ele[7][13] != ele[7][14];
    ele[7][13] != ele[7][15];
    ele[7][13] != ele[7][16];
    ele[7][13] != ele[7][17];
    ele[7][13] != ele[7][18];
    ele[7][13] != ele[7][19];
    ele[7][13] != ele[7][20];
    ele[7][13] != ele[7][21];
    ele[7][13] != ele[7][22];
    ele[7][13] != ele[7][23];
    ele[7][13] != ele[7][24];
    ele[7][13] != ele[8][10];
    ele[7][13] != ele[8][11];
    ele[7][13] != ele[8][12];
    ele[7][13] != ele[8][13];
    ele[7][13] != ele[8][14];
    ele[7][13] != ele[9][10];
    ele[7][13] != ele[9][11];
    ele[7][13] != ele[9][12];
    ele[7][13] != ele[9][13];
    ele[7][13] != ele[9][14];
    ele[7][14] != ele[10][14];
    ele[7][14] != ele[11][14];
    ele[7][14] != ele[12][14];
    ele[7][14] != ele[13][14];
    ele[7][14] != ele[14][14];
    ele[7][14] != ele[15][14];
    ele[7][14] != ele[16][14];
    ele[7][14] != ele[17][14];
    ele[7][14] != ele[18][14];
    ele[7][14] != ele[19][14];
    ele[7][14] != ele[20][14];
    ele[7][14] != ele[21][14];
    ele[7][14] != ele[22][14];
    ele[7][14] != ele[23][14];
    ele[7][14] != ele[24][14];
    ele[7][14] != ele[7][15];
    ele[7][14] != ele[7][16];
    ele[7][14] != ele[7][17];
    ele[7][14] != ele[7][18];
    ele[7][14] != ele[7][19];
    ele[7][14] != ele[7][20];
    ele[7][14] != ele[7][21];
    ele[7][14] != ele[7][22];
    ele[7][14] != ele[7][23];
    ele[7][14] != ele[7][24];
    ele[7][14] != ele[8][10];
    ele[7][14] != ele[8][11];
    ele[7][14] != ele[8][12];
    ele[7][14] != ele[8][13];
    ele[7][14] != ele[8][14];
    ele[7][14] != ele[9][10];
    ele[7][14] != ele[9][11];
    ele[7][14] != ele[9][12];
    ele[7][14] != ele[9][13];
    ele[7][14] != ele[9][14];
    ele[7][15] != ele[10][15];
    ele[7][15] != ele[11][15];
    ele[7][15] != ele[12][15];
    ele[7][15] != ele[13][15];
    ele[7][15] != ele[14][15];
    ele[7][15] != ele[15][15];
    ele[7][15] != ele[16][15];
    ele[7][15] != ele[17][15];
    ele[7][15] != ele[18][15];
    ele[7][15] != ele[19][15];
    ele[7][15] != ele[20][15];
    ele[7][15] != ele[21][15];
    ele[7][15] != ele[22][15];
    ele[7][15] != ele[23][15];
    ele[7][15] != ele[24][15];
    ele[7][15] != ele[7][16];
    ele[7][15] != ele[7][17];
    ele[7][15] != ele[7][18];
    ele[7][15] != ele[7][19];
    ele[7][15] != ele[7][20];
    ele[7][15] != ele[7][21];
    ele[7][15] != ele[7][22];
    ele[7][15] != ele[7][23];
    ele[7][15] != ele[7][24];
    ele[7][15] != ele[8][15];
    ele[7][15] != ele[8][16];
    ele[7][15] != ele[8][17];
    ele[7][15] != ele[8][18];
    ele[7][15] != ele[8][19];
    ele[7][15] != ele[9][15];
    ele[7][15] != ele[9][16];
    ele[7][15] != ele[9][17];
    ele[7][15] != ele[9][18];
    ele[7][15] != ele[9][19];
    ele[7][16] != ele[10][16];
    ele[7][16] != ele[11][16];
    ele[7][16] != ele[12][16];
    ele[7][16] != ele[13][16];
    ele[7][16] != ele[14][16];
    ele[7][16] != ele[15][16];
    ele[7][16] != ele[16][16];
    ele[7][16] != ele[17][16];
    ele[7][16] != ele[18][16];
    ele[7][16] != ele[19][16];
    ele[7][16] != ele[20][16];
    ele[7][16] != ele[21][16];
    ele[7][16] != ele[22][16];
    ele[7][16] != ele[23][16];
    ele[7][16] != ele[24][16];
    ele[7][16] != ele[7][17];
    ele[7][16] != ele[7][18];
    ele[7][16] != ele[7][19];
    ele[7][16] != ele[7][20];
    ele[7][16] != ele[7][21];
    ele[7][16] != ele[7][22];
    ele[7][16] != ele[7][23];
    ele[7][16] != ele[7][24];
    ele[7][16] != ele[8][15];
    ele[7][16] != ele[8][16];
    ele[7][16] != ele[8][17];
    ele[7][16] != ele[8][18];
    ele[7][16] != ele[8][19];
    ele[7][16] != ele[9][15];
    ele[7][16] != ele[9][16];
    ele[7][16] != ele[9][17];
    ele[7][16] != ele[9][18];
    ele[7][16] != ele[9][19];
    ele[7][17] != ele[10][17];
    ele[7][17] != ele[11][17];
    ele[7][17] != ele[12][17];
    ele[7][17] != ele[13][17];
    ele[7][17] != ele[14][17];
    ele[7][17] != ele[15][17];
    ele[7][17] != ele[16][17];
    ele[7][17] != ele[17][17];
    ele[7][17] != ele[18][17];
    ele[7][17] != ele[19][17];
    ele[7][17] != ele[20][17];
    ele[7][17] != ele[21][17];
    ele[7][17] != ele[22][17];
    ele[7][17] != ele[23][17];
    ele[7][17] != ele[24][17];
    ele[7][17] != ele[7][18];
    ele[7][17] != ele[7][19];
    ele[7][17] != ele[7][20];
    ele[7][17] != ele[7][21];
    ele[7][17] != ele[7][22];
    ele[7][17] != ele[7][23];
    ele[7][17] != ele[7][24];
    ele[7][17] != ele[8][15];
    ele[7][17] != ele[8][16];
    ele[7][17] != ele[8][17];
    ele[7][17] != ele[8][18];
    ele[7][17] != ele[8][19];
    ele[7][17] != ele[9][15];
    ele[7][17] != ele[9][16];
    ele[7][17] != ele[9][17];
    ele[7][17] != ele[9][18];
    ele[7][17] != ele[9][19];
    ele[7][18] != ele[10][18];
    ele[7][18] != ele[11][18];
    ele[7][18] != ele[12][18];
    ele[7][18] != ele[13][18];
    ele[7][18] != ele[14][18];
    ele[7][18] != ele[15][18];
    ele[7][18] != ele[16][18];
    ele[7][18] != ele[17][18];
    ele[7][18] != ele[18][18];
    ele[7][18] != ele[19][18];
    ele[7][18] != ele[20][18];
    ele[7][18] != ele[21][18];
    ele[7][18] != ele[22][18];
    ele[7][18] != ele[23][18];
    ele[7][18] != ele[24][18];
    ele[7][18] != ele[7][19];
    ele[7][18] != ele[7][20];
    ele[7][18] != ele[7][21];
    ele[7][18] != ele[7][22];
    ele[7][18] != ele[7][23];
    ele[7][18] != ele[7][24];
    ele[7][18] != ele[8][15];
    ele[7][18] != ele[8][16];
    ele[7][18] != ele[8][17];
    ele[7][18] != ele[8][18];
    ele[7][18] != ele[8][19];
    ele[7][18] != ele[9][15];
    ele[7][18] != ele[9][16];
    ele[7][18] != ele[9][17];
    ele[7][18] != ele[9][18];
    ele[7][18] != ele[9][19];
    ele[7][19] != ele[10][19];
    ele[7][19] != ele[11][19];
    ele[7][19] != ele[12][19];
    ele[7][19] != ele[13][19];
    ele[7][19] != ele[14][19];
    ele[7][19] != ele[15][19];
    ele[7][19] != ele[16][19];
    ele[7][19] != ele[17][19];
    ele[7][19] != ele[18][19];
    ele[7][19] != ele[19][19];
    ele[7][19] != ele[20][19];
    ele[7][19] != ele[21][19];
    ele[7][19] != ele[22][19];
    ele[7][19] != ele[23][19];
    ele[7][19] != ele[24][19];
    ele[7][19] != ele[7][20];
    ele[7][19] != ele[7][21];
    ele[7][19] != ele[7][22];
    ele[7][19] != ele[7][23];
    ele[7][19] != ele[7][24];
    ele[7][19] != ele[8][15];
    ele[7][19] != ele[8][16];
    ele[7][19] != ele[8][17];
    ele[7][19] != ele[8][18];
    ele[7][19] != ele[8][19];
    ele[7][19] != ele[9][15];
    ele[7][19] != ele[9][16];
    ele[7][19] != ele[9][17];
    ele[7][19] != ele[9][18];
    ele[7][19] != ele[9][19];
    ele[7][2] != ele[10][2];
    ele[7][2] != ele[11][2];
    ele[7][2] != ele[12][2];
    ele[7][2] != ele[13][2];
    ele[7][2] != ele[14][2];
    ele[7][2] != ele[15][2];
    ele[7][2] != ele[16][2];
    ele[7][2] != ele[17][2];
    ele[7][2] != ele[18][2];
    ele[7][2] != ele[19][2];
    ele[7][2] != ele[20][2];
    ele[7][2] != ele[21][2];
    ele[7][2] != ele[22][2];
    ele[7][2] != ele[23][2];
    ele[7][2] != ele[24][2];
    ele[7][2] != ele[7][10];
    ele[7][2] != ele[7][11];
    ele[7][2] != ele[7][12];
    ele[7][2] != ele[7][13];
    ele[7][2] != ele[7][14];
    ele[7][2] != ele[7][15];
    ele[7][2] != ele[7][16];
    ele[7][2] != ele[7][17];
    ele[7][2] != ele[7][18];
    ele[7][2] != ele[7][19];
    ele[7][2] != ele[7][20];
    ele[7][2] != ele[7][21];
    ele[7][2] != ele[7][22];
    ele[7][2] != ele[7][23];
    ele[7][2] != ele[7][24];
    ele[7][2] != ele[7][3];
    ele[7][2] != ele[7][4];
    ele[7][2] != ele[7][5];
    ele[7][2] != ele[7][6];
    ele[7][2] != ele[7][7];
    ele[7][2] != ele[7][8];
    ele[7][2] != ele[7][9];
    ele[7][2] != ele[8][0];
    ele[7][2] != ele[8][1];
    ele[7][2] != ele[8][2];
    ele[7][2] != ele[8][3];
    ele[7][2] != ele[8][4];
    ele[7][2] != ele[9][0];
    ele[7][2] != ele[9][1];
    ele[7][2] != ele[9][2];
    ele[7][2] != ele[9][3];
    ele[7][2] != ele[9][4];
    ele[7][20] != ele[10][20];
    ele[7][20] != ele[11][20];
    ele[7][20] != ele[12][20];
    ele[7][20] != ele[13][20];
    ele[7][20] != ele[14][20];
    ele[7][20] != ele[15][20];
    ele[7][20] != ele[16][20];
    ele[7][20] != ele[17][20];
    ele[7][20] != ele[18][20];
    ele[7][20] != ele[19][20];
    ele[7][20] != ele[20][20];
    ele[7][20] != ele[21][20];
    ele[7][20] != ele[22][20];
    ele[7][20] != ele[23][20];
    ele[7][20] != ele[24][20];
    ele[7][20] != ele[7][21];
    ele[7][20] != ele[7][22];
    ele[7][20] != ele[7][23];
    ele[7][20] != ele[7][24];
    ele[7][20] != ele[8][20];
    ele[7][20] != ele[8][21];
    ele[7][20] != ele[8][22];
    ele[7][20] != ele[8][23];
    ele[7][20] != ele[8][24];
    ele[7][20] != ele[9][20];
    ele[7][20] != ele[9][21];
    ele[7][20] != ele[9][22];
    ele[7][20] != ele[9][23];
    ele[7][20] != ele[9][24];
    ele[7][21] != ele[10][21];
    ele[7][21] != ele[11][21];
    ele[7][21] != ele[12][21];
    ele[7][21] != ele[13][21];
    ele[7][21] != ele[14][21];
    ele[7][21] != ele[15][21];
    ele[7][21] != ele[16][21];
    ele[7][21] != ele[17][21];
    ele[7][21] != ele[18][21];
    ele[7][21] != ele[19][21];
    ele[7][21] != ele[20][21];
    ele[7][21] != ele[21][21];
    ele[7][21] != ele[22][21];
    ele[7][21] != ele[23][21];
    ele[7][21] != ele[24][21];
    ele[7][21] != ele[7][22];
    ele[7][21] != ele[7][23];
    ele[7][21] != ele[7][24];
    ele[7][21] != ele[8][20];
    ele[7][21] != ele[8][21];
    ele[7][21] != ele[8][22];
    ele[7][21] != ele[8][23];
    ele[7][21] != ele[8][24];
    ele[7][21] != ele[9][20];
    ele[7][21] != ele[9][21];
    ele[7][21] != ele[9][22];
    ele[7][21] != ele[9][23];
    ele[7][21] != ele[9][24];
    ele[7][22] != ele[10][22];
    ele[7][22] != ele[11][22];
    ele[7][22] != ele[12][22];
    ele[7][22] != ele[13][22];
    ele[7][22] != ele[14][22];
    ele[7][22] != ele[15][22];
    ele[7][22] != ele[16][22];
    ele[7][22] != ele[17][22];
    ele[7][22] != ele[18][22];
    ele[7][22] != ele[19][22];
    ele[7][22] != ele[20][22];
    ele[7][22] != ele[21][22];
    ele[7][22] != ele[22][22];
    ele[7][22] != ele[23][22];
    ele[7][22] != ele[24][22];
    ele[7][22] != ele[7][23];
    ele[7][22] != ele[7][24];
    ele[7][22] != ele[8][20];
    ele[7][22] != ele[8][21];
    ele[7][22] != ele[8][22];
    ele[7][22] != ele[8][23];
    ele[7][22] != ele[8][24];
    ele[7][22] != ele[9][20];
    ele[7][22] != ele[9][21];
    ele[7][22] != ele[9][22];
    ele[7][22] != ele[9][23];
    ele[7][22] != ele[9][24];
    ele[7][23] != ele[10][23];
    ele[7][23] != ele[11][23];
    ele[7][23] != ele[12][23];
    ele[7][23] != ele[13][23];
    ele[7][23] != ele[14][23];
    ele[7][23] != ele[15][23];
    ele[7][23] != ele[16][23];
    ele[7][23] != ele[17][23];
    ele[7][23] != ele[18][23];
    ele[7][23] != ele[19][23];
    ele[7][23] != ele[20][23];
    ele[7][23] != ele[21][23];
    ele[7][23] != ele[22][23];
    ele[7][23] != ele[23][23];
    ele[7][23] != ele[24][23];
    ele[7][23] != ele[7][24];
    ele[7][23] != ele[8][20];
    ele[7][23] != ele[8][21];
    ele[7][23] != ele[8][22];
    ele[7][23] != ele[8][23];
    ele[7][23] != ele[8][24];
    ele[7][23] != ele[9][20];
    ele[7][23] != ele[9][21];
    ele[7][23] != ele[9][22];
    ele[7][23] != ele[9][23];
    ele[7][23] != ele[9][24];
    ele[7][24] != ele[10][24];
    ele[7][24] != ele[11][24];
    ele[7][24] != ele[12][24];
    ele[7][24] != ele[13][24];
    ele[7][24] != ele[14][24];
    ele[7][24] != ele[15][24];
    ele[7][24] != ele[16][24];
    ele[7][24] != ele[17][24];
    ele[7][24] != ele[18][24];
    ele[7][24] != ele[19][24];
    ele[7][24] != ele[20][24];
    ele[7][24] != ele[21][24];
    ele[7][24] != ele[22][24];
    ele[7][24] != ele[23][24];
    ele[7][24] != ele[24][24];
    ele[7][24] != ele[8][20];
    ele[7][24] != ele[8][21];
    ele[7][24] != ele[8][22];
    ele[7][24] != ele[8][23];
    ele[7][24] != ele[8][24];
    ele[7][24] != ele[9][20];
    ele[7][24] != ele[9][21];
    ele[7][24] != ele[9][22];
    ele[7][24] != ele[9][23];
    ele[7][24] != ele[9][24];
    ele[7][3] != ele[10][3];
    ele[7][3] != ele[11][3];
    ele[7][3] != ele[12][3];
    ele[7][3] != ele[13][3];
    ele[7][3] != ele[14][3];
    ele[7][3] != ele[15][3];
    ele[7][3] != ele[16][3];
    ele[7][3] != ele[17][3];
    ele[7][3] != ele[18][3];
    ele[7][3] != ele[19][3];
    ele[7][3] != ele[20][3];
    ele[7][3] != ele[21][3];
    ele[7][3] != ele[22][3];
    ele[7][3] != ele[23][3];
    ele[7][3] != ele[24][3];
    ele[7][3] != ele[7][10];
    ele[7][3] != ele[7][11];
    ele[7][3] != ele[7][12];
    ele[7][3] != ele[7][13];
    ele[7][3] != ele[7][14];
    ele[7][3] != ele[7][15];
    ele[7][3] != ele[7][16];
    ele[7][3] != ele[7][17];
    ele[7][3] != ele[7][18];
    ele[7][3] != ele[7][19];
    ele[7][3] != ele[7][20];
    ele[7][3] != ele[7][21];
    ele[7][3] != ele[7][22];
    ele[7][3] != ele[7][23];
    ele[7][3] != ele[7][24];
    ele[7][3] != ele[7][4];
    ele[7][3] != ele[7][5];
    ele[7][3] != ele[7][6];
    ele[7][3] != ele[7][7];
    ele[7][3] != ele[7][8];
    ele[7][3] != ele[7][9];
    ele[7][3] != ele[8][0];
    ele[7][3] != ele[8][1];
    ele[7][3] != ele[8][2];
    ele[7][3] != ele[8][3];
    ele[7][3] != ele[8][4];
    ele[7][3] != ele[9][0];
    ele[7][3] != ele[9][1];
    ele[7][3] != ele[9][2];
    ele[7][3] != ele[9][3];
    ele[7][3] != ele[9][4];
    ele[7][4] != ele[10][4];
    ele[7][4] != ele[11][4];
    ele[7][4] != ele[12][4];
    ele[7][4] != ele[13][4];
    ele[7][4] != ele[14][4];
    ele[7][4] != ele[15][4];
    ele[7][4] != ele[16][4];
    ele[7][4] != ele[17][4];
    ele[7][4] != ele[18][4];
    ele[7][4] != ele[19][4];
    ele[7][4] != ele[20][4];
    ele[7][4] != ele[21][4];
    ele[7][4] != ele[22][4];
    ele[7][4] != ele[23][4];
    ele[7][4] != ele[24][4];
    ele[7][4] != ele[7][10];
    ele[7][4] != ele[7][11];
    ele[7][4] != ele[7][12];
    ele[7][4] != ele[7][13];
    ele[7][4] != ele[7][14];
    ele[7][4] != ele[7][15];
    ele[7][4] != ele[7][16];
    ele[7][4] != ele[7][17];
    ele[7][4] != ele[7][18];
    ele[7][4] != ele[7][19];
    ele[7][4] != ele[7][20];
    ele[7][4] != ele[7][21];
    ele[7][4] != ele[7][22];
    ele[7][4] != ele[7][23];
    ele[7][4] != ele[7][24];
    ele[7][4] != ele[7][5];
    ele[7][4] != ele[7][6];
    ele[7][4] != ele[7][7];
    ele[7][4] != ele[7][8];
    ele[7][4] != ele[7][9];
    ele[7][4] != ele[8][0];
    ele[7][4] != ele[8][1];
    ele[7][4] != ele[8][2];
    ele[7][4] != ele[8][3];
    ele[7][4] != ele[8][4];
    ele[7][4] != ele[9][0];
    ele[7][4] != ele[9][1];
    ele[7][4] != ele[9][2];
    ele[7][4] != ele[9][3];
    ele[7][4] != ele[9][4];
    ele[7][5] != ele[10][5];
    ele[7][5] != ele[11][5];
    ele[7][5] != ele[12][5];
    ele[7][5] != ele[13][5];
    ele[7][5] != ele[14][5];
    ele[7][5] != ele[15][5];
    ele[7][5] != ele[16][5];
    ele[7][5] != ele[17][5];
    ele[7][5] != ele[18][5];
    ele[7][5] != ele[19][5];
    ele[7][5] != ele[20][5];
    ele[7][5] != ele[21][5];
    ele[7][5] != ele[22][5];
    ele[7][5] != ele[23][5];
    ele[7][5] != ele[24][5];
    ele[7][5] != ele[7][10];
    ele[7][5] != ele[7][11];
    ele[7][5] != ele[7][12];
    ele[7][5] != ele[7][13];
    ele[7][5] != ele[7][14];
    ele[7][5] != ele[7][15];
    ele[7][5] != ele[7][16];
    ele[7][5] != ele[7][17];
    ele[7][5] != ele[7][18];
    ele[7][5] != ele[7][19];
    ele[7][5] != ele[7][20];
    ele[7][5] != ele[7][21];
    ele[7][5] != ele[7][22];
    ele[7][5] != ele[7][23];
    ele[7][5] != ele[7][24];
    ele[7][5] != ele[7][6];
    ele[7][5] != ele[7][7];
    ele[7][5] != ele[7][8];
    ele[7][5] != ele[7][9];
    ele[7][5] != ele[8][5];
    ele[7][5] != ele[8][6];
    ele[7][5] != ele[8][7];
    ele[7][5] != ele[8][8];
    ele[7][5] != ele[8][9];
    ele[7][5] != ele[9][5];
    ele[7][5] != ele[9][6];
    ele[7][5] != ele[9][7];
    ele[7][5] != ele[9][8];
    ele[7][5] != ele[9][9];
    ele[7][6] != ele[10][6];
    ele[7][6] != ele[11][6];
    ele[7][6] != ele[12][6];
    ele[7][6] != ele[13][6];
    ele[7][6] != ele[14][6];
    ele[7][6] != ele[15][6];
    ele[7][6] != ele[16][6];
    ele[7][6] != ele[17][6];
    ele[7][6] != ele[18][6];
    ele[7][6] != ele[19][6];
    ele[7][6] != ele[20][6];
    ele[7][6] != ele[21][6];
    ele[7][6] != ele[22][6];
    ele[7][6] != ele[23][6];
    ele[7][6] != ele[24][6];
    ele[7][6] != ele[7][10];
    ele[7][6] != ele[7][11];
    ele[7][6] != ele[7][12];
    ele[7][6] != ele[7][13];
    ele[7][6] != ele[7][14];
    ele[7][6] != ele[7][15];
    ele[7][6] != ele[7][16];
    ele[7][6] != ele[7][17];
    ele[7][6] != ele[7][18];
    ele[7][6] != ele[7][19];
    ele[7][6] != ele[7][20];
    ele[7][6] != ele[7][21];
    ele[7][6] != ele[7][22];
    ele[7][6] != ele[7][23];
    ele[7][6] != ele[7][24];
    ele[7][6] != ele[7][7];
    ele[7][6] != ele[7][8];
    ele[7][6] != ele[7][9];
    ele[7][6] != ele[8][5];
    ele[7][6] != ele[8][6];
    ele[7][6] != ele[8][7];
    ele[7][6] != ele[8][8];
    ele[7][6] != ele[8][9];
    ele[7][6] != ele[9][5];
    ele[7][6] != ele[9][6];
    ele[7][6] != ele[9][7];
    ele[7][6] != ele[9][8];
    ele[7][6] != ele[9][9];
    ele[7][7] != ele[10][7];
    ele[7][7] != ele[11][7];
    ele[7][7] != ele[12][7];
    ele[7][7] != ele[13][7];
    ele[7][7] != ele[14][7];
    ele[7][7] != ele[15][7];
    ele[7][7] != ele[16][7];
    ele[7][7] != ele[17][7];
    ele[7][7] != ele[18][7];
    ele[7][7] != ele[19][7];
    ele[7][7] != ele[20][7];
    ele[7][7] != ele[21][7];
    ele[7][7] != ele[22][7];
    ele[7][7] != ele[23][7];
    ele[7][7] != ele[24][7];
    ele[7][7] != ele[7][10];
    ele[7][7] != ele[7][11];
    ele[7][7] != ele[7][12];
    ele[7][7] != ele[7][13];
    ele[7][7] != ele[7][14];
    ele[7][7] != ele[7][15];
    ele[7][7] != ele[7][16];
    ele[7][7] != ele[7][17];
    ele[7][7] != ele[7][18];
    ele[7][7] != ele[7][19];
    ele[7][7] != ele[7][20];
    ele[7][7] != ele[7][21];
    ele[7][7] != ele[7][22];
    ele[7][7] != ele[7][23];
    ele[7][7] != ele[7][24];
    ele[7][7] != ele[7][8];
    ele[7][7] != ele[7][9];
    ele[7][7] != ele[8][5];
    ele[7][7] != ele[8][6];
    ele[7][7] != ele[8][7];
    ele[7][7] != ele[8][8];
    ele[7][7] != ele[8][9];
    ele[7][7] != ele[9][5];
    ele[7][7] != ele[9][6];
    ele[7][7] != ele[9][7];
    ele[7][7] != ele[9][8];
    ele[7][7] != ele[9][9];
    ele[7][8] != ele[10][8];
    ele[7][8] != ele[11][8];
    ele[7][8] != ele[12][8];
    ele[7][8] != ele[13][8];
    ele[7][8] != ele[14][8];
    ele[7][8] != ele[15][8];
    ele[7][8] != ele[16][8];
    ele[7][8] != ele[17][8];
    ele[7][8] != ele[18][8];
    ele[7][8] != ele[19][8];
    ele[7][8] != ele[20][8];
    ele[7][8] != ele[21][8];
    ele[7][8] != ele[22][8];
    ele[7][8] != ele[23][8];
    ele[7][8] != ele[24][8];
    ele[7][8] != ele[7][10];
    ele[7][8] != ele[7][11];
    ele[7][8] != ele[7][12];
    ele[7][8] != ele[7][13];
    ele[7][8] != ele[7][14];
    ele[7][8] != ele[7][15];
    ele[7][8] != ele[7][16];
    ele[7][8] != ele[7][17];
    ele[7][8] != ele[7][18];
    ele[7][8] != ele[7][19];
    ele[7][8] != ele[7][20];
    ele[7][8] != ele[7][21];
    ele[7][8] != ele[7][22];
    ele[7][8] != ele[7][23];
    ele[7][8] != ele[7][24];
    ele[7][8] != ele[7][9];
    ele[7][8] != ele[8][5];
    ele[7][8] != ele[8][6];
    ele[7][8] != ele[8][7];
    ele[7][8] != ele[8][8];
    ele[7][8] != ele[8][9];
    ele[7][8] != ele[9][5];
    ele[7][8] != ele[9][6];
    ele[7][8] != ele[9][7];
    ele[7][8] != ele[9][8];
    ele[7][8] != ele[9][9];
    ele[7][9] != ele[10][9];
    ele[7][9] != ele[11][9];
    ele[7][9] != ele[12][9];
    ele[7][9] != ele[13][9];
    ele[7][9] != ele[14][9];
    ele[7][9] != ele[15][9];
    ele[7][9] != ele[16][9];
    ele[7][9] != ele[17][9];
    ele[7][9] != ele[18][9];
    ele[7][9] != ele[19][9];
    ele[7][9] != ele[20][9];
    ele[7][9] != ele[21][9];
    ele[7][9] != ele[22][9];
    ele[7][9] != ele[23][9];
    ele[7][9] != ele[24][9];
    ele[7][9] != ele[7][10];
    ele[7][9] != ele[7][11];
    ele[7][9] != ele[7][12];
    ele[7][9] != ele[7][13];
    ele[7][9] != ele[7][14];
    ele[7][9] != ele[7][15];
    ele[7][9] != ele[7][16];
    ele[7][9] != ele[7][17];
    ele[7][9] != ele[7][18];
    ele[7][9] != ele[7][19];
    ele[7][9] != ele[7][20];
    ele[7][9] != ele[7][21];
    ele[7][9] != ele[7][22];
    ele[7][9] != ele[7][23];
    ele[7][9] != ele[7][24];
    ele[7][9] != ele[8][5];
    ele[7][9] != ele[8][6];
    ele[7][9] != ele[8][7];
    ele[7][9] != ele[8][8];
    ele[7][9] != ele[8][9];
    ele[7][9] != ele[9][5];
    ele[7][9] != ele[9][6];
    ele[7][9] != ele[9][7];
    ele[7][9] != ele[9][8];
    ele[7][9] != ele[9][9];
    ele[8][0] != ele[10][0];
    ele[8][0] != ele[11][0];
    ele[8][0] != ele[12][0];
    ele[8][0] != ele[13][0];
    ele[8][0] != ele[14][0];
    ele[8][0] != ele[15][0];
    ele[8][0] != ele[16][0];
    ele[8][0] != ele[17][0];
    ele[8][0] != ele[18][0];
    ele[8][0] != ele[19][0];
    ele[8][0] != ele[20][0];
    ele[8][0] != ele[21][0];
    ele[8][0] != ele[22][0];
    ele[8][0] != ele[23][0];
    ele[8][0] != ele[24][0];
    ele[8][0] != ele[8][1];
    ele[8][0] != ele[8][10];
    ele[8][0] != ele[8][11];
    ele[8][0] != ele[8][12];
    ele[8][0] != ele[8][13];
    ele[8][0] != ele[8][14];
    ele[8][0] != ele[8][15];
    ele[8][0] != ele[8][16];
    ele[8][0] != ele[8][17];
    ele[8][0] != ele[8][18];
    ele[8][0] != ele[8][19];
    ele[8][0] != ele[8][2];
    ele[8][0] != ele[8][20];
    ele[8][0] != ele[8][21];
    ele[8][0] != ele[8][22];
    ele[8][0] != ele[8][23];
    ele[8][0] != ele[8][24];
    ele[8][0] != ele[8][3];
    ele[8][0] != ele[8][4];
    ele[8][0] != ele[8][5];
    ele[8][0] != ele[8][6];
    ele[8][0] != ele[8][7];
    ele[8][0] != ele[8][8];
    ele[8][0] != ele[8][9];
    ele[8][0] != ele[9][0];
    ele[8][0] != ele[9][1];
    ele[8][0] != ele[9][2];
    ele[8][0] != ele[9][3];
    ele[8][0] != ele[9][4];
    ele[8][1] != ele[10][1];
    ele[8][1] != ele[11][1];
    ele[8][1] != ele[12][1];
    ele[8][1] != ele[13][1];
    ele[8][1] != ele[14][1];
    ele[8][1] != ele[15][1];
    ele[8][1] != ele[16][1];
    ele[8][1] != ele[17][1];
    ele[8][1] != ele[18][1];
    ele[8][1] != ele[19][1];
    ele[8][1] != ele[20][1];
    ele[8][1] != ele[21][1];
    ele[8][1] != ele[22][1];
    ele[8][1] != ele[23][1];
    ele[8][1] != ele[24][1];
    ele[8][1] != ele[8][10];
    ele[8][1] != ele[8][11];
    ele[8][1] != ele[8][12];
    ele[8][1] != ele[8][13];
    ele[8][1] != ele[8][14];
    ele[8][1] != ele[8][15];
    ele[8][1] != ele[8][16];
    ele[8][1] != ele[8][17];
    ele[8][1] != ele[8][18];
    ele[8][1] != ele[8][19];
    ele[8][1] != ele[8][2];
    ele[8][1] != ele[8][20];
    ele[8][1] != ele[8][21];
    ele[8][1] != ele[8][22];
    ele[8][1] != ele[8][23];
    ele[8][1] != ele[8][24];
    ele[8][1] != ele[8][3];
    ele[8][1] != ele[8][4];
    ele[8][1] != ele[8][5];
    ele[8][1] != ele[8][6];
    ele[8][1] != ele[8][7];
    ele[8][1] != ele[8][8];
    ele[8][1] != ele[8][9];
    ele[8][1] != ele[9][0];
    ele[8][1] != ele[9][1];
    ele[8][1] != ele[9][2];
    ele[8][1] != ele[9][3];
    ele[8][1] != ele[9][4];
    ele[8][10] != ele[10][10];
    ele[8][10] != ele[11][10];
    ele[8][10] != ele[12][10];
    ele[8][10] != ele[13][10];
    ele[8][10] != ele[14][10];
    ele[8][10] != ele[15][10];
    ele[8][10] != ele[16][10];
    ele[8][10] != ele[17][10];
    ele[8][10] != ele[18][10];
    ele[8][10] != ele[19][10];
    ele[8][10] != ele[20][10];
    ele[8][10] != ele[21][10];
    ele[8][10] != ele[22][10];
    ele[8][10] != ele[23][10];
    ele[8][10] != ele[24][10];
    ele[8][10] != ele[8][11];
    ele[8][10] != ele[8][12];
    ele[8][10] != ele[8][13];
    ele[8][10] != ele[8][14];
    ele[8][10] != ele[8][15];
    ele[8][10] != ele[8][16];
    ele[8][10] != ele[8][17];
    ele[8][10] != ele[8][18];
    ele[8][10] != ele[8][19];
    ele[8][10] != ele[8][20];
    ele[8][10] != ele[8][21];
    ele[8][10] != ele[8][22];
    ele[8][10] != ele[8][23];
    ele[8][10] != ele[8][24];
    ele[8][10] != ele[9][10];
    ele[8][10] != ele[9][11];
    ele[8][10] != ele[9][12];
    ele[8][10] != ele[9][13];
    ele[8][10] != ele[9][14];
    ele[8][11] != ele[10][11];
    ele[8][11] != ele[11][11];
    ele[8][11] != ele[12][11];
    ele[8][11] != ele[13][11];
    ele[8][11] != ele[14][11];
    ele[8][11] != ele[15][11];
    ele[8][11] != ele[16][11];
    ele[8][11] != ele[17][11];
    ele[8][11] != ele[18][11];
    ele[8][11] != ele[19][11];
    ele[8][11] != ele[20][11];
    ele[8][11] != ele[21][11];
    ele[8][11] != ele[22][11];
    ele[8][11] != ele[23][11];
    ele[8][11] != ele[24][11];
    ele[8][11] != ele[8][12];
    ele[8][11] != ele[8][13];
    ele[8][11] != ele[8][14];
    ele[8][11] != ele[8][15];
    ele[8][11] != ele[8][16];
    ele[8][11] != ele[8][17];
    ele[8][11] != ele[8][18];
    ele[8][11] != ele[8][19];
    ele[8][11] != ele[8][20];
    ele[8][11] != ele[8][21];
    ele[8][11] != ele[8][22];
    ele[8][11] != ele[8][23];
    ele[8][11] != ele[8][24];
    ele[8][11] != ele[9][10];
    ele[8][11] != ele[9][11];
    ele[8][11] != ele[9][12];
    ele[8][11] != ele[9][13];
    ele[8][11] != ele[9][14];
    ele[8][12] != ele[10][12];
    ele[8][12] != ele[11][12];
    ele[8][12] != ele[12][12];
    ele[8][12] != ele[13][12];
    ele[8][12] != ele[14][12];
    ele[8][12] != ele[15][12];
    ele[8][12] != ele[16][12];
    ele[8][12] != ele[17][12];
    ele[8][12] != ele[18][12];
    ele[8][12] != ele[19][12];
    ele[8][12] != ele[20][12];
    ele[8][12] != ele[21][12];
    ele[8][12] != ele[22][12];
    ele[8][12] != ele[23][12];
    ele[8][12] != ele[24][12];
    ele[8][12] != ele[8][13];
    ele[8][12] != ele[8][14];
    ele[8][12] != ele[8][15];
    ele[8][12] != ele[8][16];
    ele[8][12] != ele[8][17];
    ele[8][12] != ele[8][18];
    ele[8][12] != ele[8][19];
    ele[8][12] != ele[8][20];
    ele[8][12] != ele[8][21];
    ele[8][12] != ele[8][22];
    ele[8][12] != ele[8][23];
    ele[8][12] != ele[8][24];
    ele[8][12] != ele[9][10];
    ele[8][12] != ele[9][11];
    ele[8][12] != ele[9][12];
    ele[8][12] != ele[9][13];
    ele[8][12] != ele[9][14];
    ele[8][13] != ele[10][13];
    ele[8][13] != ele[11][13];
    ele[8][13] != ele[12][13];
    ele[8][13] != ele[13][13];
    ele[8][13] != ele[14][13];
    ele[8][13] != ele[15][13];
    ele[8][13] != ele[16][13];
    ele[8][13] != ele[17][13];
    ele[8][13] != ele[18][13];
    ele[8][13] != ele[19][13];
    ele[8][13] != ele[20][13];
    ele[8][13] != ele[21][13];
    ele[8][13] != ele[22][13];
    ele[8][13] != ele[23][13];
    ele[8][13] != ele[24][13];
    ele[8][13] != ele[8][14];
    ele[8][13] != ele[8][15];
    ele[8][13] != ele[8][16];
    ele[8][13] != ele[8][17];
    ele[8][13] != ele[8][18];
    ele[8][13] != ele[8][19];
    ele[8][13] != ele[8][20];
    ele[8][13] != ele[8][21];
    ele[8][13] != ele[8][22];
    ele[8][13] != ele[8][23];
    ele[8][13] != ele[8][24];
    ele[8][13] != ele[9][10];
    ele[8][13] != ele[9][11];
    ele[8][13] != ele[9][12];
    ele[8][13] != ele[9][13];
    ele[8][13] != ele[9][14];
    ele[8][14] != ele[10][14];
    ele[8][14] != ele[11][14];
    ele[8][14] != ele[12][14];
    ele[8][14] != ele[13][14];
    ele[8][14] != ele[14][14];
    ele[8][14] != ele[15][14];
    ele[8][14] != ele[16][14];
    ele[8][14] != ele[17][14];
    ele[8][14] != ele[18][14];
    ele[8][14] != ele[19][14];
    ele[8][14] != ele[20][14];
    ele[8][14] != ele[21][14];
    ele[8][14] != ele[22][14];
    ele[8][14] != ele[23][14];
    ele[8][14] != ele[24][14];
    ele[8][14] != ele[8][15];
    ele[8][14] != ele[8][16];
    ele[8][14] != ele[8][17];
    ele[8][14] != ele[8][18];
    ele[8][14] != ele[8][19];
    ele[8][14] != ele[8][20];
    ele[8][14] != ele[8][21];
    ele[8][14] != ele[8][22];
    ele[8][14] != ele[8][23];
    ele[8][14] != ele[8][24];
    ele[8][14] != ele[9][10];
    ele[8][14] != ele[9][11];
    ele[8][14] != ele[9][12];
    ele[8][14] != ele[9][13];
    ele[8][14] != ele[9][14];
    ele[8][15] != ele[10][15];
    ele[8][15] != ele[11][15];
    ele[8][15] != ele[12][15];
    ele[8][15] != ele[13][15];
    ele[8][15] != ele[14][15];
    ele[8][15] != ele[15][15];
    ele[8][15] != ele[16][15];
    ele[8][15] != ele[17][15];
    ele[8][15] != ele[18][15];
    ele[8][15] != ele[19][15];
    ele[8][15] != ele[20][15];
    ele[8][15] != ele[21][15];
    ele[8][15] != ele[22][15];
    ele[8][15] != ele[23][15];
    ele[8][15] != ele[24][15];
    ele[8][15] != ele[8][16];
    ele[8][15] != ele[8][17];
    ele[8][15] != ele[8][18];
    ele[8][15] != ele[8][19];
    ele[8][15] != ele[8][20];
    ele[8][15] != ele[8][21];
    ele[8][15] != ele[8][22];
    ele[8][15] != ele[8][23];
    ele[8][15] != ele[8][24];
    ele[8][15] != ele[9][15];
    ele[8][15] != ele[9][16];
    ele[8][15] != ele[9][17];
    ele[8][15] != ele[9][18];
    ele[8][15] != ele[9][19];
    ele[8][16] != ele[10][16];
    ele[8][16] != ele[11][16];
    ele[8][16] != ele[12][16];
    ele[8][16] != ele[13][16];
    ele[8][16] != ele[14][16];
    ele[8][16] != ele[15][16];
    ele[8][16] != ele[16][16];
    ele[8][16] != ele[17][16];
    ele[8][16] != ele[18][16];
    ele[8][16] != ele[19][16];
    ele[8][16] != ele[20][16];
    ele[8][16] != ele[21][16];
    ele[8][16] != ele[22][16];
    ele[8][16] != ele[23][16];
    ele[8][16] != ele[24][16];
    ele[8][16] != ele[8][17];
    ele[8][16] != ele[8][18];
    ele[8][16] != ele[8][19];
    ele[8][16] != ele[8][20];
    ele[8][16] != ele[8][21];
    ele[8][16] != ele[8][22];
    ele[8][16] != ele[8][23];
    ele[8][16] != ele[8][24];
    ele[8][16] != ele[9][15];
    ele[8][16] != ele[9][16];
    ele[8][16] != ele[9][17];
    ele[8][16] != ele[9][18];
    ele[8][16] != ele[9][19];
    ele[8][17] != ele[10][17];
    ele[8][17] != ele[11][17];
    ele[8][17] != ele[12][17];
    ele[8][17] != ele[13][17];
    ele[8][17] != ele[14][17];
    ele[8][17] != ele[15][17];
    ele[8][17] != ele[16][17];
    ele[8][17] != ele[17][17];
    ele[8][17] != ele[18][17];
    ele[8][17] != ele[19][17];
    ele[8][17] != ele[20][17];
    ele[8][17] != ele[21][17];
    ele[8][17] != ele[22][17];
    ele[8][17] != ele[23][17];
    ele[8][17] != ele[24][17];
    ele[8][17] != ele[8][18];
    ele[8][17] != ele[8][19];
    ele[8][17] != ele[8][20];
    ele[8][17] != ele[8][21];
    ele[8][17] != ele[8][22];
    ele[8][17] != ele[8][23];
    ele[8][17] != ele[8][24];
    ele[8][17] != ele[9][15];
    ele[8][17] != ele[9][16];
    ele[8][17] != ele[9][17];
    ele[8][17] != ele[9][18];
    ele[8][17] != ele[9][19];
    ele[8][18] != ele[10][18];
    ele[8][18] != ele[11][18];
    ele[8][18] != ele[12][18];
    ele[8][18] != ele[13][18];
    ele[8][18] != ele[14][18];
    ele[8][18] != ele[15][18];
    ele[8][18] != ele[16][18];
    ele[8][18] != ele[17][18];
    ele[8][18] != ele[18][18];
    ele[8][18] != ele[19][18];
    ele[8][18] != ele[20][18];
    ele[8][18] != ele[21][18];
    ele[8][18] != ele[22][18];
    ele[8][18] != ele[23][18];
    ele[8][18] != ele[24][18];
    ele[8][18] != ele[8][19];
    ele[8][18] != ele[8][20];
    ele[8][18] != ele[8][21];
    ele[8][18] != ele[8][22];
    ele[8][18] != ele[8][23];
    ele[8][18] != ele[8][24];
    ele[8][18] != ele[9][15];
    ele[8][18] != ele[9][16];
    ele[8][18] != ele[9][17];
    ele[8][18] != ele[9][18];
    ele[8][18] != ele[9][19];
    ele[8][19] != ele[10][19];
    ele[8][19] != ele[11][19];
    ele[8][19] != ele[12][19];
    ele[8][19] != ele[13][19];
    ele[8][19] != ele[14][19];
    ele[8][19] != ele[15][19];
    ele[8][19] != ele[16][19];
    ele[8][19] != ele[17][19];
    ele[8][19] != ele[18][19];
    ele[8][19] != ele[19][19];
    ele[8][19] != ele[20][19];
    ele[8][19] != ele[21][19];
    ele[8][19] != ele[22][19];
    ele[8][19] != ele[23][19];
    ele[8][19] != ele[24][19];
    ele[8][19] != ele[8][20];
    ele[8][19] != ele[8][21];
    ele[8][19] != ele[8][22];
    ele[8][19] != ele[8][23];
    ele[8][19] != ele[8][24];
    ele[8][19] != ele[9][15];
    ele[8][19] != ele[9][16];
    ele[8][19] != ele[9][17];
    ele[8][19] != ele[9][18];
    ele[8][19] != ele[9][19];
    ele[8][2] != ele[10][2];
    ele[8][2] != ele[11][2];
    ele[8][2] != ele[12][2];
    ele[8][2] != ele[13][2];
    ele[8][2] != ele[14][2];
    ele[8][2] != ele[15][2];
    ele[8][2] != ele[16][2];
    ele[8][2] != ele[17][2];
    ele[8][2] != ele[18][2];
    ele[8][2] != ele[19][2];
    ele[8][2] != ele[20][2];
    ele[8][2] != ele[21][2];
    ele[8][2] != ele[22][2];
    ele[8][2] != ele[23][2];
    ele[8][2] != ele[24][2];
    ele[8][2] != ele[8][10];
    ele[8][2] != ele[8][11];
    ele[8][2] != ele[8][12];
    ele[8][2] != ele[8][13];
    ele[8][2] != ele[8][14];
    ele[8][2] != ele[8][15];
    ele[8][2] != ele[8][16];
    ele[8][2] != ele[8][17];
    ele[8][2] != ele[8][18];
    ele[8][2] != ele[8][19];
    ele[8][2] != ele[8][20];
    ele[8][2] != ele[8][21];
    ele[8][2] != ele[8][22];
    ele[8][2] != ele[8][23];
    ele[8][2] != ele[8][24];
    ele[8][2] != ele[8][3];
    ele[8][2] != ele[8][4];
    ele[8][2] != ele[8][5];
    ele[8][2] != ele[8][6];
    ele[8][2] != ele[8][7];
    ele[8][2] != ele[8][8];
    ele[8][2] != ele[8][9];
    ele[8][2] != ele[9][0];
    ele[8][2] != ele[9][1];
    ele[8][2] != ele[9][2];
    ele[8][2] != ele[9][3];
    ele[8][2] != ele[9][4];
    ele[8][20] != ele[10][20];
    ele[8][20] != ele[11][20];
    ele[8][20] != ele[12][20];
    ele[8][20] != ele[13][20];
    ele[8][20] != ele[14][20];
    ele[8][20] != ele[15][20];
    ele[8][20] != ele[16][20];
    ele[8][20] != ele[17][20];
    ele[8][20] != ele[18][20];
    ele[8][20] != ele[19][20];
    ele[8][20] != ele[20][20];
    ele[8][20] != ele[21][20];
    ele[8][20] != ele[22][20];
    ele[8][20] != ele[23][20];
    ele[8][20] != ele[24][20];
    ele[8][20] != ele[8][21];
    ele[8][20] != ele[8][22];
    ele[8][20] != ele[8][23];
    ele[8][20] != ele[8][24];
    ele[8][20] != ele[9][20];
    ele[8][20] != ele[9][21];
    ele[8][20] != ele[9][22];
    ele[8][20] != ele[9][23];
    ele[8][20] != ele[9][24];
    ele[8][21] != ele[10][21];
    ele[8][21] != ele[11][21];
    ele[8][21] != ele[12][21];
    ele[8][21] != ele[13][21];
    ele[8][21] != ele[14][21];
    ele[8][21] != ele[15][21];
    ele[8][21] != ele[16][21];
    ele[8][21] != ele[17][21];
    ele[8][21] != ele[18][21];
    ele[8][21] != ele[19][21];
    ele[8][21] != ele[20][21];
    ele[8][21] != ele[21][21];
    ele[8][21] != ele[22][21];
    ele[8][21] != ele[23][21];
    ele[8][21] != ele[24][21];
    ele[8][21] != ele[8][22];
    ele[8][21] != ele[8][23];
    ele[8][21] != ele[8][24];
    ele[8][21] != ele[9][20];
    ele[8][21] != ele[9][21];
    ele[8][21] != ele[9][22];
    ele[8][21] != ele[9][23];
    ele[8][21] != ele[9][24];
    ele[8][22] != ele[10][22];
    ele[8][22] != ele[11][22];
    ele[8][22] != ele[12][22];
    ele[8][22] != ele[13][22];
    ele[8][22] != ele[14][22];
    ele[8][22] != ele[15][22];
    ele[8][22] != ele[16][22];
    ele[8][22] != ele[17][22];
    ele[8][22] != ele[18][22];
    ele[8][22] != ele[19][22];
    ele[8][22] != ele[20][22];
    ele[8][22] != ele[21][22];
    ele[8][22] != ele[22][22];
    ele[8][22] != ele[23][22];
    ele[8][22] != ele[24][22];
    ele[8][22] != ele[8][23];
    ele[8][22] != ele[8][24];
    ele[8][22] != ele[9][20];
    ele[8][22] != ele[9][21];
    ele[8][22] != ele[9][22];
    ele[8][22] != ele[9][23];
    ele[8][22] != ele[9][24];
    ele[8][23] != ele[10][23];
    ele[8][23] != ele[11][23];
    ele[8][23] != ele[12][23];
    ele[8][23] != ele[13][23];
    ele[8][23] != ele[14][23];
    ele[8][23] != ele[15][23];
    ele[8][23] != ele[16][23];
    ele[8][23] != ele[17][23];
    ele[8][23] != ele[18][23];
    ele[8][23] != ele[19][23];
    ele[8][23] != ele[20][23];
    ele[8][23] != ele[21][23];
    ele[8][23] != ele[22][23];
    ele[8][23] != ele[23][23];
    ele[8][23] != ele[24][23];
    ele[8][23] != ele[8][24];
    ele[8][23] != ele[9][20];
    ele[8][23] != ele[9][21];
    ele[8][23] != ele[9][22];
    ele[8][23] != ele[9][23];
    ele[8][23] != ele[9][24];
    ele[8][24] != ele[10][24];
    ele[8][24] != ele[11][24];
    ele[8][24] != ele[12][24];
    ele[8][24] != ele[13][24];
    ele[8][24] != ele[14][24];
    ele[8][24] != ele[15][24];
    ele[8][24] != ele[16][24];
    ele[8][24] != ele[17][24];
    ele[8][24] != ele[18][24];
    ele[8][24] != ele[19][24];
    ele[8][24] != ele[20][24];
    ele[8][24] != ele[21][24];
    ele[8][24] != ele[22][24];
    ele[8][24] != ele[23][24];
    ele[8][24] != ele[24][24];
    ele[8][24] != ele[9][20];
    ele[8][24] != ele[9][21];
    ele[8][24] != ele[9][22];
    ele[8][24] != ele[9][23];
    ele[8][24] != ele[9][24];
    ele[8][3] != ele[10][3];
    ele[8][3] != ele[11][3];
    ele[8][3] != ele[12][3];
    ele[8][3] != ele[13][3];
    ele[8][3] != ele[14][3];
    ele[8][3] != ele[15][3];
    ele[8][3] != ele[16][3];
    ele[8][3] != ele[17][3];
    ele[8][3] != ele[18][3];
    ele[8][3] != ele[19][3];
    ele[8][3] != ele[20][3];
    ele[8][3] != ele[21][3];
    ele[8][3] != ele[22][3];
    ele[8][3] != ele[23][3];
    ele[8][3] != ele[24][3];
    ele[8][3] != ele[8][10];
    ele[8][3] != ele[8][11];
    ele[8][3] != ele[8][12];
    ele[8][3] != ele[8][13];
    ele[8][3] != ele[8][14];
    ele[8][3] != ele[8][15];
    ele[8][3] != ele[8][16];
    ele[8][3] != ele[8][17];
    ele[8][3] != ele[8][18];
    ele[8][3] != ele[8][19];
    ele[8][3] != ele[8][20];
    ele[8][3] != ele[8][21];
    ele[8][3] != ele[8][22];
    ele[8][3] != ele[8][23];
    ele[8][3] != ele[8][24];
    ele[8][3] != ele[8][4];
    ele[8][3] != ele[8][5];
    ele[8][3] != ele[8][6];
    ele[8][3] != ele[8][7];
    ele[8][3] != ele[8][8];
    ele[8][3] != ele[8][9];
    ele[8][3] != ele[9][0];
    ele[8][3] != ele[9][1];
    ele[8][3] != ele[9][2];
    ele[8][3] != ele[9][3];
    ele[8][3] != ele[9][4];
    ele[8][4] != ele[10][4];
    ele[8][4] != ele[11][4];
    ele[8][4] != ele[12][4];
    ele[8][4] != ele[13][4];
    ele[8][4] != ele[14][4];
    ele[8][4] != ele[15][4];
    ele[8][4] != ele[16][4];
    ele[8][4] != ele[17][4];
    ele[8][4] != ele[18][4];
    ele[8][4] != ele[19][4];
    ele[8][4] != ele[20][4];
    ele[8][4] != ele[21][4];
    ele[8][4] != ele[22][4];
    ele[8][4] != ele[23][4];
    ele[8][4] != ele[24][4];
    ele[8][4] != ele[8][10];
    ele[8][4] != ele[8][11];
    ele[8][4] != ele[8][12];
    ele[8][4] != ele[8][13];
    ele[8][4] != ele[8][14];
    ele[8][4] != ele[8][15];
    ele[8][4] != ele[8][16];
    ele[8][4] != ele[8][17];
    ele[8][4] != ele[8][18];
    ele[8][4] != ele[8][19];
    ele[8][4] != ele[8][20];
    ele[8][4] != ele[8][21];
    ele[8][4] != ele[8][22];
    ele[8][4] != ele[8][23];
    ele[8][4] != ele[8][24];
    ele[8][4] != ele[8][5];
    ele[8][4] != ele[8][6];
    ele[8][4] != ele[8][7];
    ele[8][4] != ele[8][8];
    ele[8][4] != ele[8][9];
    ele[8][4] != ele[9][0];
    ele[8][4] != ele[9][1];
    ele[8][4] != ele[9][2];
    ele[8][4] != ele[9][3];
    ele[8][4] != ele[9][4];
    ele[8][5] != ele[10][5];
    ele[8][5] != ele[11][5];
    ele[8][5] != ele[12][5];
    ele[8][5] != ele[13][5];
    ele[8][5] != ele[14][5];
    ele[8][5] != ele[15][5];
    ele[8][5] != ele[16][5];
    ele[8][5] != ele[17][5];
    ele[8][5] != ele[18][5];
    ele[8][5] != ele[19][5];
    ele[8][5] != ele[20][5];
    ele[8][5] != ele[21][5];
    ele[8][5] != ele[22][5];
    ele[8][5] != ele[23][5];
    ele[8][5] != ele[24][5];
    ele[8][5] != ele[8][10];
    ele[8][5] != ele[8][11];
    ele[8][5] != ele[8][12];
    ele[8][5] != ele[8][13];
    ele[8][5] != ele[8][14];
    ele[8][5] != ele[8][15];
    ele[8][5] != ele[8][16];
    ele[8][5] != ele[8][17];
    ele[8][5] != ele[8][18];
    ele[8][5] != ele[8][19];
    ele[8][5] != ele[8][20];
    ele[8][5] != ele[8][21];
    ele[8][5] != ele[8][22];
    ele[8][5] != ele[8][23];
    ele[8][5] != ele[8][24];
    ele[8][5] != ele[8][6];
    ele[8][5] != ele[8][7];
    ele[8][5] != ele[8][8];
    ele[8][5] != ele[8][9];
    ele[8][5] != ele[9][5];
    ele[8][5] != ele[9][6];
    ele[8][5] != ele[9][7];
    ele[8][5] != ele[9][8];
    ele[8][5] != ele[9][9];
    ele[8][6] != ele[10][6];
    ele[8][6] != ele[11][6];
    ele[8][6] != ele[12][6];
    ele[8][6] != ele[13][6];
    ele[8][6] != ele[14][6];
    ele[8][6] != ele[15][6];
    ele[8][6] != ele[16][6];
    ele[8][6] != ele[17][6];
    ele[8][6] != ele[18][6];
    ele[8][6] != ele[19][6];
    ele[8][6] != ele[20][6];
    ele[8][6] != ele[21][6];
    ele[8][6] != ele[22][6];
    ele[8][6] != ele[23][6];
    ele[8][6] != ele[24][6];
    ele[8][6] != ele[8][10];
    ele[8][6] != ele[8][11];
    ele[8][6] != ele[8][12];
    ele[8][6] != ele[8][13];
    ele[8][6] != ele[8][14];
    ele[8][6] != ele[8][15];
    ele[8][6] != ele[8][16];
    ele[8][6] != ele[8][17];
    ele[8][6] != ele[8][18];
    ele[8][6] != ele[8][19];
    ele[8][6] != ele[8][20];
    ele[8][6] != ele[8][21];
    ele[8][6] != ele[8][22];
    ele[8][6] != ele[8][23];
    ele[8][6] != ele[8][24];
    ele[8][6] != ele[8][7];
    ele[8][6] != ele[8][8];
    ele[8][6] != ele[8][9];
    ele[8][6] != ele[9][5];
    ele[8][6] != ele[9][6];
    ele[8][6] != ele[9][7];
    ele[8][6] != ele[9][8];
    ele[8][6] != ele[9][9];
    ele[8][7] != ele[10][7];
    ele[8][7] != ele[11][7];
    ele[8][7] != ele[12][7];
    ele[8][7] != ele[13][7];
    ele[8][7] != ele[14][7];
    ele[8][7] != ele[15][7];
    ele[8][7] != ele[16][7];
    ele[8][7] != ele[17][7];
    ele[8][7] != ele[18][7];
    ele[8][7] != ele[19][7];
    ele[8][7] != ele[20][7];
    ele[8][7] != ele[21][7];
    ele[8][7] != ele[22][7];
    ele[8][7] != ele[23][7];
    ele[8][7] != ele[24][7];
    ele[8][7] != ele[8][10];
    ele[8][7] != ele[8][11];
    ele[8][7] != ele[8][12];
    ele[8][7] != ele[8][13];
    ele[8][7] != ele[8][14];
    ele[8][7] != ele[8][15];
    ele[8][7] != ele[8][16];
    ele[8][7] != ele[8][17];
    ele[8][7] != ele[8][18];
    ele[8][7] != ele[8][19];
    ele[8][7] != ele[8][20];
    ele[8][7] != ele[8][21];
    ele[8][7] != ele[8][22];
    ele[8][7] != ele[8][23];
    ele[8][7] != ele[8][24];
    ele[8][7] != ele[8][8];
    ele[8][7] != ele[8][9];
    ele[8][7] != ele[9][5];
    ele[8][7] != ele[9][6];
    ele[8][7] != ele[9][7];
    ele[8][7] != ele[9][8];
    ele[8][7] != ele[9][9];
    ele[8][8] != ele[10][8];
    ele[8][8] != ele[11][8];
    ele[8][8] != ele[12][8];
    ele[8][8] != ele[13][8];
    ele[8][8] != ele[14][8];
    ele[8][8] != ele[15][8];
    ele[8][8] != ele[16][8];
    ele[8][8] != ele[17][8];
    ele[8][8] != ele[18][8];
    ele[8][8] != ele[19][8];
    ele[8][8] != ele[20][8];
    ele[8][8] != ele[21][8];
    ele[8][8] != ele[22][8];
    ele[8][8] != ele[23][8];
    ele[8][8] != ele[24][8];
    ele[8][8] != ele[8][10];
    ele[8][8] != ele[8][11];
    ele[8][8] != ele[8][12];
    ele[8][8] != ele[8][13];
    ele[8][8] != ele[8][14];
    ele[8][8] != ele[8][15];
    ele[8][8] != ele[8][16];
    ele[8][8] != ele[8][17];
    ele[8][8] != ele[8][18];
    ele[8][8] != ele[8][19];
    ele[8][8] != ele[8][20];
    ele[8][8] != ele[8][21];
    ele[8][8] != ele[8][22];
    ele[8][8] != ele[8][23];
    ele[8][8] != ele[8][24];
    ele[8][8] != ele[8][9];
    ele[8][8] != ele[9][5];
    ele[8][8] != ele[9][6];
    ele[8][8] != ele[9][7];
    ele[8][8] != ele[9][8];
    ele[8][8] != ele[9][9];
    ele[8][9] != ele[10][9];
    ele[8][9] != ele[11][9];
    ele[8][9] != ele[12][9];
    ele[8][9] != ele[13][9];
    ele[8][9] != ele[14][9];
    ele[8][9] != ele[15][9];
    ele[8][9] != ele[16][9];
    ele[8][9] != ele[17][9];
    ele[8][9] != ele[18][9];
    ele[8][9] != ele[19][9];
    ele[8][9] != ele[20][9];
    ele[8][9] != ele[21][9];
    ele[8][9] != ele[22][9];
    ele[8][9] != ele[23][9];
    ele[8][9] != ele[24][9];
    ele[8][9] != ele[8][10];
    ele[8][9] != ele[8][11];
    ele[8][9] != ele[8][12];
    ele[8][9] != ele[8][13];
    ele[8][9] != ele[8][14];
    ele[8][9] != ele[8][15];
    ele[8][9] != ele[8][16];
    ele[8][9] != ele[8][17];
    ele[8][9] != ele[8][18];
    ele[8][9] != ele[8][19];
    ele[8][9] != ele[8][20];
    ele[8][9] != ele[8][21];
    ele[8][9] != ele[8][22];
    ele[8][9] != ele[8][23];
    ele[8][9] != ele[8][24];
    ele[8][9] != ele[9][5];
    ele[8][9] != ele[9][6];
    ele[8][9] != ele[9][7];
    ele[8][9] != ele[9][8];
    ele[8][9] != ele[9][9];
    ele[9][0] != ele[10][0];
    ele[9][0] != ele[11][0];
    ele[9][0] != ele[12][0];
    ele[9][0] != ele[13][0];
    ele[9][0] != ele[14][0];
    ele[9][0] != ele[15][0];
    ele[9][0] != ele[16][0];
    ele[9][0] != ele[17][0];
    ele[9][0] != ele[18][0];
    ele[9][0] != ele[19][0];
    ele[9][0] != ele[20][0];
    ele[9][0] != ele[21][0];
    ele[9][0] != ele[22][0];
    ele[9][0] != ele[23][0];
    ele[9][0] != ele[24][0];
    ele[9][0] != ele[9][1];
    ele[9][0] != ele[9][10];
    ele[9][0] != ele[9][11];
    ele[9][0] != ele[9][12];
    ele[9][0] != ele[9][13];
    ele[9][0] != ele[9][14];
    ele[9][0] != ele[9][15];
    ele[9][0] != ele[9][16];
    ele[9][0] != ele[9][17];
    ele[9][0] != ele[9][18];
    ele[9][0] != ele[9][19];
    ele[9][0] != ele[9][2];
    ele[9][0] != ele[9][20];
    ele[9][0] != ele[9][21];
    ele[9][0] != ele[9][22];
    ele[9][0] != ele[9][23];
    ele[9][0] != ele[9][24];
    ele[9][0] != ele[9][3];
    ele[9][0] != ele[9][4];
    ele[9][0] != ele[9][5];
    ele[9][0] != ele[9][6];
    ele[9][0] != ele[9][7];
    ele[9][0] != ele[9][8];
    ele[9][0] != ele[9][9];
    ele[9][1] != ele[10][1];
    ele[9][1] != ele[11][1];
    ele[9][1] != ele[12][1];
    ele[9][1] != ele[13][1];
    ele[9][1] != ele[14][1];
    ele[9][1] != ele[15][1];
    ele[9][1] != ele[16][1];
    ele[9][1] != ele[17][1];
    ele[9][1] != ele[18][1];
    ele[9][1] != ele[19][1];
    ele[9][1] != ele[20][1];
    ele[9][1] != ele[21][1];
    ele[9][1] != ele[22][1];
    ele[9][1] != ele[23][1];
    ele[9][1] != ele[24][1];
    ele[9][1] != ele[9][10];
    ele[9][1] != ele[9][11];
    ele[9][1] != ele[9][12];
    ele[9][1] != ele[9][13];
    ele[9][1] != ele[9][14];
    ele[9][1] != ele[9][15];
    ele[9][1] != ele[9][16];
    ele[9][1] != ele[9][17];
    ele[9][1] != ele[9][18];
    ele[9][1] != ele[9][19];
    ele[9][1] != ele[9][2];
    ele[9][1] != ele[9][20];
    ele[9][1] != ele[9][21];
    ele[9][1] != ele[9][22];
    ele[9][1] != ele[9][23];
    ele[9][1] != ele[9][24];
    ele[9][1] != ele[9][3];
    ele[9][1] != ele[9][4];
    ele[9][1] != ele[9][5];
    ele[9][1] != ele[9][6];
    ele[9][1] != ele[9][7];
    ele[9][1] != ele[9][8];
    ele[9][1] != ele[9][9];
    ele[9][10] != ele[10][10];
    ele[9][10] != ele[11][10];
    ele[9][10] != ele[12][10];
    ele[9][10] != ele[13][10];
    ele[9][10] != ele[14][10];
    ele[9][10] != ele[15][10];
    ele[9][10] != ele[16][10];
    ele[9][10] != ele[17][10];
    ele[9][10] != ele[18][10];
    ele[9][10] != ele[19][10];
    ele[9][10] != ele[20][10];
    ele[9][10] != ele[21][10];
    ele[9][10] != ele[22][10];
    ele[9][10] != ele[23][10];
    ele[9][10] != ele[24][10];
    ele[9][10] != ele[9][11];
    ele[9][10] != ele[9][12];
    ele[9][10] != ele[9][13];
    ele[9][10] != ele[9][14];
    ele[9][10] != ele[9][15];
    ele[9][10] != ele[9][16];
    ele[9][10] != ele[9][17];
    ele[9][10] != ele[9][18];
    ele[9][10] != ele[9][19];
    ele[9][10] != ele[9][20];
    ele[9][10] != ele[9][21];
    ele[9][10] != ele[9][22];
    ele[9][10] != ele[9][23];
    ele[9][10] != ele[9][24];
    ele[9][11] != ele[10][11];
    ele[9][11] != ele[11][11];
    ele[9][11] != ele[12][11];
    ele[9][11] != ele[13][11];
    ele[9][11] != ele[14][11];
    ele[9][11] != ele[15][11];
    ele[9][11] != ele[16][11];
    ele[9][11] != ele[17][11];
    ele[9][11] != ele[18][11];
    ele[9][11] != ele[19][11];
    ele[9][11] != ele[20][11];
    ele[9][11] != ele[21][11];
    ele[9][11] != ele[22][11];
    ele[9][11] != ele[23][11];
    ele[9][11] != ele[24][11];
    ele[9][11] != ele[9][12];
    ele[9][11] != ele[9][13];
    ele[9][11] != ele[9][14];
    ele[9][11] != ele[9][15];
    ele[9][11] != ele[9][16];
    ele[9][11] != ele[9][17];
    ele[9][11] != ele[9][18];
    ele[9][11] != ele[9][19];
    ele[9][11] != ele[9][20];
    ele[9][11] != ele[9][21];
    ele[9][11] != ele[9][22];
    ele[9][11] != ele[9][23];
    ele[9][11] != ele[9][24];
    ele[9][12] != ele[10][12];
    ele[9][12] != ele[11][12];
    ele[9][12] != ele[12][12];
    ele[9][12] != ele[13][12];
    ele[9][12] != ele[14][12];
    ele[9][12] != ele[15][12];
    ele[9][12] != ele[16][12];
    ele[9][12] != ele[17][12];
    ele[9][12] != ele[18][12];
    ele[9][12] != ele[19][12];
    ele[9][12] != ele[20][12];
    ele[9][12] != ele[21][12];
    ele[9][12] != ele[22][12];
    ele[9][12] != ele[23][12];
    ele[9][12] != ele[24][12];
    ele[9][12] != ele[9][13];
    ele[9][12] != ele[9][14];
    ele[9][12] != ele[9][15];
    ele[9][12] != ele[9][16];
    ele[9][12] != ele[9][17];
    ele[9][12] != ele[9][18];
    ele[9][12] != ele[9][19];
    ele[9][12] != ele[9][20];
    ele[9][12] != ele[9][21];
    ele[9][12] != ele[9][22];
    ele[9][12] != ele[9][23];
    ele[9][12] != ele[9][24];
    ele[9][13] != ele[10][13];
    ele[9][13] != ele[11][13];
    ele[9][13] != ele[12][13];
    ele[9][13] != ele[13][13];
    ele[9][13] != ele[14][13];
    ele[9][13] != ele[15][13];
    ele[9][13] != ele[16][13];
    ele[9][13] != ele[17][13];
    ele[9][13] != ele[18][13];
    ele[9][13] != ele[19][13];
    ele[9][13] != ele[20][13];
    ele[9][13] != ele[21][13];
    ele[9][13] != ele[22][13];
    ele[9][13] != ele[23][13];
    ele[9][13] != ele[24][13];
    ele[9][13] != ele[9][14];
    ele[9][13] != ele[9][15];
    ele[9][13] != ele[9][16];
    ele[9][13] != ele[9][17];
    ele[9][13] != ele[9][18];
    ele[9][13] != ele[9][19];
    ele[9][13] != ele[9][20];
    ele[9][13] != ele[9][21];
    ele[9][13] != ele[9][22];
    ele[9][13] != ele[9][23];
    ele[9][13] != ele[9][24];
    ele[9][14] != ele[10][14];
    ele[9][14] != ele[11][14];
    ele[9][14] != ele[12][14];
    ele[9][14] != ele[13][14];
    ele[9][14] != ele[14][14];
    ele[9][14] != ele[15][14];
    ele[9][14] != ele[16][14];
    ele[9][14] != ele[17][14];
    ele[9][14] != ele[18][14];
    ele[9][14] != ele[19][14];
    ele[9][14] != ele[20][14];
    ele[9][14] != ele[21][14];
    ele[9][14] != ele[22][14];
    ele[9][14] != ele[23][14];
    ele[9][14] != ele[24][14];
    ele[9][14] != ele[9][15];
    ele[9][14] != ele[9][16];
    ele[9][14] != ele[9][17];
    ele[9][14] != ele[9][18];
    ele[9][14] != ele[9][19];
    ele[9][14] != ele[9][20];
    ele[9][14] != ele[9][21];
    ele[9][14] != ele[9][22];
    ele[9][14] != ele[9][23];
    ele[9][14] != ele[9][24];
    ele[9][15] != ele[10][15];
    ele[9][15] != ele[11][15];
    ele[9][15] != ele[12][15];
    ele[9][15] != ele[13][15];
    ele[9][15] != ele[14][15];
    ele[9][15] != ele[15][15];
    ele[9][15] != ele[16][15];
    ele[9][15] != ele[17][15];
    ele[9][15] != ele[18][15];
    ele[9][15] != ele[19][15];
    ele[9][15] != ele[20][15];
    ele[9][15] != ele[21][15];
    ele[9][15] != ele[22][15];
    ele[9][15] != ele[23][15];
    ele[9][15] != ele[24][15];
    ele[9][15] != ele[9][16];
    ele[9][15] != ele[9][17];
    ele[9][15] != ele[9][18];
    ele[9][15] != ele[9][19];
    ele[9][15] != ele[9][20];
    ele[9][15] != ele[9][21];
    ele[9][15] != ele[9][22];
    ele[9][15] != ele[9][23];
    ele[9][15] != ele[9][24];
    ele[9][16] != ele[10][16];
    ele[9][16] != ele[11][16];
    ele[9][16] != ele[12][16];
    ele[9][16] != ele[13][16];
    ele[9][16] != ele[14][16];
    ele[9][16] != ele[15][16];
    ele[9][16] != ele[16][16];
    ele[9][16] != ele[17][16];
    ele[9][16] != ele[18][16];
    ele[9][16] != ele[19][16];
    ele[9][16] != ele[20][16];
    ele[9][16] != ele[21][16];
    ele[9][16] != ele[22][16];
    ele[9][16] != ele[23][16];
    ele[9][16] != ele[24][16];
    ele[9][16] != ele[9][17];
    ele[9][16] != ele[9][18];
    ele[9][16] != ele[9][19];
    ele[9][16] != ele[9][20];
    ele[9][16] != ele[9][21];
    ele[9][16] != ele[9][22];
    ele[9][16] != ele[9][23];
    ele[9][16] != ele[9][24];
    ele[9][17] != ele[10][17];
    ele[9][17] != ele[11][17];
    ele[9][17] != ele[12][17];
    ele[9][17] != ele[13][17];
    ele[9][17] != ele[14][17];
    ele[9][17] != ele[15][17];
    ele[9][17] != ele[16][17];
    ele[9][17] != ele[17][17];
    ele[9][17] != ele[18][17];
    ele[9][17] != ele[19][17];
    ele[9][17] != ele[20][17];
    ele[9][17] != ele[21][17];
    ele[9][17] != ele[22][17];
    ele[9][17] != ele[23][17];
    ele[9][17] != ele[24][17];
    ele[9][17] != ele[9][18];
    ele[9][17] != ele[9][19];
    ele[9][17] != ele[9][20];
    ele[9][17] != ele[9][21];
    ele[9][17] != ele[9][22];
    ele[9][17] != ele[9][23];
    ele[9][17] != ele[9][24];
    ele[9][18] != ele[10][18];
    ele[9][18] != ele[11][18];
    ele[9][18] != ele[12][18];
    ele[9][18] != ele[13][18];
    ele[9][18] != ele[14][18];
    ele[9][18] != ele[15][18];
    ele[9][18] != ele[16][18];
    ele[9][18] != ele[17][18];
    ele[9][18] != ele[18][18];
    ele[9][18] != ele[19][18];
    ele[9][18] != ele[20][18];
    ele[9][18] != ele[21][18];
    ele[9][18] != ele[22][18];
    ele[9][18] != ele[23][18];
    ele[9][18] != ele[24][18];
    ele[9][18] != ele[9][19];
    ele[9][18] != ele[9][20];
    ele[9][18] != ele[9][21];
    ele[9][18] != ele[9][22];
    ele[9][18] != ele[9][23];
    ele[9][18] != ele[9][24];
    ele[9][19] != ele[10][19];
    ele[9][19] != ele[11][19];
    ele[9][19] != ele[12][19];
    ele[9][19] != ele[13][19];
    ele[9][19] != ele[14][19];
    ele[9][19] != ele[15][19];
    ele[9][19] != ele[16][19];
    ele[9][19] != ele[17][19];
    ele[9][19] != ele[18][19];
    ele[9][19] != ele[19][19];
    ele[9][19] != ele[20][19];
    ele[9][19] != ele[21][19];
    ele[9][19] != ele[22][19];
    ele[9][19] != ele[23][19];
    ele[9][19] != ele[24][19];
    ele[9][19] != ele[9][20];
    ele[9][19] != ele[9][21];
    ele[9][19] != ele[9][22];
    ele[9][19] != ele[9][23];
    ele[9][19] != ele[9][24];
    ele[9][2] != ele[10][2];
    ele[9][2] != ele[11][2];
    ele[9][2] != ele[12][2];
    ele[9][2] != ele[13][2];
    ele[9][2] != ele[14][2];
    ele[9][2] != ele[15][2];
    ele[9][2] != ele[16][2];
    ele[9][2] != ele[17][2];
    ele[9][2] != ele[18][2];
    ele[9][2] != ele[19][2];
    ele[9][2] != ele[20][2];
    ele[9][2] != ele[21][2];
    ele[9][2] != ele[22][2];
    ele[9][2] != ele[23][2];
    ele[9][2] != ele[24][2];
    ele[9][2] != ele[9][10];
    ele[9][2] != ele[9][11];
    ele[9][2] != ele[9][12];
    ele[9][2] != ele[9][13];
    ele[9][2] != ele[9][14];
    ele[9][2] != ele[9][15];
    ele[9][2] != ele[9][16];
    ele[9][2] != ele[9][17];
    ele[9][2] != ele[9][18];
    ele[9][2] != ele[9][19];
    ele[9][2] != ele[9][20];
    ele[9][2] != ele[9][21];
    ele[9][2] != ele[9][22];
    ele[9][2] != ele[9][23];
    ele[9][2] != ele[9][24];
    ele[9][2] != ele[9][3];
    ele[9][2] != ele[9][4];
    ele[9][2] != ele[9][5];
    ele[9][2] != ele[9][6];
    ele[9][2] != ele[9][7];
    ele[9][2] != ele[9][8];
    ele[9][2] != ele[9][9];
    ele[9][20] != ele[10][20];
    ele[9][20] != ele[11][20];
    ele[9][20] != ele[12][20];
    ele[9][20] != ele[13][20];
    ele[9][20] != ele[14][20];
    ele[9][20] != ele[15][20];
    ele[9][20] != ele[16][20];
    ele[9][20] != ele[17][20];
    ele[9][20] != ele[18][20];
    ele[9][20] != ele[19][20];
    ele[9][20] != ele[20][20];
    ele[9][20] != ele[21][20];
    ele[9][20] != ele[22][20];
    ele[9][20] != ele[23][20];
    ele[9][20] != ele[24][20];
    ele[9][20] != ele[9][21];
    ele[9][20] != ele[9][22];
    ele[9][20] != ele[9][23];
    ele[9][20] != ele[9][24];
    ele[9][21] != ele[10][21];
    ele[9][21] != ele[11][21];
    ele[9][21] != ele[12][21];
    ele[9][21] != ele[13][21];
    ele[9][21] != ele[14][21];
    ele[9][21] != ele[15][21];
    ele[9][21] != ele[16][21];
    ele[9][21] != ele[17][21];
    ele[9][21] != ele[18][21];
    ele[9][21] != ele[19][21];
    ele[9][21] != ele[20][21];
    ele[9][21] != ele[21][21];
    ele[9][21] != ele[22][21];
    ele[9][21] != ele[23][21];
    ele[9][21] != ele[24][21];
    ele[9][21] != ele[9][22];
    ele[9][21] != ele[9][23];
    ele[9][21] != ele[9][24];
    ele[9][22] != ele[10][22];
    ele[9][22] != ele[11][22];
    ele[9][22] != ele[12][22];
    ele[9][22] != ele[13][22];
    ele[9][22] != ele[14][22];
    ele[9][22] != ele[15][22];
    ele[9][22] != ele[16][22];
    ele[9][22] != ele[17][22];
    ele[9][22] != ele[18][22];
    ele[9][22] != ele[19][22];
    ele[9][22] != ele[20][22];
    ele[9][22] != ele[21][22];
    ele[9][22] != ele[22][22];
    ele[9][22] != ele[23][22];
    ele[9][22] != ele[24][22];
    ele[9][22] != ele[9][23];
    ele[9][22] != ele[9][24];
    ele[9][23] != ele[10][23];
    ele[9][23] != ele[11][23];
    ele[9][23] != ele[12][23];
    ele[9][23] != ele[13][23];
    ele[9][23] != ele[14][23];
    ele[9][23] != ele[15][23];
    ele[9][23] != ele[16][23];
    ele[9][23] != ele[17][23];
    ele[9][23] != ele[18][23];
    ele[9][23] != ele[19][23];
    ele[9][23] != ele[20][23];
    ele[9][23] != ele[21][23];
    ele[9][23] != ele[22][23];
    ele[9][23] != ele[23][23];
    ele[9][23] != ele[24][23];
    ele[9][23] != ele[9][24];
    ele[9][24] != ele[10][24];
    ele[9][24] != ele[11][24];
    ele[9][24] != ele[12][24];
    ele[9][24] != ele[13][24];
    ele[9][24] != ele[14][24];
    ele[9][24] != ele[15][24];
    ele[9][24] != ele[16][24];
    ele[9][24] != ele[17][24];
    ele[9][24] != ele[18][24];
    ele[9][24] != ele[19][24];
    ele[9][24] != ele[20][24];
    ele[9][24] != ele[21][24];
    ele[9][24] != ele[22][24];
    ele[9][24] != ele[23][24];
    ele[9][24] != ele[24][24];
    ele[9][3] != ele[10][3];
    ele[9][3] != ele[11][3];
    ele[9][3] != ele[12][3];
    ele[9][3] != ele[13][3];
    ele[9][3] != ele[14][3];
    ele[9][3] != ele[15][3];
    ele[9][3] != ele[16][3];
    ele[9][3] != ele[17][3];
    ele[9][3] != ele[18][3];
    ele[9][3] != ele[19][3];
    ele[9][3] != ele[20][3];
    ele[9][3] != ele[21][3];
    ele[9][3] != ele[22][3];
    ele[9][3] != ele[23][3];
    ele[9][3] != ele[24][3];
    ele[9][3] != ele[9][10];
    ele[9][3] != ele[9][11];
    ele[9][3] != ele[9][12];
    ele[9][3] != ele[9][13];
    ele[9][3] != ele[9][14];
    ele[9][3] != ele[9][15];
    ele[9][3] != ele[9][16];
    ele[9][3] != ele[9][17];
    ele[9][3] != ele[9][18];
    ele[9][3] != ele[9][19];
    ele[9][3] != ele[9][20];
    ele[9][3] != ele[9][21];
    ele[9][3] != ele[9][22];
    ele[9][3] != ele[9][23];
    ele[9][3] != ele[9][24];
    ele[9][3] != ele[9][4];
    ele[9][3] != ele[9][5];
    ele[9][3] != ele[9][6];
    ele[9][3] != ele[9][7];
    ele[9][3] != ele[9][8];
    ele[9][3] != ele[9][9];
    ele[9][4] != ele[10][4];
    ele[9][4] != ele[11][4];
    ele[9][4] != ele[12][4];
    ele[9][4] != ele[13][4];
    ele[9][4] != ele[14][4];
    ele[9][4] != ele[15][4];
    ele[9][4] != ele[16][4];
    ele[9][4] != ele[17][4];
    ele[9][4] != ele[18][4];
    ele[9][4] != ele[19][4];
    ele[9][4] != ele[20][4];
    ele[9][4] != ele[21][4];
    ele[9][4] != ele[22][4];
    ele[9][4] != ele[23][4];
    ele[9][4] != ele[24][4];
    ele[9][4] != ele[9][10];
    ele[9][4] != ele[9][11];
    ele[9][4] != ele[9][12];
    ele[9][4] != ele[9][13];
    ele[9][4] != ele[9][14];
    ele[9][4] != ele[9][15];
    ele[9][4] != ele[9][16];
    ele[9][4] != ele[9][17];
    ele[9][4] != ele[9][18];
    ele[9][4] != ele[9][19];
    ele[9][4] != ele[9][20];
    ele[9][4] != ele[9][21];
    ele[9][4] != ele[9][22];
    ele[9][4] != ele[9][23];
    ele[9][4] != ele[9][24];
    ele[9][4] != ele[9][5];
    ele[9][4] != ele[9][6];
    ele[9][4] != ele[9][7];
    ele[9][4] != ele[9][8];
    ele[9][4] != ele[9][9];
    ele[9][5] != ele[10][5];
    ele[9][5] != ele[11][5];
    ele[9][5] != ele[12][5];
    ele[9][5] != ele[13][5];
    ele[9][5] != ele[14][5];
    ele[9][5] != ele[15][5];
    ele[9][5] != ele[16][5];
    ele[9][5] != ele[17][5];
    ele[9][5] != ele[18][5];
    ele[9][5] != ele[19][5];
    ele[9][5] != ele[20][5];
    ele[9][5] != ele[21][5];
    ele[9][5] != ele[22][5];
    ele[9][5] != ele[23][5];
    ele[9][5] != ele[24][5];
    ele[9][5] != ele[9][10];
    ele[9][5] != ele[9][11];
    ele[9][5] != ele[9][12];
    ele[9][5] != ele[9][13];
    ele[9][5] != ele[9][14];
    ele[9][5] != ele[9][15];
    ele[9][5] != ele[9][16];
    ele[9][5] != ele[9][17];
    ele[9][5] != ele[9][18];
    ele[9][5] != ele[9][19];
    ele[9][5] != ele[9][20];
    ele[9][5] != ele[9][21];
    ele[9][5] != ele[9][22];
    ele[9][5] != ele[9][23];
    ele[9][5] != ele[9][24];
    ele[9][5] != ele[9][6];
    ele[9][5] != ele[9][7];
    ele[9][5] != ele[9][8];
    ele[9][5] != ele[9][9];
    ele[9][6] != ele[10][6];
    ele[9][6] != ele[11][6];
    ele[9][6] != ele[12][6];
    ele[9][6] != ele[13][6];
    ele[9][6] != ele[14][6];
    ele[9][6] != ele[15][6];
    ele[9][6] != ele[16][6];
    ele[9][6] != ele[17][6];
    ele[9][6] != ele[18][6];
    ele[9][6] != ele[19][6];
    ele[9][6] != ele[20][6];
    ele[9][6] != ele[21][6];
    ele[9][6] != ele[22][6];
    ele[9][6] != ele[23][6];
    ele[9][6] != ele[24][6];
    ele[9][6] != ele[9][10];
    ele[9][6] != ele[9][11];
    ele[9][6] != ele[9][12];
    ele[9][6] != ele[9][13];
    ele[9][6] != ele[9][14];
    ele[9][6] != ele[9][15];
    ele[9][6] != ele[9][16];
    ele[9][6] != ele[9][17];
    ele[9][6] != ele[9][18];
    ele[9][6] != ele[9][19];
    ele[9][6] != ele[9][20];
    ele[9][6] != ele[9][21];
    ele[9][6] != ele[9][22];
    ele[9][6] != ele[9][23];
    ele[9][6] != ele[9][24];
    ele[9][6] != ele[9][7];
    ele[9][6] != ele[9][8];
    ele[9][6] != ele[9][9];
    ele[9][7] != ele[10][7];
    ele[9][7] != ele[11][7];
    ele[9][7] != ele[12][7];
    ele[9][7] != ele[13][7];
    ele[9][7] != ele[14][7];
    ele[9][7] != ele[15][7];
    ele[9][7] != ele[16][7];
    ele[9][7] != ele[17][7];
    ele[9][7] != ele[18][7];
    ele[9][7] != ele[19][7];
    ele[9][7] != ele[20][7];
    ele[9][7] != ele[21][7];
    ele[9][7] != ele[22][7];
    ele[9][7] != ele[23][7];
    ele[9][7] != ele[24][7];
    ele[9][7] != ele[9][10];
    ele[9][7] != ele[9][11];
    ele[9][7] != ele[9][12];
    ele[9][7] != ele[9][13];
    ele[9][7] != ele[9][14];
    ele[9][7] != ele[9][15];
    ele[9][7] != ele[9][16];
    ele[9][7] != ele[9][17];
    ele[9][7] != ele[9][18];
    ele[9][7] != ele[9][19];
    ele[9][7] != ele[9][20];
    ele[9][7] != ele[9][21];
    ele[9][7] != ele[9][22];
    ele[9][7] != ele[9][23];
    ele[9][7] != ele[9][24];
    ele[9][7] != ele[9][8];
    ele[9][7] != ele[9][9];
    ele[9][8] != ele[10][8];
    ele[9][8] != ele[11][8];
    ele[9][8] != ele[12][8];
    ele[9][8] != ele[13][8];
    ele[9][8] != ele[14][8];
    ele[9][8] != ele[15][8];
    ele[9][8] != ele[16][8];
    ele[9][8] != ele[17][8];
    ele[9][8] != ele[18][8];
    ele[9][8] != ele[19][8];
    ele[9][8] != ele[20][8];
    ele[9][8] != ele[21][8];
    ele[9][8] != ele[22][8];
    ele[9][8] != ele[23][8];
    ele[9][8] != ele[24][8];
    ele[9][8] != ele[9][10];
    ele[9][8] != ele[9][11];
    ele[9][8] != ele[9][12];
    ele[9][8] != ele[9][13];
    ele[9][8] != ele[9][14];
    ele[9][8] != ele[9][15];
    ele[9][8] != ele[9][16];
    ele[9][8] != ele[9][17];
    ele[9][8] != ele[9][18];
    ele[9][8] != ele[9][19];
    ele[9][8] != ele[9][20];
    ele[9][8] != ele[9][21];
    ele[9][8] != ele[9][22];
    ele[9][8] != ele[9][23];
    ele[9][8] != ele[9][24];
    ele[9][8] != ele[9][9];
    ele[9][9] != ele[10][9];
    ele[9][9] != ele[11][9];
    ele[9][9] != ele[12][9];
    ele[9][9] != ele[13][9];
    ele[9][9] != ele[14][9];
    ele[9][9] != ele[15][9];
    ele[9][9] != ele[16][9];
    ele[9][9] != ele[17][9];
    ele[9][9] != ele[18][9];
    ele[9][9] != ele[19][9];
    ele[9][9] != ele[20][9];
    ele[9][9] != ele[21][9];
    ele[9][9] != ele[22][9];
    ele[9][9] != ele[23][9];
    ele[9][9] != ele[24][9];
    ele[9][9] != ele[9][10];
    ele[9][9] != ele[9][11];
    ele[9][9] != ele[9][12];
    ele[9][9] != ele[9][13];
    ele[9][9] != ele[9][14];
    ele[9][9] != ele[9][15];
    ele[9][9] != ele[9][16];
    ele[9][9] != ele[9][17];
    ele[9][9] != ele[9][18];
    ele[9][9] != ele[9][19];
    ele[9][9] != ele[9][20];
    ele[9][9] != ele[9][21];
    ele[9][9] != ele[9][22];
    ele[9][9] != ele[9][23];
    ele[9][9] != ele[9][24];
  // NUMBER OF CONSTRAINTS: 20000
  }
  function new ();
    if (! this.randomize ()) begin
      $display ("ERROR: Randomization failed...!!!");
    end
  endfunction: new
  function show ();
    $display (ele[0][0], ele[0][1], ele[0][2], ele[0][3], ele[0][4], ele[0][5], ele[0][6], ele[0][7], ele[0][8], ele[0][9], ele[0][10], ele[0][11], ele[0][12], ele[0][13], ele[0][14], ele[0][15], ele[0][16], ele[0][17], ele[0][18], ele[0][19], ele[0][20], ele[0][21], ele[0][22], ele[0][23], ele[0][24]);
    $display (ele[1][0], ele[1][1], ele[1][2], ele[1][3], ele[1][4], ele[1][5], ele[1][6], ele[1][7], ele[1][8], ele[1][9], ele[1][10], ele[1][11], ele[1][12], ele[1][13], ele[1][14], ele[1][15], ele[1][16], ele[1][17], ele[1][18], ele[1][19], ele[1][20], ele[1][21], ele[1][22], ele[1][23], ele[1][24]);
    $display (ele[2][0], ele[2][1], ele[2][2], ele[2][3], ele[2][4], ele[2][5], ele[2][6], ele[2][7], ele[2][8], ele[2][9], ele[2][10], ele[2][11], ele[2][12], ele[2][13], ele[2][14], ele[2][15], ele[2][16], ele[2][17], ele[2][18], ele[2][19], ele[2][20], ele[2][21], ele[2][22], ele[2][23], ele[2][24]);
    $display (ele[3][0], ele[3][1], ele[3][2], ele[3][3], ele[3][4], ele[3][5], ele[3][6], ele[3][7], ele[3][8], ele[3][9], ele[3][10], ele[3][11], ele[3][12], ele[3][13], ele[3][14], ele[3][15], ele[3][16], ele[3][17], ele[3][18], ele[3][19], ele[3][20], ele[3][21], ele[3][22], ele[3][23], ele[3][24]);
    $display (ele[4][0], ele[4][1], ele[4][2], ele[4][3], ele[4][4], ele[4][5], ele[4][6], ele[4][7], ele[4][8], ele[4][9], ele[4][10], ele[4][11], ele[4][12], ele[4][13], ele[4][14], ele[4][15], ele[4][16], ele[4][17], ele[4][18], ele[4][19], ele[4][20], ele[4][21], ele[4][22], ele[4][23], ele[4][24]);
    $display (ele[5][0], ele[5][1], ele[5][2], ele[5][3], ele[5][4], ele[5][5], ele[5][6], ele[5][7], ele[5][8], ele[5][9], ele[5][10], ele[5][11], ele[5][12], ele[5][13], ele[5][14], ele[5][15], ele[5][16], ele[5][17], ele[5][18], ele[5][19], ele[5][20], ele[5][21], ele[5][22], ele[5][23], ele[5][24]);
    $display (ele[6][0], ele[6][1], ele[6][2], ele[6][3], ele[6][4], ele[6][5], ele[6][6], ele[6][7], ele[6][8], ele[6][9], ele[6][10], ele[6][11], ele[6][12], ele[6][13], ele[6][14], ele[6][15], ele[6][16], ele[6][17], ele[6][18], ele[6][19], ele[6][20], ele[6][21], ele[6][22], ele[6][23], ele[6][24]);
    $display (ele[7][0], ele[7][1], ele[7][2], ele[7][3], ele[7][4], ele[7][5], ele[7][6], ele[7][7], ele[7][8], ele[7][9], ele[7][10], ele[7][11], ele[7][12], ele[7][13], ele[7][14], ele[7][15], ele[7][16], ele[7][17], ele[7][18], ele[7][19], ele[7][20], ele[7][21], ele[7][22], ele[7][23], ele[7][24]);
    $display (ele[8][0], ele[8][1], ele[8][2], ele[8][3], ele[8][4], ele[8][5], ele[8][6], ele[8][7], ele[8][8], ele[8][9], ele[8][10], ele[8][11], ele[8][12], ele[8][13], ele[8][14], ele[8][15], ele[8][16], ele[8][17], ele[8][18], ele[8][19], ele[8][20], ele[8][21], ele[8][22], ele[8][23], ele[8][24]);
    $display (ele[9][0], ele[9][1], ele[9][2], ele[9][3], ele[9][4], ele[9][5], ele[9][6], ele[9][7], ele[9][8], ele[9][9], ele[9][10], ele[9][11], ele[9][12], ele[9][13], ele[9][14], ele[9][15], ele[9][16], ele[9][17], ele[9][18], ele[9][19], ele[9][20], ele[9][21], ele[9][22], ele[9][23], ele[9][24]);
    $display (ele[10][0], ele[10][1], ele[10][2], ele[10][3], ele[10][4], ele[10][5], ele[10][6], ele[10][7], ele[10][8], ele[10][9], ele[10][10], ele[10][11], ele[10][12], ele[10][13], ele[10][14], ele[10][15], ele[10][16], ele[10][17], ele[10][18], ele[10][19], ele[10][20], ele[10][21], ele[10][22], ele[10][23], ele[10][24]);
    $display (ele[11][0], ele[11][1], ele[11][2], ele[11][3], ele[11][4], ele[11][5], ele[11][6], ele[11][7], ele[11][8], ele[11][9], ele[11][10], ele[11][11], ele[11][12], ele[11][13], ele[11][14], ele[11][15], ele[11][16], ele[11][17], ele[11][18], ele[11][19], ele[11][20], ele[11][21], ele[11][22], ele[11][23], ele[11][24]);
    $display (ele[12][0], ele[12][1], ele[12][2], ele[12][3], ele[12][4], ele[12][5], ele[12][6], ele[12][7], ele[12][8], ele[12][9], ele[12][10], ele[12][11], ele[12][12], ele[12][13], ele[12][14], ele[12][15], ele[12][16], ele[12][17], ele[12][18], ele[12][19], ele[12][20], ele[12][21], ele[12][22], ele[12][23], ele[12][24]);
    $display (ele[13][0], ele[13][1], ele[13][2], ele[13][3], ele[13][4], ele[13][5], ele[13][6], ele[13][7], ele[13][8], ele[13][9], ele[13][10], ele[13][11], ele[13][12], ele[13][13], ele[13][14], ele[13][15], ele[13][16], ele[13][17], ele[13][18], ele[13][19], ele[13][20], ele[13][21], ele[13][22], ele[13][23], ele[13][24]);
    $display (ele[14][0], ele[14][1], ele[14][2], ele[14][3], ele[14][4], ele[14][5], ele[14][6], ele[14][7], ele[14][8], ele[14][9], ele[14][10], ele[14][11], ele[14][12], ele[14][13], ele[14][14], ele[14][15], ele[14][16], ele[14][17], ele[14][18], ele[14][19], ele[14][20], ele[14][21], ele[14][22], ele[14][23], ele[14][24]);
    $display (ele[15][0], ele[15][1], ele[15][2], ele[15][3], ele[15][4], ele[15][5], ele[15][6], ele[15][7], ele[15][8], ele[15][9], ele[15][10], ele[15][11], ele[15][12], ele[15][13], ele[15][14], ele[15][15], ele[15][16], ele[15][17], ele[15][18], ele[15][19], ele[15][20], ele[15][21], ele[15][22], ele[15][23], ele[15][24]);
    $display (ele[16][0], ele[16][1], ele[16][2], ele[16][3], ele[16][4], ele[16][5], ele[16][6], ele[16][7], ele[16][8], ele[16][9], ele[16][10], ele[16][11], ele[16][12], ele[16][13], ele[16][14], ele[16][15], ele[16][16], ele[16][17], ele[16][18], ele[16][19], ele[16][20], ele[16][21], ele[16][22], ele[16][23], ele[16][24]);
    $display (ele[17][0], ele[17][1], ele[17][2], ele[17][3], ele[17][4], ele[17][5], ele[17][6], ele[17][7], ele[17][8], ele[17][9], ele[17][10], ele[17][11], ele[17][12], ele[17][13], ele[17][14], ele[17][15], ele[17][16], ele[17][17], ele[17][18], ele[17][19], ele[17][20], ele[17][21], ele[17][22], ele[17][23], ele[17][24]);
    $display (ele[18][0], ele[18][1], ele[18][2], ele[18][3], ele[18][4], ele[18][5], ele[18][6], ele[18][7], ele[18][8], ele[18][9], ele[18][10], ele[18][11], ele[18][12], ele[18][13], ele[18][14], ele[18][15], ele[18][16], ele[18][17], ele[18][18], ele[18][19], ele[18][20], ele[18][21], ele[18][22], ele[18][23], ele[18][24]);
    $display (ele[19][0], ele[19][1], ele[19][2], ele[19][3], ele[19][4], ele[19][5], ele[19][6], ele[19][7], ele[19][8], ele[19][9], ele[19][10], ele[19][11], ele[19][12], ele[19][13], ele[19][14], ele[19][15], ele[19][16], ele[19][17], ele[19][18], ele[19][19], ele[19][20], ele[19][21], ele[19][22], ele[19][23], ele[19][24]);
    $display (ele[20][0], ele[20][1], ele[20][2], ele[20][3], ele[20][4], ele[20][5], ele[20][6], ele[20][7], ele[20][8], ele[20][9], ele[20][10], ele[20][11], ele[20][12], ele[20][13], ele[20][14], ele[20][15], ele[20][16], ele[20][17], ele[20][18], ele[20][19], ele[20][20], ele[20][21], ele[20][22], ele[20][23], ele[20][24]);
    $display (ele[21][0], ele[21][1], ele[21][2], ele[21][3], ele[21][4], ele[21][5], ele[21][6], ele[21][7], ele[21][8], ele[21][9], ele[21][10], ele[21][11], ele[21][12], ele[21][13], ele[21][14], ele[21][15], ele[21][16], ele[21][17], ele[21][18], ele[21][19], ele[21][20], ele[21][21], ele[21][22], ele[21][23], ele[21][24]);
    $display (ele[22][0], ele[22][1], ele[22][2], ele[22][3], ele[22][4], ele[22][5], ele[22][6], ele[22][7], ele[22][8], ele[22][9], ele[22][10], ele[22][11], ele[22][12], ele[22][13], ele[22][14], ele[22][15], ele[22][16], ele[22][17], ele[22][18], ele[22][19], ele[22][20], ele[22][21], ele[22][22], ele[22][23], ele[22][24]);
    $display (ele[23][0], ele[23][1], ele[23][2], ele[23][3], ele[23][4], ele[23][5], ele[23][6], ele[23][7], ele[23][8], ele[23][9], ele[23][10], ele[23][11], ele[23][12], ele[23][13], ele[23][14], ele[23][15], ele[23][16], ele[23][17], ele[23][18], ele[23][19], ele[23][20], ele[23][21], ele[23][22], ele[23][23], ele[23][24]);
    $display (ele[24][0], ele[24][1], ele[24][2], ele[24][3], ele[24][4], ele[24][5], ele[24][6], ele[24][7], ele[24][8], ele[24][9], ele[24][10], ele[24][11], ele[24][12], ele[24][13], ele[24][14], ele[24][15], ele[24][16], ele[24][17], ele[24][18], ele[24][19], ele[24][20], ele[24][21], ele[24][22], ele[24][23], ele[24][24]);
  endfunction: show
endclass: board
