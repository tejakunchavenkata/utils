class board;
  typedef enum {
    AAA=1,
    AAB=2,
    AAC=3,
    AAD=4,
    AAE=5,
    AAF=6,
    AAG=7,
    AAH=8,
    AAI
  } elements;
  rand elements ele[9][9];
  constraint all {
    ele[0][0] != ele[0][1];
    ele[0][0] != ele[0][2];
    ele[0][0] != ele[0][3];
    ele[0][0] != ele[0][4];
    ele[0][0] != ele[0][5];
    ele[0][0] != ele[0][6];
    ele[0][0] != ele[0][7];
    ele[0][0] != ele[0][8];
    ele[0][0] != ele[1][0];
    ele[0][0] != ele[1][1];
    ele[0][0] != ele[1][2];
    ele[0][0] != ele[2][0];
    ele[0][0] != ele[2][1];
    ele[0][0] != ele[2][2];
    ele[0][0] != ele[3][0];
    ele[0][0] != ele[4][0];
    ele[0][0] != ele[5][0];
    ele[0][0] != ele[6][0];
    ele[0][0] != ele[7][0];
    ele[0][0] != ele[8][0];
    ele[0][1] != ele[0][2];
    ele[0][1] != ele[0][3];
    ele[0][1] != ele[0][4];
    ele[0][1] != ele[0][5];
    ele[0][1] != ele[0][6];
    ele[0][1] != ele[0][7];
    ele[0][1] != ele[0][8];
    ele[0][1] != ele[1][0];
    ele[0][1] != ele[1][1];
    ele[0][1] != ele[1][2];
    ele[0][1] != ele[2][0];
    ele[0][1] != ele[2][1];
    ele[0][1] != ele[2][2];
    ele[0][1] != ele[3][1];
    ele[0][1] != ele[4][1];
    ele[0][1] != ele[5][1];
    ele[0][1] != ele[6][1];
    ele[0][1] != ele[7][1];
    ele[0][1] != ele[8][1];
    ele[0][2] != ele[0][3];
    ele[0][2] != ele[0][4];
    ele[0][2] != ele[0][5];
    ele[0][2] != ele[0][6];
    ele[0][2] != ele[0][7];
    ele[0][2] != ele[0][8];
    ele[0][2] != ele[1][0];
    ele[0][2] != ele[1][1];
    ele[0][2] != ele[1][2];
    ele[0][2] != ele[2][0];
    ele[0][2] != ele[2][1];
    ele[0][2] != ele[2][2];
    ele[0][2] != ele[3][2];
    ele[0][2] != ele[4][2];
    ele[0][2] != ele[5][2];
    ele[0][2] != ele[6][2];
    ele[0][2] != ele[7][2];
    ele[0][2] != ele[8][2];
    ele[0][3] != ele[0][4];
    ele[0][3] != ele[0][5];
    ele[0][3] != ele[0][6];
    ele[0][3] != ele[0][7];
    ele[0][3] != ele[0][8];
    ele[0][3] != ele[1][3];
    ele[0][3] != ele[1][4];
    ele[0][3] != ele[1][5];
    ele[0][3] != ele[2][3];
    ele[0][3] != ele[2][4];
    ele[0][3] != ele[2][5];
    ele[0][3] != ele[3][3];
    ele[0][3] != ele[4][3];
    ele[0][3] != ele[5][3];
    ele[0][3] != ele[6][3];
    ele[0][3] != ele[7][3];
    ele[0][3] != ele[8][3];
    ele[0][4] != ele[0][5];
    ele[0][4] != ele[0][6];
    ele[0][4] != ele[0][7];
    ele[0][4] != ele[0][8];
    ele[0][4] != ele[1][3];
    ele[0][4] != ele[1][4];
    ele[0][4] != ele[1][5];
    ele[0][4] != ele[2][3];
    ele[0][4] != ele[2][4];
    ele[0][4] != ele[2][5];
    ele[0][4] != ele[3][4];
    ele[0][4] != ele[4][4];
    ele[0][4] != ele[5][4];
    ele[0][4] != ele[6][4];
    ele[0][4] != ele[7][4];
    ele[0][4] != ele[8][4];
    ele[0][5] != ele[0][6];
    ele[0][5] != ele[0][7];
    ele[0][5] != ele[0][8];
    ele[0][5] != ele[1][3];
    ele[0][5] != ele[1][4];
    ele[0][5] != ele[1][5];
    ele[0][5] != ele[2][3];
    ele[0][5] != ele[2][4];
    ele[0][5] != ele[2][5];
    ele[0][5] != ele[3][5];
    ele[0][5] != ele[4][5];
    ele[0][5] != ele[5][5];
    ele[0][5] != ele[6][5];
    ele[0][5] != ele[7][5];
    ele[0][5] != ele[8][5];
    ele[0][6] != ele[0][7];
    ele[0][6] != ele[0][8];
    ele[0][6] != ele[1][6];
    ele[0][6] != ele[1][7];
    ele[0][6] != ele[1][8];
    ele[0][6] != ele[2][6];
    ele[0][6] != ele[2][7];
    ele[0][6] != ele[2][8];
    ele[0][6] != ele[3][6];
    ele[0][6] != ele[4][6];
    ele[0][6] != ele[5][6];
    ele[0][6] != ele[6][6];
    ele[0][6] != ele[7][6];
    ele[0][6] != ele[8][6];
    ele[0][7] != ele[0][8];
    ele[0][7] != ele[1][6];
    ele[0][7] != ele[1][7];
    ele[0][7] != ele[1][8];
    ele[0][7] != ele[2][6];
    ele[0][7] != ele[2][7];
    ele[0][7] != ele[2][8];
    ele[0][7] != ele[3][7];
    ele[0][7] != ele[4][7];
    ele[0][7] != ele[5][7];
    ele[0][7] != ele[6][7];
    ele[0][7] != ele[7][7];
    ele[0][7] != ele[8][7];
    ele[0][8] != ele[1][6];
    ele[0][8] != ele[1][7];
    ele[0][8] != ele[1][8];
    ele[0][8] != ele[2][6];
    ele[0][8] != ele[2][7];
    ele[0][8] != ele[2][8];
    ele[0][8] != ele[3][8];
    ele[0][8] != ele[4][8];
    ele[0][8] != ele[5][8];
    ele[0][8] != ele[6][8];
    ele[0][8] != ele[7][8];
    ele[0][8] != ele[8][8];
    ele[1][0] != ele[1][1];
    ele[1][0] != ele[1][2];
    ele[1][0] != ele[1][3];
    ele[1][0] != ele[1][4];
    ele[1][0] != ele[1][5];
    ele[1][0] != ele[1][6];
    ele[1][0] != ele[1][7];
    ele[1][0] != ele[1][8];
    ele[1][0] != ele[2][0];
    ele[1][0] != ele[2][1];
    ele[1][0] != ele[2][2];
    ele[1][0] != ele[3][0];
    ele[1][0] != ele[4][0];
    ele[1][0] != ele[5][0];
    ele[1][0] != ele[6][0];
    ele[1][0] != ele[7][0];
    ele[1][0] != ele[8][0];
    ele[1][1] != ele[1][2];
    ele[1][1] != ele[1][3];
    ele[1][1] != ele[1][4];
    ele[1][1] != ele[1][5];
    ele[1][1] != ele[1][6];
    ele[1][1] != ele[1][7];
    ele[1][1] != ele[1][8];
    ele[1][1] != ele[2][0];
    ele[1][1] != ele[2][1];
    ele[1][1] != ele[2][2];
    ele[1][1] != ele[3][1];
    ele[1][1] != ele[4][1];
    ele[1][1] != ele[5][1];
    ele[1][1] != ele[6][1];
    ele[1][1] != ele[7][1];
    ele[1][1] != ele[8][1];
    ele[1][2] != ele[1][3];
    ele[1][2] != ele[1][4];
    ele[1][2] != ele[1][5];
    ele[1][2] != ele[1][6];
    ele[1][2] != ele[1][7];
    ele[1][2] != ele[1][8];
    ele[1][2] != ele[2][0];
    ele[1][2] != ele[2][1];
    ele[1][2] != ele[2][2];
    ele[1][2] != ele[3][2];
    ele[1][2] != ele[4][2];
    ele[1][2] != ele[5][2];
    ele[1][2] != ele[6][2];
    ele[1][2] != ele[7][2];
    ele[1][2] != ele[8][2];
    ele[1][3] != ele[1][4];
    ele[1][3] != ele[1][5];
    ele[1][3] != ele[1][6];
    ele[1][3] != ele[1][7];
    ele[1][3] != ele[1][8];
    ele[1][3] != ele[2][3];
    ele[1][3] != ele[2][4];
    ele[1][3] != ele[2][5];
    ele[1][3] != ele[3][3];
    ele[1][3] != ele[4][3];
    ele[1][3] != ele[5][3];
    ele[1][3] != ele[6][3];
    ele[1][3] != ele[7][3];
    ele[1][3] != ele[8][3];
    ele[1][4] != ele[1][5];
    ele[1][4] != ele[1][6];
    ele[1][4] != ele[1][7];
    ele[1][4] != ele[1][8];
    ele[1][4] != ele[2][3];
    ele[1][4] != ele[2][4];
    ele[1][4] != ele[2][5];
    ele[1][4] != ele[3][4];
    ele[1][4] != ele[4][4];
    ele[1][4] != ele[5][4];
    ele[1][4] != ele[6][4];
    ele[1][4] != ele[7][4];
    ele[1][4] != ele[8][4];
    ele[1][5] != ele[1][6];
    ele[1][5] != ele[1][7];
    ele[1][5] != ele[1][8];
    ele[1][5] != ele[2][3];
    ele[1][5] != ele[2][4];
    ele[1][5] != ele[2][5];
    ele[1][5] != ele[3][5];
    ele[1][5] != ele[4][5];
    ele[1][5] != ele[5][5];
    ele[1][5] != ele[6][5];
    ele[1][5] != ele[7][5];
    ele[1][5] != ele[8][5];
    ele[1][6] != ele[1][7];
    ele[1][6] != ele[1][8];
    ele[1][6] != ele[2][6];
    ele[1][6] != ele[2][7];
    ele[1][6] != ele[2][8];
    ele[1][6] != ele[3][6];
    ele[1][6] != ele[4][6];
    ele[1][6] != ele[5][6];
    ele[1][6] != ele[6][6];
    ele[1][6] != ele[7][6];
    ele[1][6] != ele[8][6];
    ele[1][7] != ele[1][8];
    ele[1][7] != ele[2][6];
    ele[1][7] != ele[2][7];
    ele[1][7] != ele[2][8];
    ele[1][7] != ele[3][7];
    ele[1][7] != ele[4][7];
    ele[1][7] != ele[5][7];
    ele[1][7] != ele[6][7];
    ele[1][7] != ele[7][7];
    ele[1][7] != ele[8][7];
    ele[1][8] != ele[2][6];
    ele[1][8] != ele[2][7];
    ele[1][8] != ele[2][8];
    ele[1][8] != ele[3][8];
    ele[1][8] != ele[4][8];
    ele[1][8] != ele[5][8];
    ele[1][8] != ele[6][8];
    ele[1][8] != ele[7][8];
    ele[1][8] != ele[8][8];
    ele[2][0] != ele[2][1];
    ele[2][0] != ele[2][2];
    ele[2][0] != ele[2][3];
    ele[2][0] != ele[2][4];
    ele[2][0] != ele[2][5];
    ele[2][0] != ele[2][6];
    ele[2][0] != ele[2][7];
    ele[2][0] != ele[2][8];
    ele[2][0] != ele[3][0];
    ele[2][0] != ele[4][0];
    ele[2][0] != ele[5][0];
    ele[2][0] != ele[6][0];
    ele[2][0] != ele[7][0];
    ele[2][0] != ele[8][0];
    ele[2][1] != ele[2][2];
    ele[2][1] != ele[2][3];
    ele[2][1] != ele[2][4];
    ele[2][1] != ele[2][5];
    ele[2][1] != ele[2][6];
    ele[2][1] != ele[2][7];
    ele[2][1] != ele[2][8];
    ele[2][1] != ele[3][1];
    ele[2][1] != ele[4][1];
    ele[2][1] != ele[5][1];
    ele[2][1] != ele[6][1];
    ele[2][1] != ele[7][1];
    ele[2][1] != ele[8][1];
    ele[2][2] != ele[2][3];
    ele[2][2] != ele[2][4];
    ele[2][2] != ele[2][5];
    ele[2][2] != ele[2][6];
    ele[2][2] != ele[2][7];
    ele[2][2] != ele[2][8];
    ele[2][2] != ele[3][2];
    ele[2][2] != ele[4][2];
    ele[2][2] != ele[5][2];
    ele[2][2] != ele[6][2];
    ele[2][2] != ele[7][2];
    ele[2][2] != ele[8][2];
    ele[2][3] != ele[2][4];
    ele[2][3] != ele[2][5];
    ele[2][3] != ele[2][6];
    ele[2][3] != ele[2][7];
    ele[2][3] != ele[2][8];
    ele[2][3] != ele[3][3];
    ele[2][3] != ele[4][3];
    ele[2][3] != ele[5][3];
    ele[2][3] != ele[6][3];
    ele[2][3] != ele[7][3];
    ele[2][3] != ele[8][3];
    ele[2][4] != ele[2][5];
    ele[2][4] != ele[2][6];
    ele[2][4] != ele[2][7];
    ele[2][4] != ele[2][8];
    ele[2][4] != ele[3][4];
    ele[2][4] != ele[4][4];
    ele[2][4] != ele[5][4];
    ele[2][4] != ele[6][4];
    ele[2][4] != ele[7][4];
    ele[2][4] != ele[8][4];
    ele[2][5] != ele[2][6];
    ele[2][5] != ele[2][7];
    ele[2][5] != ele[2][8];
    ele[2][5] != ele[3][5];
    ele[2][5] != ele[4][5];
    ele[2][5] != ele[5][5];
    ele[2][5] != ele[6][5];
    ele[2][5] != ele[7][5];
    ele[2][5] != ele[8][5];
    ele[2][6] != ele[2][7];
    ele[2][6] != ele[2][8];
    ele[2][6] != ele[3][6];
    ele[2][6] != ele[4][6];
    ele[2][6] != ele[5][6];
    ele[2][6] != ele[6][6];
    ele[2][6] != ele[7][6];
    ele[2][6] != ele[8][6];
    ele[2][7] != ele[2][8];
    ele[2][7] != ele[3][7];
    ele[2][7] != ele[4][7];
    ele[2][7] != ele[5][7];
    ele[2][7] != ele[6][7];
    ele[2][7] != ele[7][7];
    ele[2][7] != ele[8][7];
    ele[2][8] != ele[3][8];
    ele[2][8] != ele[4][8];
    ele[2][8] != ele[5][8];
    ele[2][8] != ele[6][8];
    ele[2][8] != ele[7][8];
    ele[2][8] != ele[8][8];
    ele[3][0] != ele[3][1];
    ele[3][0] != ele[3][2];
    ele[3][0] != ele[3][3];
    ele[3][0] != ele[3][4];
    ele[3][0] != ele[3][5];
    ele[3][0] != ele[3][6];
    ele[3][0] != ele[3][7];
    ele[3][0] != ele[3][8];
    ele[3][0] != ele[4][0];
    ele[3][0] != ele[4][1];
    ele[3][0] != ele[4][2];
    ele[3][0] != ele[5][0];
    ele[3][0] != ele[5][1];
    ele[3][0] != ele[5][2];
    ele[3][0] != ele[6][0];
    ele[3][0] != ele[7][0];
    ele[3][0] != ele[8][0];
    ele[3][1] != ele[3][2];
    ele[3][1] != ele[3][3];
    ele[3][1] != ele[3][4];
    ele[3][1] != ele[3][5];
    ele[3][1] != ele[3][6];
    ele[3][1] != ele[3][7];
    ele[3][1] != ele[3][8];
    ele[3][1] != ele[4][0];
    ele[3][1] != ele[4][1];
    ele[3][1] != ele[4][2];
    ele[3][1] != ele[5][0];
    ele[3][1] != ele[5][1];
    ele[3][1] != ele[5][2];
    ele[3][1] != ele[6][1];
    ele[3][1] != ele[7][1];
    ele[3][1] != ele[8][1];
    ele[3][2] != ele[3][3];
    ele[3][2] != ele[3][4];
    ele[3][2] != ele[3][5];
    ele[3][2] != ele[3][6];
    ele[3][2] != ele[3][7];
    ele[3][2] != ele[3][8];
    ele[3][2] != ele[4][0];
    ele[3][2] != ele[4][1];
    ele[3][2] != ele[4][2];
    ele[3][2] != ele[5][0];
    ele[3][2] != ele[5][1];
    ele[3][2] != ele[5][2];
    ele[3][2] != ele[6][2];
    ele[3][2] != ele[7][2];
    ele[3][2] != ele[8][2];
    ele[3][3] != ele[3][4];
    ele[3][3] != ele[3][5];
    ele[3][3] != ele[3][6];
    ele[3][3] != ele[3][7];
    ele[3][3] != ele[3][8];
    ele[3][3] != ele[4][3];
    ele[3][3] != ele[4][4];
    ele[3][3] != ele[4][5];
    ele[3][3] != ele[5][3];
    ele[3][3] != ele[5][4];
    ele[3][3] != ele[5][5];
    ele[3][3] != ele[6][3];
    ele[3][3] != ele[7][3];
    ele[3][3] != ele[8][3];
    ele[3][4] != ele[3][5];
    ele[3][4] != ele[3][6];
    ele[3][4] != ele[3][7];
    ele[3][4] != ele[3][8];
    ele[3][4] != ele[4][3];
    ele[3][4] != ele[4][4];
    ele[3][4] != ele[4][5];
    ele[3][4] != ele[5][3];
    ele[3][4] != ele[5][4];
    ele[3][4] != ele[5][5];
    ele[3][4] != ele[6][4];
    ele[3][4] != ele[7][4];
    ele[3][4] != ele[8][4];
    ele[3][5] != ele[3][6];
    ele[3][5] != ele[3][7];
    ele[3][5] != ele[3][8];
    ele[3][5] != ele[4][3];
    ele[3][5] != ele[4][4];
    ele[3][5] != ele[4][5];
    ele[3][5] != ele[5][3];
    ele[3][5] != ele[5][4];
    ele[3][5] != ele[5][5];
    ele[3][5] != ele[6][5];
    ele[3][5] != ele[7][5];
    ele[3][5] != ele[8][5];
    ele[3][6] != ele[3][7];
    ele[3][6] != ele[3][8];
    ele[3][6] != ele[4][6];
    ele[3][6] != ele[4][7];
    ele[3][6] != ele[4][8];
    ele[3][6] != ele[5][6];
    ele[3][6] != ele[5][7];
    ele[3][6] != ele[5][8];
    ele[3][6] != ele[6][6];
    ele[3][6] != ele[7][6];
    ele[3][6] != ele[8][6];
    ele[3][7] != ele[3][8];
    ele[3][7] != ele[4][6];
    ele[3][7] != ele[4][7];
    ele[3][7] != ele[4][8];
    ele[3][7] != ele[5][6];
    ele[3][7] != ele[5][7];
    ele[3][7] != ele[5][8];
    ele[3][7] != ele[6][7];
    ele[3][7] != ele[7][7];
    ele[3][7] != ele[8][7];
    ele[3][8] != ele[4][6];
    ele[3][8] != ele[4][7];
    ele[3][8] != ele[4][8];
    ele[3][8] != ele[5][6];
    ele[3][8] != ele[5][7];
    ele[3][8] != ele[5][8];
    ele[3][8] != ele[6][8];
    ele[3][8] != ele[7][8];
    ele[3][8] != ele[8][8];
    ele[4][0] != ele[4][1];
    ele[4][0] != ele[4][2];
    ele[4][0] != ele[4][3];
    ele[4][0] != ele[4][4];
    ele[4][0] != ele[4][5];
    ele[4][0] != ele[4][6];
    ele[4][0] != ele[4][7];
    ele[4][0] != ele[4][8];
    ele[4][0] != ele[5][0];
    ele[4][0] != ele[5][1];
    ele[4][0] != ele[5][2];
    ele[4][0] != ele[6][0];
    ele[4][0] != ele[7][0];
    ele[4][0] != ele[8][0];
    ele[4][1] != ele[4][2];
    ele[4][1] != ele[4][3];
    ele[4][1] != ele[4][4];
    ele[4][1] != ele[4][5];
    ele[4][1] != ele[4][6];
    ele[4][1] != ele[4][7];
    ele[4][1] != ele[4][8];
    ele[4][1] != ele[5][0];
    ele[4][1] != ele[5][1];
    ele[4][1] != ele[5][2];
    ele[4][1] != ele[6][1];
    ele[4][1] != ele[7][1];
    ele[4][1] != ele[8][1];
    ele[4][2] != ele[4][3];
    ele[4][2] != ele[4][4];
    ele[4][2] != ele[4][5];
    ele[4][2] != ele[4][6];
    ele[4][2] != ele[4][7];
    ele[4][2] != ele[4][8];
    ele[4][2] != ele[5][0];
    ele[4][2] != ele[5][1];
    ele[4][2] != ele[5][2];
    ele[4][2] != ele[6][2];
    ele[4][2] != ele[7][2];
    ele[4][2] != ele[8][2];
    ele[4][3] != ele[4][4];
    ele[4][3] != ele[4][5];
    ele[4][3] != ele[4][6];
    ele[4][3] != ele[4][7];
    ele[4][3] != ele[4][8];
    ele[4][3] != ele[5][3];
    ele[4][3] != ele[5][4];
    ele[4][3] != ele[5][5];
    ele[4][3] != ele[6][3];
    ele[4][3] != ele[7][3];
    ele[4][3] != ele[8][3];
    ele[4][4] != ele[4][5];
    ele[4][4] != ele[4][6];
    ele[4][4] != ele[4][7];
    ele[4][4] != ele[4][8];
    ele[4][4] != ele[5][3];
    ele[4][4] != ele[5][4];
    ele[4][4] != ele[5][5];
    ele[4][4] != ele[6][4];
    ele[4][4] != ele[7][4];
    ele[4][4] != ele[8][4];
    ele[4][5] != ele[4][6];
    ele[4][5] != ele[4][7];
    ele[4][5] != ele[4][8];
    ele[4][5] != ele[5][3];
    ele[4][5] != ele[5][4];
    ele[4][5] != ele[5][5];
    ele[4][5] != ele[6][5];
    ele[4][5] != ele[7][5];
    ele[4][5] != ele[8][5];
    ele[4][6] != ele[4][7];
    ele[4][6] != ele[4][8];
    ele[4][6] != ele[5][6];
    ele[4][6] != ele[5][7];
    ele[4][6] != ele[5][8];
    ele[4][6] != ele[6][6];
    ele[4][6] != ele[7][6];
    ele[4][6] != ele[8][6];
    ele[4][7] != ele[4][8];
    ele[4][7] != ele[5][6];
    ele[4][7] != ele[5][7];
    ele[4][7] != ele[5][8];
    ele[4][7] != ele[6][7];
    ele[4][7] != ele[7][7];
    ele[4][7] != ele[8][7];
    ele[4][8] != ele[5][6];
    ele[4][8] != ele[5][7];
    ele[4][8] != ele[5][8];
    ele[4][8] != ele[6][8];
    ele[4][8] != ele[7][8];
    ele[4][8] != ele[8][8];
    ele[5][0] != ele[5][1];
    ele[5][0] != ele[5][2];
    ele[5][0] != ele[5][3];
    ele[5][0] != ele[5][4];
    ele[5][0] != ele[5][5];
    ele[5][0] != ele[5][6];
    ele[5][0] != ele[5][7];
    ele[5][0] != ele[5][8];
    ele[5][0] != ele[6][0];
    ele[5][0] != ele[7][0];
    ele[5][0] != ele[8][0];
    ele[5][1] != ele[5][2];
    ele[5][1] != ele[5][3];
    ele[5][1] != ele[5][4];
    ele[5][1] != ele[5][5];
    ele[5][1] != ele[5][6];
    ele[5][1] != ele[5][7];
    ele[5][1] != ele[5][8];
    ele[5][1] != ele[6][1];
    ele[5][1] != ele[7][1];
    ele[5][1] != ele[8][1];
    ele[5][2] != ele[5][3];
    ele[5][2] != ele[5][4];
    ele[5][2] != ele[5][5];
    ele[5][2] != ele[5][6];
    ele[5][2] != ele[5][7];
    ele[5][2] != ele[5][8];
    ele[5][2] != ele[6][2];
    ele[5][2] != ele[7][2];
    ele[5][2] != ele[8][2];
    ele[5][3] != ele[5][4];
    ele[5][3] != ele[5][5];
    ele[5][3] != ele[5][6];
    ele[5][3] != ele[5][7];
    ele[5][3] != ele[5][8];
    ele[5][3] != ele[6][3];
    ele[5][3] != ele[7][3];
    ele[5][3] != ele[8][3];
    ele[5][4] != ele[5][5];
    ele[5][4] != ele[5][6];
    ele[5][4] != ele[5][7];
    ele[5][4] != ele[5][8];
    ele[5][4] != ele[6][4];
    ele[5][4] != ele[7][4];
    ele[5][4] != ele[8][4];
    ele[5][5] != ele[5][6];
    ele[5][5] != ele[5][7];
    ele[5][5] != ele[5][8];
    ele[5][5] != ele[6][5];
    ele[5][5] != ele[7][5];
    ele[5][5] != ele[8][5];
    ele[5][6] != ele[5][7];
    ele[5][6] != ele[5][8];
    ele[5][6] != ele[6][6];
    ele[5][6] != ele[7][6];
    ele[5][6] != ele[8][6];
    ele[5][7] != ele[5][8];
    ele[5][7] != ele[6][7];
    ele[5][7] != ele[7][7];
    ele[5][7] != ele[8][7];
    ele[5][8] != ele[6][8];
    ele[5][8] != ele[7][8];
    ele[5][8] != ele[8][8];
    ele[6][0] != ele[6][1];
    ele[6][0] != ele[6][2];
    ele[6][0] != ele[6][3];
    ele[6][0] != ele[6][4];
    ele[6][0] != ele[6][5];
    ele[6][0] != ele[6][6];
    ele[6][0] != ele[6][7];
    ele[6][0] != ele[6][8];
    ele[6][0] != ele[7][0];
    ele[6][0] != ele[7][1];
    ele[6][0] != ele[7][2];
    ele[6][0] != ele[8][0];
    ele[6][0] != ele[8][1];
    ele[6][0] != ele[8][2];
    ele[6][1] != ele[6][2];
    ele[6][1] != ele[6][3];
    ele[6][1] != ele[6][4];
    ele[6][1] != ele[6][5];
    ele[6][1] != ele[6][6];
    ele[6][1] != ele[6][7];
    ele[6][1] != ele[6][8];
    ele[6][1] != ele[7][0];
    ele[6][1] != ele[7][1];
    ele[6][1] != ele[7][2];
    ele[6][1] != ele[8][0];
    ele[6][1] != ele[8][1];
    ele[6][1] != ele[8][2];
    ele[6][2] != ele[6][3];
    ele[6][2] != ele[6][4];
    ele[6][2] != ele[6][5];
    ele[6][2] != ele[6][6];
    ele[6][2] != ele[6][7];
    ele[6][2] != ele[6][8];
    ele[6][2] != ele[7][0];
    ele[6][2] != ele[7][1];
    ele[6][2] != ele[7][2];
    ele[6][2] != ele[8][0];
    ele[6][2] != ele[8][1];
    ele[6][2] != ele[8][2];
    ele[6][3] != ele[6][4];
    ele[6][3] != ele[6][5];
    ele[6][3] != ele[6][6];
    ele[6][3] != ele[6][7];
    ele[6][3] != ele[6][8];
    ele[6][3] != ele[7][3];
    ele[6][3] != ele[7][4];
    ele[6][3] != ele[7][5];
    ele[6][3] != ele[8][3];
    ele[6][3] != ele[8][4];
    ele[6][3] != ele[8][5];
    ele[6][4] != ele[6][5];
    ele[6][4] != ele[6][6];
    ele[6][4] != ele[6][7];
    ele[6][4] != ele[6][8];
    ele[6][4] != ele[7][3];
    ele[6][4] != ele[7][4];
    ele[6][4] != ele[7][5];
    ele[6][4] != ele[8][3];
    ele[6][4] != ele[8][4];
    ele[6][4] != ele[8][5];
    ele[6][5] != ele[6][6];
    ele[6][5] != ele[6][7];
    ele[6][5] != ele[6][8];
    ele[6][5] != ele[7][3];
    ele[6][5] != ele[7][4];
    ele[6][5] != ele[7][5];
    ele[6][5] != ele[8][3];
    ele[6][5] != ele[8][4];
    ele[6][5] != ele[8][5];
    ele[6][6] != ele[6][7];
    ele[6][6] != ele[6][8];
    ele[6][6] != ele[7][6];
    ele[6][6] != ele[7][7];
    ele[6][6] != ele[7][8];
    ele[6][6] != ele[8][6];
    ele[6][6] != ele[8][7];
    ele[6][6] != ele[8][8];
    ele[6][7] != ele[6][8];
    ele[6][7] != ele[7][6];
    ele[6][7] != ele[7][7];
    ele[6][7] != ele[7][8];
    ele[6][7] != ele[8][6];
    ele[6][7] != ele[8][7];
    ele[6][7] != ele[8][8];
    ele[6][8] != ele[7][6];
    ele[6][8] != ele[7][7];
    ele[6][8] != ele[7][8];
    ele[6][8] != ele[8][6];
    ele[6][8] != ele[8][7];
    ele[6][8] != ele[8][8];
    ele[7][0] != ele[7][1];
    ele[7][0] != ele[7][2];
    ele[7][0] != ele[7][3];
    ele[7][0] != ele[7][4];
    ele[7][0] != ele[7][5];
    ele[7][0] != ele[7][6];
    ele[7][0] != ele[7][7];
    ele[7][0] != ele[7][8];
    ele[7][0] != ele[8][0];
    ele[7][0] != ele[8][1];
    ele[7][0] != ele[8][2];
    ele[7][1] != ele[7][2];
    ele[7][1] != ele[7][3];
    ele[7][1] != ele[7][4];
    ele[7][1] != ele[7][5];
    ele[7][1] != ele[7][6];
    ele[7][1] != ele[7][7];
    ele[7][1] != ele[7][8];
    ele[7][1] != ele[8][0];
    ele[7][1] != ele[8][1];
    ele[7][1] != ele[8][2];
    ele[7][2] != ele[7][3];
    ele[7][2] != ele[7][4];
    ele[7][2] != ele[7][5];
    ele[7][2] != ele[7][6];
    ele[7][2] != ele[7][7];
    ele[7][2] != ele[7][8];
    ele[7][2] != ele[8][0];
    ele[7][2] != ele[8][1];
    ele[7][2] != ele[8][2];
    ele[7][3] != ele[7][4];
    ele[7][3] != ele[7][5];
    ele[7][3] != ele[7][6];
    ele[7][3] != ele[7][7];
    ele[7][3] != ele[7][8];
    ele[7][3] != ele[8][3];
    ele[7][3] != ele[8][4];
    ele[7][3] != ele[8][5];
    ele[7][4] != ele[7][5];
    ele[7][4] != ele[7][6];
    ele[7][4] != ele[7][7];
    ele[7][4] != ele[7][8];
    ele[7][4] != ele[8][3];
    ele[7][4] != ele[8][4];
    ele[7][4] != ele[8][5];
    ele[7][5] != ele[7][6];
    ele[7][5] != ele[7][7];
    ele[7][5] != ele[7][8];
    ele[7][5] != ele[8][3];
    ele[7][5] != ele[8][4];
    ele[7][5] != ele[8][5];
    ele[7][6] != ele[7][7];
    ele[7][6] != ele[7][8];
    ele[7][6] != ele[8][6];
    ele[7][6] != ele[8][7];
    ele[7][6] != ele[8][8];
    ele[7][7] != ele[7][8];
    ele[7][7] != ele[8][6];
    ele[7][7] != ele[8][7];
    ele[7][7] != ele[8][8];
    ele[7][8] != ele[8][6];
    ele[7][8] != ele[8][7];
    ele[7][8] != ele[8][8];
    ele[8][0] != ele[8][1];
    ele[8][0] != ele[8][2];
    ele[8][0] != ele[8][3];
    ele[8][0] != ele[8][4];
    ele[8][0] != ele[8][5];
    ele[8][0] != ele[8][6];
    ele[8][0] != ele[8][7];
    ele[8][0] != ele[8][8];
    ele[8][1] != ele[8][2];
    ele[8][1] != ele[8][3];
    ele[8][1] != ele[8][4];
    ele[8][1] != ele[8][5];
    ele[8][1] != ele[8][6];
    ele[8][1] != ele[8][7];
    ele[8][1] != ele[8][8];
    ele[8][2] != ele[8][3];
    ele[8][2] != ele[8][4];
    ele[8][2] != ele[8][5];
    ele[8][2] != ele[8][6];
    ele[8][2] != ele[8][7];
    ele[8][2] != ele[8][8];
    ele[8][3] != ele[8][4];
    ele[8][3] != ele[8][5];
    ele[8][3] != ele[8][6];
    ele[8][3] != ele[8][7];
    ele[8][3] != ele[8][8];
    ele[8][4] != ele[8][5];
    ele[8][4] != ele[8][6];
    ele[8][4] != ele[8][7];
    ele[8][4] != ele[8][8];
    ele[8][5] != ele[8][6];
    ele[8][5] != ele[8][7];
    ele[8][5] != ele[8][8];
    ele[8][6] != ele[8][7];
    ele[8][6] != ele[8][8];
    ele[8][7] != ele[8][8];
  // NUMBER OF CONSTRAINTS: 810
  }
  function new ();
    if (! this.randomize ()) begin
      $display ("ERROR: Randomization failed...!!!");
    end
  endfunction: new
  function show ();
    $display (ele[0][0], ele[0][1], ele[0][2], ele[0][3], ele[0][4], ele[0][5], ele[0][6], ele[0][7], ele[0][8]);
    $display (ele[1][0], ele[1][1], ele[1][2], ele[1][3], ele[1][4], ele[1][5], ele[1][6], ele[1][7], ele[1][8]);
    $display (ele[2][0], ele[2][1], ele[2][2], ele[2][3], ele[2][4], ele[2][5], ele[2][6], ele[2][7], ele[2][8]);
    $display (ele[3][0], ele[3][1], ele[3][2], ele[3][3], ele[3][4], ele[3][5], ele[3][6], ele[3][7], ele[3][8]);
    $display (ele[4][0], ele[4][1], ele[4][2], ele[4][3], ele[4][4], ele[4][5], ele[4][6], ele[4][7], ele[4][8]);
    $display (ele[5][0], ele[5][1], ele[5][2], ele[5][3], ele[5][4], ele[5][5], ele[5][6], ele[5][7], ele[5][8]);
    $display (ele[6][0], ele[6][1], ele[6][2], ele[6][3], ele[6][4], ele[6][5], ele[6][6], ele[6][7], ele[6][8]);
    $display (ele[7][0], ele[7][1], ele[7][2], ele[7][3], ele[7][4], ele[7][5], ele[7][6], ele[7][7], ele[7][8]);
    $display (ele[8][0], ele[8][1], ele[8][2], ele[8][3], ele[8][4], ele[8][5], ele[8][6], ele[8][7], ele[8][8]);
  endfunction: show
endclass: board
