program core (
        input clk,
        input rst, 
        core_cache_if.core_p cache_if
);


endprogram
