module cache (input clk, input rst, core_cache_if.cache_p core_if);

endmodule
