class board;
  typedef enum {
    AAA=1,
    AAB=2,
    AAC=3,
    AAD=4,
    AAE=5,
    AAF=6,
    AAG=7,
    AAH=8,
    AAI=9,
    AAJ=10,
    AAK=11,
    AAL=12,
    AAM=13,
    AAN=14,
    AAO=15,
    AAP
  } elements;
  rand elements ele[16][16];
  constraint all {
    ele[0][0] != ele[0][1];
    ele[0][0] != ele[0][10];
    ele[0][0] != ele[0][11];
    ele[0][0] != ele[0][12];
    ele[0][0] != ele[0][13];
    ele[0][0] != ele[0][14];
    ele[0][0] != ele[0][15];
    ele[0][0] != ele[0][2];
    ele[0][0] != ele[0][3];
    ele[0][0] != ele[0][4];
    ele[0][0] != ele[0][5];
    ele[0][0] != ele[0][6];
    ele[0][0] != ele[0][7];
    ele[0][0] != ele[0][8];
    ele[0][0] != ele[0][9];
    ele[0][0] != ele[1][0];
    ele[0][0] != ele[1][1];
    ele[0][0] != ele[1][2];
    ele[0][0] != ele[1][3];
    ele[0][0] != ele[10][0];
    ele[0][0] != ele[11][0];
    ele[0][0] != ele[12][0];
    ele[0][0] != ele[13][0];
    ele[0][0] != ele[14][0];
    ele[0][0] != ele[15][0];
    ele[0][0] != ele[2][0];
    ele[0][0] != ele[2][1];
    ele[0][0] != ele[2][2];
    ele[0][0] != ele[2][3];
    ele[0][0] != ele[3][0];
    ele[0][0] != ele[3][1];
    ele[0][0] != ele[3][2];
    ele[0][0] != ele[3][3];
    ele[0][0] != ele[4][0];
    ele[0][0] != ele[5][0];
    ele[0][0] != ele[6][0];
    ele[0][0] != ele[7][0];
    ele[0][0] != ele[8][0];
    ele[0][0] != ele[9][0];
    ele[0][1] != ele[0][10];
    ele[0][1] != ele[0][11];
    ele[0][1] != ele[0][12];
    ele[0][1] != ele[0][13];
    ele[0][1] != ele[0][14];
    ele[0][1] != ele[0][15];
    ele[0][1] != ele[0][2];
    ele[0][1] != ele[0][3];
    ele[0][1] != ele[0][4];
    ele[0][1] != ele[0][5];
    ele[0][1] != ele[0][6];
    ele[0][1] != ele[0][7];
    ele[0][1] != ele[0][8];
    ele[0][1] != ele[0][9];
    ele[0][1] != ele[1][0];
    ele[0][1] != ele[1][1];
    ele[0][1] != ele[1][2];
    ele[0][1] != ele[1][3];
    ele[0][1] != ele[10][1];
    ele[0][1] != ele[11][1];
    ele[0][1] != ele[12][1];
    ele[0][1] != ele[13][1];
    ele[0][1] != ele[14][1];
    ele[0][1] != ele[15][1];
    ele[0][1] != ele[2][0];
    ele[0][1] != ele[2][1];
    ele[0][1] != ele[2][2];
    ele[0][1] != ele[2][3];
    ele[0][1] != ele[3][0];
    ele[0][1] != ele[3][1];
    ele[0][1] != ele[3][2];
    ele[0][1] != ele[3][3];
    ele[0][1] != ele[4][1];
    ele[0][1] != ele[5][1];
    ele[0][1] != ele[6][1];
    ele[0][1] != ele[7][1];
    ele[0][1] != ele[8][1];
    ele[0][1] != ele[9][1];
    ele[0][10] != ele[0][11];
    ele[0][10] != ele[0][12];
    ele[0][10] != ele[0][13];
    ele[0][10] != ele[0][14];
    ele[0][10] != ele[0][15];
    ele[0][10] != ele[1][10];
    ele[0][10] != ele[1][11];
    ele[0][10] != ele[1][8];
    ele[0][10] != ele[1][9];
    ele[0][10] != ele[10][10];
    ele[0][10] != ele[11][10];
    ele[0][10] != ele[12][10];
    ele[0][10] != ele[13][10];
    ele[0][10] != ele[14][10];
    ele[0][10] != ele[15][10];
    ele[0][10] != ele[2][10];
    ele[0][10] != ele[2][11];
    ele[0][10] != ele[2][8];
    ele[0][10] != ele[2][9];
    ele[0][10] != ele[3][10];
    ele[0][10] != ele[3][11];
    ele[0][10] != ele[3][8];
    ele[0][10] != ele[3][9];
    ele[0][10] != ele[4][10];
    ele[0][10] != ele[5][10];
    ele[0][10] != ele[6][10];
    ele[0][10] != ele[7][10];
    ele[0][10] != ele[8][10];
    ele[0][10] != ele[9][10];
    ele[0][11] != ele[0][12];
    ele[0][11] != ele[0][13];
    ele[0][11] != ele[0][14];
    ele[0][11] != ele[0][15];
    ele[0][11] != ele[1][10];
    ele[0][11] != ele[1][11];
    ele[0][11] != ele[1][8];
    ele[0][11] != ele[1][9];
    ele[0][11] != ele[10][11];
    ele[0][11] != ele[11][11];
    ele[0][11] != ele[12][11];
    ele[0][11] != ele[13][11];
    ele[0][11] != ele[14][11];
    ele[0][11] != ele[15][11];
    ele[0][11] != ele[2][10];
    ele[0][11] != ele[2][11];
    ele[0][11] != ele[2][8];
    ele[0][11] != ele[2][9];
    ele[0][11] != ele[3][10];
    ele[0][11] != ele[3][11];
    ele[0][11] != ele[3][8];
    ele[0][11] != ele[3][9];
    ele[0][11] != ele[4][11];
    ele[0][11] != ele[5][11];
    ele[0][11] != ele[6][11];
    ele[0][11] != ele[7][11];
    ele[0][11] != ele[8][11];
    ele[0][11] != ele[9][11];
    ele[0][12] != ele[0][13];
    ele[0][12] != ele[0][14];
    ele[0][12] != ele[0][15];
    ele[0][12] != ele[1][12];
    ele[0][12] != ele[1][13];
    ele[0][12] != ele[1][14];
    ele[0][12] != ele[1][15];
    ele[0][12] != ele[10][12];
    ele[0][12] != ele[11][12];
    ele[0][12] != ele[12][12];
    ele[0][12] != ele[13][12];
    ele[0][12] != ele[14][12];
    ele[0][12] != ele[15][12];
    ele[0][12] != ele[2][12];
    ele[0][12] != ele[2][13];
    ele[0][12] != ele[2][14];
    ele[0][12] != ele[2][15];
    ele[0][12] != ele[3][12];
    ele[0][12] != ele[3][13];
    ele[0][12] != ele[3][14];
    ele[0][12] != ele[3][15];
    ele[0][12] != ele[4][12];
    ele[0][12] != ele[5][12];
    ele[0][12] != ele[6][12];
    ele[0][12] != ele[7][12];
    ele[0][12] != ele[8][12];
    ele[0][12] != ele[9][12];
    ele[0][13] != ele[0][14];
    ele[0][13] != ele[0][15];
    ele[0][13] != ele[1][12];
    ele[0][13] != ele[1][13];
    ele[0][13] != ele[1][14];
    ele[0][13] != ele[1][15];
    ele[0][13] != ele[10][13];
    ele[0][13] != ele[11][13];
    ele[0][13] != ele[12][13];
    ele[0][13] != ele[13][13];
    ele[0][13] != ele[14][13];
    ele[0][13] != ele[15][13];
    ele[0][13] != ele[2][12];
    ele[0][13] != ele[2][13];
    ele[0][13] != ele[2][14];
    ele[0][13] != ele[2][15];
    ele[0][13] != ele[3][12];
    ele[0][13] != ele[3][13];
    ele[0][13] != ele[3][14];
    ele[0][13] != ele[3][15];
    ele[0][13] != ele[4][13];
    ele[0][13] != ele[5][13];
    ele[0][13] != ele[6][13];
    ele[0][13] != ele[7][13];
    ele[0][13] != ele[8][13];
    ele[0][13] != ele[9][13];
    ele[0][14] != ele[0][15];
    ele[0][14] != ele[1][12];
    ele[0][14] != ele[1][13];
    ele[0][14] != ele[1][14];
    ele[0][14] != ele[1][15];
    ele[0][14] != ele[10][14];
    ele[0][14] != ele[11][14];
    ele[0][14] != ele[12][14];
    ele[0][14] != ele[13][14];
    ele[0][14] != ele[14][14];
    ele[0][14] != ele[15][14];
    ele[0][14] != ele[2][12];
    ele[0][14] != ele[2][13];
    ele[0][14] != ele[2][14];
    ele[0][14] != ele[2][15];
    ele[0][14] != ele[3][12];
    ele[0][14] != ele[3][13];
    ele[0][14] != ele[3][14];
    ele[0][14] != ele[3][15];
    ele[0][14] != ele[4][14];
    ele[0][14] != ele[5][14];
    ele[0][14] != ele[6][14];
    ele[0][14] != ele[7][14];
    ele[0][14] != ele[8][14];
    ele[0][14] != ele[9][14];
    ele[0][15] != ele[1][12];
    ele[0][15] != ele[1][13];
    ele[0][15] != ele[1][14];
    ele[0][15] != ele[1][15];
    ele[0][15] != ele[10][15];
    ele[0][15] != ele[11][15];
    ele[0][15] != ele[12][15];
    ele[0][15] != ele[13][15];
    ele[0][15] != ele[14][15];
    ele[0][15] != ele[15][15];
    ele[0][15] != ele[2][12];
    ele[0][15] != ele[2][13];
    ele[0][15] != ele[2][14];
    ele[0][15] != ele[2][15];
    ele[0][15] != ele[3][12];
    ele[0][15] != ele[3][13];
    ele[0][15] != ele[3][14];
    ele[0][15] != ele[3][15];
    ele[0][15] != ele[4][15];
    ele[0][15] != ele[5][15];
    ele[0][15] != ele[6][15];
    ele[0][15] != ele[7][15];
    ele[0][15] != ele[8][15];
    ele[0][15] != ele[9][15];
    ele[0][2] != ele[0][10];
    ele[0][2] != ele[0][11];
    ele[0][2] != ele[0][12];
    ele[0][2] != ele[0][13];
    ele[0][2] != ele[0][14];
    ele[0][2] != ele[0][15];
    ele[0][2] != ele[0][3];
    ele[0][2] != ele[0][4];
    ele[0][2] != ele[0][5];
    ele[0][2] != ele[0][6];
    ele[0][2] != ele[0][7];
    ele[0][2] != ele[0][8];
    ele[0][2] != ele[0][9];
    ele[0][2] != ele[1][0];
    ele[0][2] != ele[1][1];
    ele[0][2] != ele[1][2];
    ele[0][2] != ele[1][3];
    ele[0][2] != ele[10][2];
    ele[0][2] != ele[11][2];
    ele[0][2] != ele[12][2];
    ele[0][2] != ele[13][2];
    ele[0][2] != ele[14][2];
    ele[0][2] != ele[15][2];
    ele[0][2] != ele[2][0];
    ele[0][2] != ele[2][1];
    ele[0][2] != ele[2][2];
    ele[0][2] != ele[2][3];
    ele[0][2] != ele[3][0];
    ele[0][2] != ele[3][1];
    ele[0][2] != ele[3][2];
    ele[0][2] != ele[3][3];
    ele[0][2] != ele[4][2];
    ele[0][2] != ele[5][2];
    ele[0][2] != ele[6][2];
    ele[0][2] != ele[7][2];
    ele[0][2] != ele[8][2];
    ele[0][2] != ele[9][2];
    ele[0][3] != ele[0][10];
    ele[0][3] != ele[0][11];
    ele[0][3] != ele[0][12];
    ele[0][3] != ele[0][13];
    ele[0][3] != ele[0][14];
    ele[0][3] != ele[0][15];
    ele[0][3] != ele[0][4];
    ele[0][3] != ele[0][5];
    ele[0][3] != ele[0][6];
    ele[0][3] != ele[0][7];
    ele[0][3] != ele[0][8];
    ele[0][3] != ele[0][9];
    ele[0][3] != ele[1][0];
    ele[0][3] != ele[1][1];
    ele[0][3] != ele[1][2];
    ele[0][3] != ele[1][3];
    ele[0][3] != ele[10][3];
    ele[0][3] != ele[11][3];
    ele[0][3] != ele[12][3];
    ele[0][3] != ele[13][3];
    ele[0][3] != ele[14][3];
    ele[0][3] != ele[15][3];
    ele[0][3] != ele[2][0];
    ele[0][3] != ele[2][1];
    ele[0][3] != ele[2][2];
    ele[0][3] != ele[2][3];
    ele[0][3] != ele[3][0];
    ele[0][3] != ele[3][1];
    ele[0][3] != ele[3][2];
    ele[0][3] != ele[3][3];
    ele[0][3] != ele[4][3];
    ele[0][3] != ele[5][3];
    ele[0][3] != ele[6][3];
    ele[0][3] != ele[7][3];
    ele[0][3] != ele[8][3];
    ele[0][3] != ele[9][3];
    ele[0][4] != ele[0][10];
    ele[0][4] != ele[0][11];
    ele[0][4] != ele[0][12];
    ele[0][4] != ele[0][13];
    ele[0][4] != ele[0][14];
    ele[0][4] != ele[0][15];
    ele[0][4] != ele[0][5];
    ele[0][4] != ele[0][6];
    ele[0][4] != ele[0][7];
    ele[0][4] != ele[0][8];
    ele[0][4] != ele[0][9];
    ele[0][4] != ele[1][4];
    ele[0][4] != ele[1][5];
    ele[0][4] != ele[1][6];
    ele[0][4] != ele[1][7];
    ele[0][4] != ele[10][4];
    ele[0][4] != ele[11][4];
    ele[0][4] != ele[12][4];
    ele[0][4] != ele[13][4];
    ele[0][4] != ele[14][4];
    ele[0][4] != ele[15][4];
    ele[0][4] != ele[2][4];
    ele[0][4] != ele[2][5];
    ele[0][4] != ele[2][6];
    ele[0][4] != ele[2][7];
    ele[0][4] != ele[3][4];
    ele[0][4] != ele[3][5];
    ele[0][4] != ele[3][6];
    ele[0][4] != ele[3][7];
    ele[0][4] != ele[4][4];
    ele[0][4] != ele[5][4];
    ele[0][4] != ele[6][4];
    ele[0][4] != ele[7][4];
    ele[0][4] != ele[8][4];
    ele[0][4] != ele[9][4];
    ele[0][5] != ele[0][10];
    ele[0][5] != ele[0][11];
    ele[0][5] != ele[0][12];
    ele[0][5] != ele[0][13];
    ele[0][5] != ele[0][14];
    ele[0][5] != ele[0][15];
    ele[0][5] != ele[0][6];
    ele[0][5] != ele[0][7];
    ele[0][5] != ele[0][8];
    ele[0][5] != ele[0][9];
    ele[0][5] != ele[1][4];
    ele[0][5] != ele[1][5];
    ele[0][5] != ele[1][6];
    ele[0][5] != ele[1][7];
    ele[0][5] != ele[10][5];
    ele[0][5] != ele[11][5];
    ele[0][5] != ele[12][5];
    ele[0][5] != ele[13][5];
    ele[0][5] != ele[14][5];
    ele[0][5] != ele[15][5];
    ele[0][5] != ele[2][4];
    ele[0][5] != ele[2][5];
    ele[0][5] != ele[2][6];
    ele[0][5] != ele[2][7];
    ele[0][5] != ele[3][4];
    ele[0][5] != ele[3][5];
    ele[0][5] != ele[3][6];
    ele[0][5] != ele[3][7];
    ele[0][5] != ele[4][5];
    ele[0][5] != ele[5][5];
    ele[0][5] != ele[6][5];
    ele[0][5] != ele[7][5];
    ele[0][5] != ele[8][5];
    ele[0][5] != ele[9][5];
    ele[0][6] != ele[0][10];
    ele[0][6] != ele[0][11];
    ele[0][6] != ele[0][12];
    ele[0][6] != ele[0][13];
    ele[0][6] != ele[0][14];
    ele[0][6] != ele[0][15];
    ele[0][6] != ele[0][7];
    ele[0][6] != ele[0][8];
    ele[0][6] != ele[0][9];
    ele[0][6] != ele[1][4];
    ele[0][6] != ele[1][5];
    ele[0][6] != ele[1][6];
    ele[0][6] != ele[1][7];
    ele[0][6] != ele[10][6];
    ele[0][6] != ele[11][6];
    ele[0][6] != ele[12][6];
    ele[0][6] != ele[13][6];
    ele[0][6] != ele[14][6];
    ele[0][6] != ele[15][6];
    ele[0][6] != ele[2][4];
    ele[0][6] != ele[2][5];
    ele[0][6] != ele[2][6];
    ele[0][6] != ele[2][7];
    ele[0][6] != ele[3][4];
    ele[0][6] != ele[3][5];
    ele[0][6] != ele[3][6];
    ele[0][6] != ele[3][7];
    ele[0][6] != ele[4][6];
    ele[0][6] != ele[5][6];
    ele[0][6] != ele[6][6];
    ele[0][6] != ele[7][6];
    ele[0][6] != ele[8][6];
    ele[0][6] != ele[9][6];
    ele[0][7] != ele[0][10];
    ele[0][7] != ele[0][11];
    ele[0][7] != ele[0][12];
    ele[0][7] != ele[0][13];
    ele[0][7] != ele[0][14];
    ele[0][7] != ele[0][15];
    ele[0][7] != ele[0][8];
    ele[0][7] != ele[0][9];
    ele[0][7] != ele[1][4];
    ele[0][7] != ele[1][5];
    ele[0][7] != ele[1][6];
    ele[0][7] != ele[1][7];
    ele[0][7] != ele[10][7];
    ele[0][7] != ele[11][7];
    ele[0][7] != ele[12][7];
    ele[0][7] != ele[13][7];
    ele[0][7] != ele[14][7];
    ele[0][7] != ele[15][7];
    ele[0][7] != ele[2][4];
    ele[0][7] != ele[2][5];
    ele[0][7] != ele[2][6];
    ele[0][7] != ele[2][7];
    ele[0][7] != ele[3][4];
    ele[0][7] != ele[3][5];
    ele[0][7] != ele[3][6];
    ele[0][7] != ele[3][7];
    ele[0][7] != ele[4][7];
    ele[0][7] != ele[5][7];
    ele[0][7] != ele[6][7];
    ele[0][7] != ele[7][7];
    ele[0][7] != ele[8][7];
    ele[0][7] != ele[9][7];
    ele[0][8] != ele[0][10];
    ele[0][8] != ele[0][11];
    ele[0][8] != ele[0][12];
    ele[0][8] != ele[0][13];
    ele[0][8] != ele[0][14];
    ele[0][8] != ele[0][15];
    ele[0][8] != ele[0][9];
    ele[0][8] != ele[1][10];
    ele[0][8] != ele[1][11];
    ele[0][8] != ele[1][8];
    ele[0][8] != ele[1][9];
    ele[0][8] != ele[10][8];
    ele[0][8] != ele[11][8];
    ele[0][8] != ele[12][8];
    ele[0][8] != ele[13][8];
    ele[0][8] != ele[14][8];
    ele[0][8] != ele[15][8];
    ele[0][8] != ele[2][10];
    ele[0][8] != ele[2][11];
    ele[0][8] != ele[2][8];
    ele[0][8] != ele[2][9];
    ele[0][8] != ele[3][10];
    ele[0][8] != ele[3][11];
    ele[0][8] != ele[3][8];
    ele[0][8] != ele[3][9];
    ele[0][8] != ele[4][8];
    ele[0][8] != ele[5][8];
    ele[0][8] != ele[6][8];
    ele[0][8] != ele[7][8];
    ele[0][8] != ele[8][8];
    ele[0][8] != ele[9][8];
    ele[0][9] != ele[0][10];
    ele[0][9] != ele[0][11];
    ele[0][9] != ele[0][12];
    ele[0][9] != ele[0][13];
    ele[0][9] != ele[0][14];
    ele[0][9] != ele[0][15];
    ele[0][9] != ele[1][10];
    ele[0][9] != ele[1][11];
    ele[0][9] != ele[1][8];
    ele[0][9] != ele[1][9];
    ele[0][9] != ele[10][9];
    ele[0][9] != ele[11][9];
    ele[0][9] != ele[12][9];
    ele[0][9] != ele[13][9];
    ele[0][9] != ele[14][9];
    ele[0][9] != ele[15][9];
    ele[0][9] != ele[2][10];
    ele[0][9] != ele[2][11];
    ele[0][9] != ele[2][8];
    ele[0][9] != ele[2][9];
    ele[0][9] != ele[3][10];
    ele[0][9] != ele[3][11];
    ele[0][9] != ele[3][8];
    ele[0][9] != ele[3][9];
    ele[0][9] != ele[4][9];
    ele[0][9] != ele[5][9];
    ele[0][9] != ele[6][9];
    ele[0][9] != ele[7][9];
    ele[0][9] != ele[8][9];
    ele[0][9] != ele[9][9];
    ele[1][0] != ele[1][1];
    ele[1][0] != ele[1][10];
    ele[1][0] != ele[1][11];
    ele[1][0] != ele[1][12];
    ele[1][0] != ele[1][13];
    ele[1][0] != ele[1][14];
    ele[1][0] != ele[1][15];
    ele[1][0] != ele[1][2];
    ele[1][0] != ele[1][3];
    ele[1][0] != ele[1][4];
    ele[1][0] != ele[1][5];
    ele[1][0] != ele[1][6];
    ele[1][0] != ele[1][7];
    ele[1][0] != ele[1][8];
    ele[1][0] != ele[1][9];
    ele[1][0] != ele[10][0];
    ele[1][0] != ele[11][0];
    ele[1][0] != ele[12][0];
    ele[1][0] != ele[13][0];
    ele[1][0] != ele[14][0];
    ele[1][0] != ele[15][0];
    ele[1][0] != ele[2][0];
    ele[1][0] != ele[2][1];
    ele[1][0] != ele[2][2];
    ele[1][0] != ele[2][3];
    ele[1][0] != ele[3][0];
    ele[1][0] != ele[3][1];
    ele[1][0] != ele[3][2];
    ele[1][0] != ele[3][3];
    ele[1][0] != ele[4][0];
    ele[1][0] != ele[5][0];
    ele[1][0] != ele[6][0];
    ele[1][0] != ele[7][0];
    ele[1][0] != ele[8][0];
    ele[1][0] != ele[9][0];
    ele[1][1] != ele[1][10];
    ele[1][1] != ele[1][11];
    ele[1][1] != ele[1][12];
    ele[1][1] != ele[1][13];
    ele[1][1] != ele[1][14];
    ele[1][1] != ele[1][15];
    ele[1][1] != ele[1][2];
    ele[1][1] != ele[1][3];
    ele[1][1] != ele[1][4];
    ele[1][1] != ele[1][5];
    ele[1][1] != ele[1][6];
    ele[1][1] != ele[1][7];
    ele[1][1] != ele[1][8];
    ele[1][1] != ele[1][9];
    ele[1][1] != ele[10][1];
    ele[1][1] != ele[11][1];
    ele[1][1] != ele[12][1];
    ele[1][1] != ele[13][1];
    ele[1][1] != ele[14][1];
    ele[1][1] != ele[15][1];
    ele[1][1] != ele[2][0];
    ele[1][1] != ele[2][1];
    ele[1][1] != ele[2][2];
    ele[1][1] != ele[2][3];
    ele[1][1] != ele[3][0];
    ele[1][1] != ele[3][1];
    ele[1][1] != ele[3][2];
    ele[1][1] != ele[3][3];
    ele[1][1] != ele[4][1];
    ele[1][1] != ele[5][1];
    ele[1][1] != ele[6][1];
    ele[1][1] != ele[7][1];
    ele[1][1] != ele[8][1];
    ele[1][1] != ele[9][1];
    ele[1][10] != ele[1][11];
    ele[1][10] != ele[1][12];
    ele[1][10] != ele[1][13];
    ele[1][10] != ele[1][14];
    ele[1][10] != ele[1][15];
    ele[1][10] != ele[10][10];
    ele[1][10] != ele[11][10];
    ele[1][10] != ele[12][10];
    ele[1][10] != ele[13][10];
    ele[1][10] != ele[14][10];
    ele[1][10] != ele[15][10];
    ele[1][10] != ele[2][10];
    ele[1][10] != ele[2][11];
    ele[1][10] != ele[2][8];
    ele[1][10] != ele[2][9];
    ele[1][10] != ele[3][10];
    ele[1][10] != ele[3][11];
    ele[1][10] != ele[3][8];
    ele[1][10] != ele[3][9];
    ele[1][10] != ele[4][10];
    ele[1][10] != ele[5][10];
    ele[1][10] != ele[6][10];
    ele[1][10] != ele[7][10];
    ele[1][10] != ele[8][10];
    ele[1][10] != ele[9][10];
    ele[1][11] != ele[1][12];
    ele[1][11] != ele[1][13];
    ele[1][11] != ele[1][14];
    ele[1][11] != ele[1][15];
    ele[1][11] != ele[10][11];
    ele[1][11] != ele[11][11];
    ele[1][11] != ele[12][11];
    ele[1][11] != ele[13][11];
    ele[1][11] != ele[14][11];
    ele[1][11] != ele[15][11];
    ele[1][11] != ele[2][10];
    ele[1][11] != ele[2][11];
    ele[1][11] != ele[2][8];
    ele[1][11] != ele[2][9];
    ele[1][11] != ele[3][10];
    ele[1][11] != ele[3][11];
    ele[1][11] != ele[3][8];
    ele[1][11] != ele[3][9];
    ele[1][11] != ele[4][11];
    ele[1][11] != ele[5][11];
    ele[1][11] != ele[6][11];
    ele[1][11] != ele[7][11];
    ele[1][11] != ele[8][11];
    ele[1][11] != ele[9][11];
    ele[1][12] != ele[1][13];
    ele[1][12] != ele[1][14];
    ele[1][12] != ele[1][15];
    ele[1][12] != ele[10][12];
    ele[1][12] != ele[11][12];
    ele[1][12] != ele[12][12];
    ele[1][12] != ele[13][12];
    ele[1][12] != ele[14][12];
    ele[1][12] != ele[15][12];
    ele[1][12] != ele[2][12];
    ele[1][12] != ele[2][13];
    ele[1][12] != ele[2][14];
    ele[1][12] != ele[2][15];
    ele[1][12] != ele[3][12];
    ele[1][12] != ele[3][13];
    ele[1][12] != ele[3][14];
    ele[1][12] != ele[3][15];
    ele[1][12] != ele[4][12];
    ele[1][12] != ele[5][12];
    ele[1][12] != ele[6][12];
    ele[1][12] != ele[7][12];
    ele[1][12] != ele[8][12];
    ele[1][12] != ele[9][12];
    ele[1][13] != ele[1][14];
    ele[1][13] != ele[1][15];
    ele[1][13] != ele[10][13];
    ele[1][13] != ele[11][13];
    ele[1][13] != ele[12][13];
    ele[1][13] != ele[13][13];
    ele[1][13] != ele[14][13];
    ele[1][13] != ele[15][13];
    ele[1][13] != ele[2][12];
    ele[1][13] != ele[2][13];
    ele[1][13] != ele[2][14];
    ele[1][13] != ele[2][15];
    ele[1][13] != ele[3][12];
    ele[1][13] != ele[3][13];
    ele[1][13] != ele[3][14];
    ele[1][13] != ele[3][15];
    ele[1][13] != ele[4][13];
    ele[1][13] != ele[5][13];
    ele[1][13] != ele[6][13];
    ele[1][13] != ele[7][13];
    ele[1][13] != ele[8][13];
    ele[1][13] != ele[9][13];
    ele[1][14] != ele[1][15];
    ele[1][14] != ele[10][14];
    ele[1][14] != ele[11][14];
    ele[1][14] != ele[12][14];
    ele[1][14] != ele[13][14];
    ele[1][14] != ele[14][14];
    ele[1][14] != ele[15][14];
    ele[1][14] != ele[2][12];
    ele[1][14] != ele[2][13];
    ele[1][14] != ele[2][14];
    ele[1][14] != ele[2][15];
    ele[1][14] != ele[3][12];
    ele[1][14] != ele[3][13];
    ele[1][14] != ele[3][14];
    ele[1][14] != ele[3][15];
    ele[1][14] != ele[4][14];
    ele[1][14] != ele[5][14];
    ele[1][14] != ele[6][14];
    ele[1][14] != ele[7][14];
    ele[1][14] != ele[8][14];
    ele[1][14] != ele[9][14];
    ele[1][15] != ele[10][15];
    ele[1][15] != ele[11][15];
    ele[1][15] != ele[12][15];
    ele[1][15] != ele[13][15];
    ele[1][15] != ele[14][15];
    ele[1][15] != ele[15][15];
    ele[1][15] != ele[2][12];
    ele[1][15] != ele[2][13];
    ele[1][15] != ele[2][14];
    ele[1][15] != ele[2][15];
    ele[1][15] != ele[3][12];
    ele[1][15] != ele[3][13];
    ele[1][15] != ele[3][14];
    ele[1][15] != ele[3][15];
    ele[1][15] != ele[4][15];
    ele[1][15] != ele[5][15];
    ele[1][15] != ele[6][15];
    ele[1][15] != ele[7][15];
    ele[1][15] != ele[8][15];
    ele[1][15] != ele[9][15];
    ele[1][2] != ele[1][10];
    ele[1][2] != ele[1][11];
    ele[1][2] != ele[1][12];
    ele[1][2] != ele[1][13];
    ele[1][2] != ele[1][14];
    ele[1][2] != ele[1][15];
    ele[1][2] != ele[1][3];
    ele[1][2] != ele[1][4];
    ele[1][2] != ele[1][5];
    ele[1][2] != ele[1][6];
    ele[1][2] != ele[1][7];
    ele[1][2] != ele[1][8];
    ele[1][2] != ele[1][9];
    ele[1][2] != ele[10][2];
    ele[1][2] != ele[11][2];
    ele[1][2] != ele[12][2];
    ele[1][2] != ele[13][2];
    ele[1][2] != ele[14][2];
    ele[1][2] != ele[15][2];
    ele[1][2] != ele[2][0];
    ele[1][2] != ele[2][1];
    ele[1][2] != ele[2][2];
    ele[1][2] != ele[2][3];
    ele[1][2] != ele[3][0];
    ele[1][2] != ele[3][1];
    ele[1][2] != ele[3][2];
    ele[1][2] != ele[3][3];
    ele[1][2] != ele[4][2];
    ele[1][2] != ele[5][2];
    ele[1][2] != ele[6][2];
    ele[1][2] != ele[7][2];
    ele[1][2] != ele[8][2];
    ele[1][2] != ele[9][2];
    ele[1][3] != ele[1][10];
    ele[1][3] != ele[1][11];
    ele[1][3] != ele[1][12];
    ele[1][3] != ele[1][13];
    ele[1][3] != ele[1][14];
    ele[1][3] != ele[1][15];
    ele[1][3] != ele[1][4];
    ele[1][3] != ele[1][5];
    ele[1][3] != ele[1][6];
    ele[1][3] != ele[1][7];
    ele[1][3] != ele[1][8];
    ele[1][3] != ele[1][9];
    ele[1][3] != ele[10][3];
    ele[1][3] != ele[11][3];
    ele[1][3] != ele[12][3];
    ele[1][3] != ele[13][3];
    ele[1][3] != ele[14][3];
    ele[1][3] != ele[15][3];
    ele[1][3] != ele[2][0];
    ele[1][3] != ele[2][1];
    ele[1][3] != ele[2][2];
    ele[1][3] != ele[2][3];
    ele[1][3] != ele[3][0];
    ele[1][3] != ele[3][1];
    ele[1][3] != ele[3][2];
    ele[1][3] != ele[3][3];
    ele[1][3] != ele[4][3];
    ele[1][3] != ele[5][3];
    ele[1][3] != ele[6][3];
    ele[1][3] != ele[7][3];
    ele[1][3] != ele[8][3];
    ele[1][3] != ele[9][3];
    ele[1][4] != ele[1][10];
    ele[1][4] != ele[1][11];
    ele[1][4] != ele[1][12];
    ele[1][4] != ele[1][13];
    ele[1][4] != ele[1][14];
    ele[1][4] != ele[1][15];
    ele[1][4] != ele[1][5];
    ele[1][4] != ele[1][6];
    ele[1][4] != ele[1][7];
    ele[1][4] != ele[1][8];
    ele[1][4] != ele[1][9];
    ele[1][4] != ele[10][4];
    ele[1][4] != ele[11][4];
    ele[1][4] != ele[12][4];
    ele[1][4] != ele[13][4];
    ele[1][4] != ele[14][4];
    ele[1][4] != ele[15][4];
    ele[1][4] != ele[2][4];
    ele[1][4] != ele[2][5];
    ele[1][4] != ele[2][6];
    ele[1][4] != ele[2][7];
    ele[1][4] != ele[3][4];
    ele[1][4] != ele[3][5];
    ele[1][4] != ele[3][6];
    ele[1][4] != ele[3][7];
    ele[1][4] != ele[4][4];
    ele[1][4] != ele[5][4];
    ele[1][4] != ele[6][4];
    ele[1][4] != ele[7][4];
    ele[1][4] != ele[8][4];
    ele[1][4] != ele[9][4];
    ele[1][5] != ele[1][10];
    ele[1][5] != ele[1][11];
    ele[1][5] != ele[1][12];
    ele[1][5] != ele[1][13];
    ele[1][5] != ele[1][14];
    ele[1][5] != ele[1][15];
    ele[1][5] != ele[1][6];
    ele[1][5] != ele[1][7];
    ele[1][5] != ele[1][8];
    ele[1][5] != ele[1][9];
    ele[1][5] != ele[10][5];
    ele[1][5] != ele[11][5];
    ele[1][5] != ele[12][5];
    ele[1][5] != ele[13][5];
    ele[1][5] != ele[14][5];
    ele[1][5] != ele[15][5];
    ele[1][5] != ele[2][4];
    ele[1][5] != ele[2][5];
    ele[1][5] != ele[2][6];
    ele[1][5] != ele[2][7];
    ele[1][5] != ele[3][4];
    ele[1][5] != ele[3][5];
    ele[1][5] != ele[3][6];
    ele[1][5] != ele[3][7];
    ele[1][5] != ele[4][5];
    ele[1][5] != ele[5][5];
    ele[1][5] != ele[6][5];
    ele[1][5] != ele[7][5];
    ele[1][5] != ele[8][5];
    ele[1][5] != ele[9][5];
    ele[1][6] != ele[1][10];
    ele[1][6] != ele[1][11];
    ele[1][6] != ele[1][12];
    ele[1][6] != ele[1][13];
    ele[1][6] != ele[1][14];
    ele[1][6] != ele[1][15];
    ele[1][6] != ele[1][7];
    ele[1][6] != ele[1][8];
    ele[1][6] != ele[1][9];
    ele[1][6] != ele[10][6];
    ele[1][6] != ele[11][6];
    ele[1][6] != ele[12][6];
    ele[1][6] != ele[13][6];
    ele[1][6] != ele[14][6];
    ele[1][6] != ele[15][6];
    ele[1][6] != ele[2][4];
    ele[1][6] != ele[2][5];
    ele[1][6] != ele[2][6];
    ele[1][6] != ele[2][7];
    ele[1][6] != ele[3][4];
    ele[1][6] != ele[3][5];
    ele[1][6] != ele[3][6];
    ele[1][6] != ele[3][7];
    ele[1][6] != ele[4][6];
    ele[1][6] != ele[5][6];
    ele[1][6] != ele[6][6];
    ele[1][6] != ele[7][6];
    ele[1][6] != ele[8][6];
    ele[1][6] != ele[9][6];
    ele[1][7] != ele[1][10];
    ele[1][7] != ele[1][11];
    ele[1][7] != ele[1][12];
    ele[1][7] != ele[1][13];
    ele[1][7] != ele[1][14];
    ele[1][7] != ele[1][15];
    ele[1][7] != ele[1][8];
    ele[1][7] != ele[1][9];
    ele[1][7] != ele[10][7];
    ele[1][7] != ele[11][7];
    ele[1][7] != ele[12][7];
    ele[1][7] != ele[13][7];
    ele[1][7] != ele[14][7];
    ele[1][7] != ele[15][7];
    ele[1][7] != ele[2][4];
    ele[1][7] != ele[2][5];
    ele[1][7] != ele[2][6];
    ele[1][7] != ele[2][7];
    ele[1][7] != ele[3][4];
    ele[1][7] != ele[3][5];
    ele[1][7] != ele[3][6];
    ele[1][7] != ele[3][7];
    ele[1][7] != ele[4][7];
    ele[1][7] != ele[5][7];
    ele[1][7] != ele[6][7];
    ele[1][7] != ele[7][7];
    ele[1][7] != ele[8][7];
    ele[1][7] != ele[9][7];
    ele[1][8] != ele[1][10];
    ele[1][8] != ele[1][11];
    ele[1][8] != ele[1][12];
    ele[1][8] != ele[1][13];
    ele[1][8] != ele[1][14];
    ele[1][8] != ele[1][15];
    ele[1][8] != ele[1][9];
    ele[1][8] != ele[10][8];
    ele[1][8] != ele[11][8];
    ele[1][8] != ele[12][8];
    ele[1][8] != ele[13][8];
    ele[1][8] != ele[14][8];
    ele[1][8] != ele[15][8];
    ele[1][8] != ele[2][10];
    ele[1][8] != ele[2][11];
    ele[1][8] != ele[2][8];
    ele[1][8] != ele[2][9];
    ele[1][8] != ele[3][10];
    ele[1][8] != ele[3][11];
    ele[1][8] != ele[3][8];
    ele[1][8] != ele[3][9];
    ele[1][8] != ele[4][8];
    ele[1][8] != ele[5][8];
    ele[1][8] != ele[6][8];
    ele[1][8] != ele[7][8];
    ele[1][8] != ele[8][8];
    ele[1][8] != ele[9][8];
    ele[1][9] != ele[1][10];
    ele[1][9] != ele[1][11];
    ele[1][9] != ele[1][12];
    ele[1][9] != ele[1][13];
    ele[1][9] != ele[1][14];
    ele[1][9] != ele[1][15];
    ele[1][9] != ele[10][9];
    ele[1][9] != ele[11][9];
    ele[1][9] != ele[12][9];
    ele[1][9] != ele[13][9];
    ele[1][9] != ele[14][9];
    ele[1][9] != ele[15][9];
    ele[1][9] != ele[2][10];
    ele[1][9] != ele[2][11];
    ele[1][9] != ele[2][8];
    ele[1][9] != ele[2][9];
    ele[1][9] != ele[3][10];
    ele[1][9] != ele[3][11];
    ele[1][9] != ele[3][8];
    ele[1][9] != ele[3][9];
    ele[1][9] != ele[4][9];
    ele[1][9] != ele[5][9];
    ele[1][9] != ele[6][9];
    ele[1][9] != ele[7][9];
    ele[1][9] != ele[8][9];
    ele[1][9] != ele[9][9];
    ele[10][0] != ele[10][1];
    ele[10][0] != ele[10][10];
    ele[10][0] != ele[10][11];
    ele[10][0] != ele[10][12];
    ele[10][0] != ele[10][13];
    ele[10][0] != ele[10][14];
    ele[10][0] != ele[10][15];
    ele[10][0] != ele[10][2];
    ele[10][0] != ele[10][3];
    ele[10][0] != ele[10][4];
    ele[10][0] != ele[10][5];
    ele[10][0] != ele[10][6];
    ele[10][0] != ele[10][7];
    ele[10][0] != ele[10][8];
    ele[10][0] != ele[10][9];
    ele[10][0] != ele[11][0];
    ele[10][0] != ele[11][1];
    ele[10][0] != ele[11][2];
    ele[10][0] != ele[11][3];
    ele[10][0] != ele[12][0];
    ele[10][0] != ele[13][0];
    ele[10][0] != ele[14][0];
    ele[10][0] != ele[15][0];
    ele[10][1] != ele[10][10];
    ele[10][1] != ele[10][11];
    ele[10][1] != ele[10][12];
    ele[10][1] != ele[10][13];
    ele[10][1] != ele[10][14];
    ele[10][1] != ele[10][15];
    ele[10][1] != ele[10][2];
    ele[10][1] != ele[10][3];
    ele[10][1] != ele[10][4];
    ele[10][1] != ele[10][5];
    ele[10][1] != ele[10][6];
    ele[10][1] != ele[10][7];
    ele[10][1] != ele[10][8];
    ele[10][1] != ele[10][9];
    ele[10][1] != ele[11][0];
    ele[10][1] != ele[11][1];
    ele[10][1] != ele[11][2];
    ele[10][1] != ele[11][3];
    ele[10][1] != ele[12][1];
    ele[10][1] != ele[13][1];
    ele[10][1] != ele[14][1];
    ele[10][1] != ele[15][1];
    ele[10][10] != ele[10][11];
    ele[10][10] != ele[10][12];
    ele[10][10] != ele[10][13];
    ele[10][10] != ele[10][14];
    ele[10][10] != ele[10][15];
    ele[10][10] != ele[11][10];
    ele[10][10] != ele[11][11];
    ele[10][10] != ele[11][8];
    ele[10][10] != ele[11][9];
    ele[10][10] != ele[12][10];
    ele[10][10] != ele[13][10];
    ele[10][10] != ele[14][10];
    ele[10][10] != ele[15][10];
    ele[10][11] != ele[10][12];
    ele[10][11] != ele[10][13];
    ele[10][11] != ele[10][14];
    ele[10][11] != ele[10][15];
    ele[10][11] != ele[11][10];
    ele[10][11] != ele[11][11];
    ele[10][11] != ele[11][8];
    ele[10][11] != ele[11][9];
    ele[10][11] != ele[12][11];
    ele[10][11] != ele[13][11];
    ele[10][11] != ele[14][11];
    ele[10][11] != ele[15][11];
    ele[10][12] != ele[10][13];
    ele[10][12] != ele[10][14];
    ele[10][12] != ele[10][15];
    ele[10][12] != ele[11][12];
    ele[10][12] != ele[11][13];
    ele[10][12] != ele[11][14];
    ele[10][12] != ele[11][15];
    ele[10][12] != ele[12][12];
    ele[10][12] != ele[13][12];
    ele[10][12] != ele[14][12];
    ele[10][12] != ele[15][12];
    ele[10][13] != ele[10][14];
    ele[10][13] != ele[10][15];
    ele[10][13] != ele[11][12];
    ele[10][13] != ele[11][13];
    ele[10][13] != ele[11][14];
    ele[10][13] != ele[11][15];
    ele[10][13] != ele[12][13];
    ele[10][13] != ele[13][13];
    ele[10][13] != ele[14][13];
    ele[10][13] != ele[15][13];
    ele[10][14] != ele[10][15];
    ele[10][14] != ele[11][12];
    ele[10][14] != ele[11][13];
    ele[10][14] != ele[11][14];
    ele[10][14] != ele[11][15];
    ele[10][14] != ele[12][14];
    ele[10][14] != ele[13][14];
    ele[10][14] != ele[14][14];
    ele[10][14] != ele[15][14];
    ele[10][15] != ele[11][12];
    ele[10][15] != ele[11][13];
    ele[10][15] != ele[11][14];
    ele[10][15] != ele[11][15];
    ele[10][15] != ele[12][15];
    ele[10][15] != ele[13][15];
    ele[10][15] != ele[14][15];
    ele[10][15] != ele[15][15];
    ele[10][2] != ele[10][10];
    ele[10][2] != ele[10][11];
    ele[10][2] != ele[10][12];
    ele[10][2] != ele[10][13];
    ele[10][2] != ele[10][14];
    ele[10][2] != ele[10][15];
    ele[10][2] != ele[10][3];
    ele[10][2] != ele[10][4];
    ele[10][2] != ele[10][5];
    ele[10][2] != ele[10][6];
    ele[10][2] != ele[10][7];
    ele[10][2] != ele[10][8];
    ele[10][2] != ele[10][9];
    ele[10][2] != ele[11][0];
    ele[10][2] != ele[11][1];
    ele[10][2] != ele[11][2];
    ele[10][2] != ele[11][3];
    ele[10][2] != ele[12][2];
    ele[10][2] != ele[13][2];
    ele[10][2] != ele[14][2];
    ele[10][2] != ele[15][2];
    ele[10][3] != ele[10][10];
    ele[10][3] != ele[10][11];
    ele[10][3] != ele[10][12];
    ele[10][3] != ele[10][13];
    ele[10][3] != ele[10][14];
    ele[10][3] != ele[10][15];
    ele[10][3] != ele[10][4];
    ele[10][3] != ele[10][5];
    ele[10][3] != ele[10][6];
    ele[10][3] != ele[10][7];
    ele[10][3] != ele[10][8];
    ele[10][3] != ele[10][9];
    ele[10][3] != ele[11][0];
    ele[10][3] != ele[11][1];
    ele[10][3] != ele[11][2];
    ele[10][3] != ele[11][3];
    ele[10][3] != ele[12][3];
    ele[10][3] != ele[13][3];
    ele[10][3] != ele[14][3];
    ele[10][3] != ele[15][3];
    ele[10][4] != ele[10][10];
    ele[10][4] != ele[10][11];
    ele[10][4] != ele[10][12];
    ele[10][4] != ele[10][13];
    ele[10][4] != ele[10][14];
    ele[10][4] != ele[10][15];
    ele[10][4] != ele[10][5];
    ele[10][4] != ele[10][6];
    ele[10][4] != ele[10][7];
    ele[10][4] != ele[10][8];
    ele[10][4] != ele[10][9];
    ele[10][4] != ele[11][4];
    ele[10][4] != ele[11][5];
    ele[10][4] != ele[11][6];
    ele[10][4] != ele[11][7];
    ele[10][4] != ele[12][4];
    ele[10][4] != ele[13][4];
    ele[10][4] != ele[14][4];
    ele[10][4] != ele[15][4];
    ele[10][5] != ele[10][10];
    ele[10][5] != ele[10][11];
    ele[10][5] != ele[10][12];
    ele[10][5] != ele[10][13];
    ele[10][5] != ele[10][14];
    ele[10][5] != ele[10][15];
    ele[10][5] != ele[10][6];
    ele[10][5] != ele[10][7];
    ele[10][5] != ele[10][8];
    ele[10][5] != ele[10][9];
    ele[10][5] != ele[11][4];
    ele[10][5] != ele[11][5];
    ele[10][5] != ele[11][6];
    ele[10][5] != ele[11][7];
    ele[10][5] != ele[12][5];
    ele[10][5] != ele[13][5];
    ele[10][5] != ele[14][5];
    ele[10][5] != ele[15][5];
    ele[10][6] != ele[10][10];
    ele[10][6] != ele[10][11];
    ele[10][6] != ele[10][12];
    ele[10][6] != ele[10][13];
    ele[10][6] != ele[10][14];
    ele[10][6] != ele[10][15];
    ele[10][6] != ele[10][7];
    ele[10][6] != ele[10][8];
    ele[10][6] != ele[10][9];
    ele[10][6] != ele[11][4];
    ele[10][6] != ele[11][5];
    ele[10][6] != ele[11][6];
    ele[10][6] != ele[11][7];
    ele[10][6] != ele[12][6];
    ele[10][6] != ele[13][6];
    ele[10][6] != ele[14][6];
    ele[10][6] != ele[15][6];
    ele[10][7] != ele[10][10];
    ele[10][7] != ele[10][11];
    ele[10][7] != ele[10][12];
    ele[10][7] != ele[10][13];
    ele[10][7] != ele[10][14];
    ele[10][7] != ele[10][15];
    ele[10][7] != ele[10][8];
    ele[10][7] != ele[10][9];
    ele[10][7] != ele[11][4];
    ele[10][7] != ele[11][5];
    ele[10][7] != ele[11][6];
    ele[10][7] != ele[11][7];
    ele[10][7] != ele[12][7];
    ele[10][7] != ele[13][7];
    ele[10][7] != ele[14][7];
    ele[10][7] != ele[15][7];
    ele[10][8] != ele[10][10];
    ele[10][8] != ele[10][11];
    ele[10][8] != ele[10][12];
    ele[10][8] != ele[10][13];
    ele[10][8] != ele[10][14];
    ele[10][8] != ele[10][15];
    ele[10][8] != ele[10][9];
    ele[10][8] != ele[11][10];
    ele[10][8] != ele[11][11];
    ele[10][8] != ele[11][8];
    ele[10][8] != ele[11][9];
    ele[10][8] != ele[12][8];
    ele[10][8] != ele[13][8];
    ele[10][8] != ele[14][8];
    ele[10][8] != ele[15][8];
    ele[10][9] != ele[10][10];
    ele[10][9] != ele[10][11];
    ele[10][9] != ele[10][12];
    ele[10][9] != ele[10][13];
    ele[10][9] != ele[10][14];
    ele[10][9] != ele[10][15];
    ele[10][9] != ele[11][10];
    ele[10][9] != ele[11][11];
    ele[10][9] != ele[11][8];
    ele[10][9] != ele[11][9];
    ele[10][9] != ele[12][9];
    ele[10][9] != ele[13][9];
    ele[10][9] != ele[14][9];
    ele[10][9] != ele[15][9];
    ele[11][0] != ele[11][1];
    ele[11][0] != ele[11][10];
    ele[11][0] != ele[11][11];
    ele[11][0] != ele[11][12];
    ele[11][0] != ele[11][13];
    ele[11][0] != ele[11][14];
    ele[11][0] != ele[11][15];
    ele[11][0] != ele[11][2];
    ele[11][0] != ele[11][3];
    ele[11][0] != ele[11][4];
    ele[11][0] != ele[11][5];
    ele[11][0] != ele[11][6];
    ele[11][0] != ele[11][7];
    ele[11][0] != ele[11][8];
    ele[11][0] != ele[11][9];
    ele[11][0] != ele[12][0];
    ele[11][0] != ele[13][0];
    ele[11][0] != ele[14][0];
    ele[11][0] != ele[15][0];
    ele[11][1] != ele[11][10];
    ele[11][1] != ele[11][11];
    ele[11][1] != ele[11][12];
    ele[11][1] != ele[11][13];
    ele[11][1] != ele[11][14];
    ele[11][1] != ele[11][15];
    ele[11][1] != ele[11][2];
    ele[11][1] != ele[11][3];
    ele[11][1] != ele[11][4];
    ele[11][1] != ele[11][5];
    ele[11][1] != ele[11][6];
    ele[11][1] != ele[11][7];
    ele[11][1] != ele[11][8];
    ele[11][1] != ele[11][9];
    ele[11][1] != ele[12][1];
    ele[11][1] != ele[13][1];
    ele[11][1] != ele[14][1];
    ele[11][1] != ele[15][1];
    ele[11][10] != ele[11][11];
    ele[11][10] != ele[11][12];
    ele[11][10] != ele[11][13];
    ele[11][10] != ele[11][14];
    ele[11][10] != ele[11][15];
    ele[11][10] != ele[12][10];
    ele[11][10] != ele[13][10];
    ele[11][10] != ele[14][10];
    ele[11][10] != ele[15][10];
    ele[11][11] != ele[11][12];
    ele[11][11] != ele[11][13];
    ele[11][11] != ele[11][14];
    ele[11][11] != ele[11][15];
    ele[11][11] != ele[12][11];
    ele[11][11] != ele[13][11];
    ele[11][11] != ele[14][11];
    ele[11][11] != ele[15][11];
    ele[11][12] != ele[11][13];
    ele[11][12] != ele[11][14];
    ele[11][12] != ele[11][15];
    ele[11][12] != ele[12][12];
    ele[11][12] != ele[13][12];
    ele[11][12] != ele[14][12];
    ele[11][12] != ele[15][12];
    ele[11][13] != ele[11][14];
    ele[11][13] != ele[11][15];
    ele[11][13] != ele[12][13];
    ele[11][13] != ele[13][13];
    ele[11][13] != ele[14][13];
    ele[11][13] != ele[15][13];
    ele[11][14] != ele[11][15];
    ele[11][14] != ele[12][14];
    ele[11][14] != ele[13][14];
    ele[11][14] != ele[14][14];
    ele[11][14] != ele[15][14];
    ele[11][15] != ele[12][15];
    ele[11][15] != ele[13][15];
    ele[11][15] != ele[14][15];
    ele[11][15] != ele[15][15];
    ele[11][2] != ele[11][10];
    ele[11][2] != ele[11][11];
    ele[11][2] != ele[11][12];
    ele[11][2] != ele[11][13];
    ele[11][2] != ele[11][14];
    ele[11][2] != ele[11][15];
    ele[11][2] != ele[11][3];
    ele[11][2] != ele[11][4];
    ele[11][2] != ele[11][5];
    ele[11][2] != ele[11][6];
    ele[11][2] != ele[11][7];
    ele[11][2] != ele[11][8];
    ele[11][2] != ele[11][9];
    ele[11][2] != ele[12][2];
    ele[11][2] != ele[13][2];
    ele[11][2] != ele[14][2];
    ele[11][2] != ele[15][2];
    ele[11][3] != ele[11][10];
    ele[11][3] != ele[11][11];
    ele[11][3] != ele[11][12];
    ele[11][3] != ele[11][13];
    ele[11][3] != ele[11][14];
    ele[11][3] != ele[11][15];
    ele[11][3] != ele[11][4];
    ele[11][3] != ele[11][5];
    ele[11][3] != ele[11][6];
    ele[11][3] != ele[11][7];
    ele[11][3] != ele[11][8];
    ele[11][3] != ele[11][9];
    ele[11][3] != ele[12][3];
    ele[11][3] != ele[13][3];
    ele[11][3] != ele[14][3];
    ele[11][3] != ele[15][3];
    ele[11][4] != ele[11][10];
    ele[11][4] != ele[11][11];
    ele[11][4] != ele[11][12];
    ele[11][4] != ele[11][13];
    ele[11][4] != ele[11][14];
    ele[11][4] != ele[11][15];
    ele[11][4] != ele[11][5];
    ele[11][4] != ele[11][6];
    ele[11][4] != ele[11][7];
    ele[11][4] != ele[11][8];
    ele[11][4] != ele[11][9];
    ele[11][4] != ele[12][4];
    ele[11][4] != ele[13][4];
    ele[11][4] != ele[14][4];
    ele[11][4] != ele[15][4];
    ele[11][5] != ele[11][10];
    ele[11][5] != ele[11][11];
    ele[11][5] != ele[11][12];
    ele[11][5] != ele[11][13];
    ele[11][5] != ele[11][14];
    ele[11][5] != ele[11][15];
    ele[11][5] != ele[11][6];
    ele[11][5] != ele[11][7];
    ele[11][5] != ele[11][8];
    ele[11][5] != ele[11][9];
    ele[11][5] != ele[12][5];
    ele[11][5] != ele[13][5];
    ele[11][5] != ele[14][5];
    ele[11][5] != ele[15][5];
    ele[11][6] != ele[11][10];
    ele[11][6] != ele[11][11];
    ele[11][6] != ele[11][12];
    ele[11][6] != ele[11][13];
    ele[11][6] != ele[11][14];
    ele[11][6] != ele[11][15];
    ele[11][6] != ele[11][7];
    ele[11][6] != ele[11][8];
    ele[11][6] != ele[11][9];
    ele[11][6] != ele[12][6];
    ele[11][6] != ele[13][6];
    ele[11][6] != ele[14][6];
    ele[11][6] != ele[15][6];
    ele[11][7] != ele[11][10];
    ele[11][7] != ele[11][11];
    ele[11][7] != ele[11][12];
    ele[11][7] != ele[11][13];
    ele[11][7] != ele[11][14];
    ele[11][7] != ele[11][15];
    ele[11][7] != ele[11][8];
    ele[11][7] != ele[11][9];
    ele[11][7] != ele[12][7];
    ele[11][7] != ele[13][7];
    ele[11][7] != ele[14][7];
    ele[11][7] != ele[15][7];
    ele[11][8] != ele[11][10];
    ele[11][8] != ele[11][11];
    ele[11][8] != ele[11][12];
    ele[11][8] != ele[11][13];
    ele[11][8] != ele[11][14];
    ele[11][8] != ele[11][15];
    ele[11][8] != ele[11][9];
    ele[11][8] != ele[12][8];
    ele[11][8] != ele[13][8];
    ele[11][8] != ele[14][8];
    ele[11][8] != ele[15][8];
    ele[11][9] != ele[11][10];
    ele[11][9] != ele[11][11];
    ele[11][9] != ele[11][12];
    ele[11][9] != ele[11][13];
    ele[11][9] != ele[11][14];
    ele[11][9] != ele[11][15];
    ele[11][9] != ele[12][9];
    ele[11][9] != ele[13][9];
    ele[11][9] != ele[14][9];
    ele[11][9] != ele[15][9];
    ele[12][0] != ele[12][1];
    ele[12][0] != ele[12][10];
    ele[12][0] != ele[12][11];
    ele[12][0] != ele[12][12];
    ele[12][0] != ele[12][13];
    ele[12][0] != ele[12][14];
    ele[12][0] != ele[12][15];
    ele[12][0] != ele[12][2];
    ele[12][0] != ele[12][3];
    ele[12][0] != ele[12][4];
    ele[12][0] != ele[12][5];
    ele[12][0] != ele[12][6];
    ele[12][0] != ele[12][7];
    ele[12][0] != ele[12][8];
    ele[12][0] != ele[12][9];
    ele[12][0] != ele[13][0];
    ele[12][0] != ele[13][1];
    ele[12][0] != ele[13][2];
    ele[12][0] != ele[13][3];
    ele[12][0] != ele[14][0];
    ele[12][0] != ele[14][1];
    ele[12][0] != ele[14][2];
    ele[12][0] != ele[14][3];
    ele[12][0] != ele[15][0];
    ele[12][0] != ele[15][1];
    ele[12][0] != ele[15][2];
    ele[12][0] != ele[15][3];
    ele[12][1] != ele[12][10];
    ele[12][1] != ele[12][11];
    ele[12][1] != ele[12][12];
    ele[12][1] != ele[12][13];
    ele[12][1] != ele[12][14];
    ele[12][1] != ele[12][15];
    ele[12][1] != ele[12][2];
    ele[12][1] != ele[12][3];
    ele[12][1] != ele[12][4];
    ele[12][1] != ele[12][5];
    ele[12][1] != ele[12][6];
    ele[12][1] != ele[12][7];
    ele[12][1] != ele[12][8];
    ele[12][1] != ele[12][9];
    ele[12][1] != ele[13][0];
    ele[12][1] != ele[13][1];
    ele[12][1] != ele[13][2];
    ele[12][1] != ele[13][3];
    ele[12][1] != ele[14][0];
    ele[12][1] != ele[14][1];
    ele[12][1] != ele[14][2];
    ele[12][1] != ele[14][3];
    ele[12][1] != ele[15][0];
    ele[12][1] != ele[15][1];
    ele[12][1] != ele[15][2];
    ele[12][1] != ele[15][3];
    ele[12][10] != ele[12][11];
    ele[12][10] != ele[12][12];
    ele[12][10] != ele[12][13];
    ele[12][10] != ele[12][14];
    ele[12][10] != ele[12][15];
    ele[12][10] != ele[13][10];
    ele[12][10] != ele[13][11];
    ele[12][10] != ele[13][8];
    ele[12][10] != ele[13][9];
    ele[12][10] != ele[14][10];
    ele[12][10] != ele[14][11];
    ele[12][10] != ele[14][8];
    ele[12][10] != ele[14][9];
    ele[12][10] != ele[15][10];
    ele[12][10] != ele[15][11];
    ele[12][10] != ele[15][8];
    ele[12][10] != ele[15][9];
    ele[12][11] != ele[12][12];
    ele[12][11] != ele[12][13];
    ele[12][11] != ele[12][14];
    ele[12][11] != ele[12][15];
    ele[12][11] != ele[13][10];
    ele[12][11] != ele[13][11];
    ele[12][11] != ele[13][8];
    ele[12][11] != ele[13][9];
    ele[12][11] != ele[14][10];
    ele[12][11] != ele[14][11];
    ele[12][11] != ele[14][8];
    ele[12][11] != ele[14][9];
    ele[12][11] != ele[15][10];
    ele[12][11] != ele[15][11];
    ele[12][11] != ele[15][8];
    ele[12][11] != ele[15][9];
    ele[12][12] != ele[12][13];
    ele[12][12] != ele[12][14];
    ele[12][12] != ele[12][15];
    ele[12][12] != ele[13][12];
    ele[12][12] != ele[13][13];
    ele[12][12] != ele[13][14];
    ele[12][12] != ele[13][15];
    ele[12][12] != ele[14][12];
    ele[12][12] != ele[14][13];
    ele[12][12] != ele[14][14];
    ele[12][12] != ele[14][15];
    ele[12][12] != ele[15][12];
    ele[12][12] != ele[15][13];
    ele[12][12] != ele[15][14];
    ele[12][12] != ele[15][15];
    ele[12][13] != ele[12][14];
    ele[12][13] != ele[12][15];
    ele[12][13] != ele[13][12];
    ele[12][13] != ele[13][13];
    ele[12][13] != ele[13][14];
    ele[12][13] != ele[13][15];
    ele[12][13] != ele[14][12];
    ele[12][13] != ele[14][13];
    ele[12][13] != ele[14][14];
    ele[12][13] != ele[14][15];
    ele[12][13] != ele[15][12];
    ele[12][13] != ele[15][13];
    ele[12][13] != ele[15][14];
    ele[12][13] != ele[15][15];
    ele[12][14] != ele[12][15];
    ele[12][14] != ele[13][12];
    ele[12][14] != ele[13][13];
    ele[12][14] != ele[13][14];
    ele[12][14] != ele[13][15];
    ele[12][14] != ele[14][12];
    ele[12][14] != ele[14][13];
    ele[12][14] != ele[14][14];
    ele[12][14] != ele[14][15];
    ele[12][14] != ele[15][12];
    ele[12][14] != ele[15][13];
    ele[12][14] != ele[15][14];
    ele[12][14] != ele[15][15];
    ele[12][15] != ele[13][12];
    ele[12][15] != ele[13][13];
    ele[12][15] != ele[13][14];
    ele[12][15] != ele[13][15];
    ele[12][15] != ele[14][12];
    ele[12][15] != ele[14][13];
    ele[12][15] != ele[14][14];
    ele[12][15] != ele[14][15];
    ele[12][15] != ele[15][12];
    ele[12][15] != ele[15][13];
    ele[12][15] != ele[15][14];
    ele[12][15] != ele[15][15];
    ele[12][2] != ele[12][10];
    ele[12][2] != ele[12][11];
    ele[12][2] != ele[12][12];
    ele[12][2] != ele[12][13];
    ele[12][2] != ele[12][14];
    ele[12][2] != ele[12][15];
    ele[12][2] != ele[12][3];
    ele[12][2] != ele[12][4];
    ele[12][2] != ele[12][5];
    ele[12][2] != ele[12][6];
    ele[12][2] != ele[12][7];
    ele[12][2] != ele[12][8];
    ele[12][2] != ele[12][9];
    ele[12][2] != ele[13][0];
    ele[12][2] != ele[13][1];
    ele[12][2] != ele[13][2];
    ele[12][2] != ele[13][3];
    ele[12][2] != ele[14][0];
    ele[12][2] != ele[14][1];
    ele[12][2] != ele[14][2];
    ele[12][2] != ele[14][3];
    ele[12][2] != ele[15][0];
    ele[12][2] != ele[15][1];
    ele[12][2] != ele[15][2];
    ele[12][2] != ele[15][3];
    ele[12][3] != ele[12][10];
    ele[12][3] != ele[12][11];
    ele[12][3] != ele[12][12];
    ele[12][3] != ele[12][13];
    ele[12][3] != ele[12][14];
    ele[12][3] != ele[12][15];
    ele[12][3] != ele[12][4];
    ele[12][3] != ele[12][5];
    ele[12][3] != ele[12][6];
    ele[12][3] != ele[12][7];
    ele[12][3] != ele[12][8];
    ele[12][3] != ele[12][9];
    ele[12][3] != ele[13][0];
    ele[12][3] != ele[13][1];
    ele[12][3] != ele[13][2];
    ele[12][3] != ele[13][3];
    ele[12][3] != ele[14][0];
    ele[12][3] != ele[14][1];
    ele[12][3] != ele[14][2];
    ele[12][3] != ele[14][3];
    ele[12][3] != ele[15][0];
    ele[12][3] != ele[15][1];
    ele[12][3] != ele[15][2];
    ele[12][3] != ele[15][3];
    ele[12][4] != ele[12][10];
    ele[12][4] != ele[12][11];
    ele[12][4] != ele[12][12];
    ele[12][4] != ele[12][13];
    ele[12][4] != ele[12][14];
    ele[12][4] != ele[12][15];
    ele[12][4] != ele[12][5];
    ele[12][4] != ele[12][6];
    ele[12][4] != ele[12][7];
    ele[12][4] != ele[12][8];
    ele[12][4] != ele[12][9];
    ele[12][4] != ele[13][4];
    ele[12][4] != ele[13][5];
    ele[12][4] != ele[13][6];
    ele[12][4] != ele[13][7];
    ele[12][4] != ele[14][4];
    ele[12][4] != ele[14][5];
    ele[12][4] != ele[14][6];
    ele[12][4] != ele[14][7];
    ele[12][4] != ele[15][4];
    ele[12][4] != ele[15][5];
    ele[12][4] != ele[15][6];
    ele[12][4] != ele[15][7];
    ele[12][5] != ele[12][10];
    ele[12][5] != ele[12][11];
    ele[12][5] != ele[12][12];
    ele[12][5] != ele[12][13];
    ele[12][5] != ele[12][14];
    ele[12][5] != ele[12][15];
    ele[12][5] != ele[12][6];
    ele[12][5] != ele[12][7];
    ele[12][5] != ele[12][8];
    ele[12][5] != ele[12][9];
    ele[12][5] != ele[13][4];
    ele[12][5] != ele[13][5];
    ele[12][5] != ele[13][6];
    ele[12][5] != ele[13][7];
    ele[12][5] != ele[14][4];
    ele[12][5] != ele[14][5];
    ele[12][5] != ele[14][6];
    ele[12][5] != ele[14][7];
    ele[12][5] != ele[15][4];
    ele[12][5] != ele[15][5];
    ele[12][5] != ele[15][6];
    ele[12][5] != ele[15][7];
    ele[12][6] != ele[12][10];
    ele[12][6] != ele[12][11];
    ele[12][6] != ele[12][12];
    ele[12][6] != ele[12][13];
    ele[12][6] != ele[12][14];
    ele[12][6] != ele[12][15];
    ele[12][6] != ele[12][7];
    ele[12][6] != ele[12][8];
    ele[12][6] != ele[12][9];
    ele[12][6] != ele[13][4];
    ele[12][6] != ele[13][5];
    ele[12][6] != ele[13][6];
    ele[12][6] != ele[13][7];
    ele[12][6] != ele[14][4];
    ele[12][6] != ele[14][5];
    ele[12][6] != ele[14][6];
    ele[12][6] != ele[14][7];
    ele[12][6] != ele[15][4];
    ele[12][6] != ele[15][5];
    ele[12][6] != ele[15][6];
    ele[12][6] != ele[15][7];
    ele[12][7] != ele[12][10];
    ele[12][7] != ele[12][11];
    ele[12][7] != ele[12][12];
    ele[12][7] != ele[12][13];
    ele[12][7] != ele[12][14];
    ele[12][7] != ele[12][15];
    ele[12][7] != ele[12][8];
    ele[12][7] != ele[12][9];
    ele[12][7] != ele[13][4];
    ele[12][7] != ele[13][5];
    ele[12][7] != ele[13][6];
    ele[12][7] != ele[13][7];
    ele[12][7] != ele[14][4];
    ele[12][7] != ele[14][5];
    ele[12][7] != ele[14][6];
    ele[12][7] != ele[14][7];
    ele[12][7] != ele[15][4];
    ele[12][7] != ele[15][5];
    ele[12][7] != ele[15][6];
    ele[12][7] != ele[15][7];
    ele[12][8] != ele[12][10];
    ele[12][8] != ele[12][11];
    ele[12][8] != ele[12][12];
    ele[12][8] != ele[12][13];
    ele[12][8] != ele[12][14];
    ele[12][8] != ele[12][15];
    ele[12][8] != ele[12][9];
    ele[12][8] != ele[13][10];
    ele[12][8] != ele[13][11];
    ele[12][8] != ele[13][8];
    ele[12][8] != ele[13][9];
    ele[12][8] != ele[14][10];
    ele[12][8] != ele[14][11];
    ele[12][8] != ele[14][8];
    ele[12][8] != ele[14][9];
    ele[12][8] != ele[15][10];
    ele[12][8] != ele[15][11];
    ele[12][8] != ele[15][8];
    ele[12][8] != ele[15][9];
    ele[12][9] != ele[12][10];
    ele[12][9] != ele[12][11];
    ele[12][9] != ele[12][12];
    ele[12][9] != ele[12][13];
    ele[12][9] != ele[12][14];
    ele[12][9] != ele[12][15];
    ele[12][9] != ele[13][10];
    ele[12][9] != ele[13][11];
    ele[12][9] != ele[13][8];
    ele[12][9] != ele[13][9];
    ele[12][9] != ele[14][10];
    ele[12][9] != ele[14][11];
    ele[12][9] != ele[14][8];
    ele[12][9] != ele[14][9];
    ele[12][9] != ele[15][10];
    ele[12][9] != ele[15][11];
    ele[12][9] != ele[15][8];
    ele[12][9] != ele[15][9];
    ele[13][0] != ele[13][1];
    ele[13][0] != ele[13][10];
    ele[13][0] != ele[13][11];
    ele[13][0] != ele[13][12];
    ele[13][0] != ele[13][13];
    ele[13][0] != ele[13][14];
    ele[13][0] != ele[13][15];
    ele[13][0] != ele[13][2];
    ele[13][0] != ele[13][3];
    ele[13][0] != ele[13][4];
    ele[13][0] != ele[13][5];
    ele[13][0] != ele[13][6];
    ele[13][0] != ele[13][7];
    ele[13][0] != ele[13][8];
    ele[13][0] != ele[13][9];
    ele[13][0] != ele[14][0];
    ele[13][0] != ele[14][1];
    ele[13][0] != ele[14][2];
    ele[13][0] != ele[14][3];
    ele[13][0] != ele[15][0];
    ele[13][0] != ele[15][1];
    ele[13][0] != ele[15][2];
    ele[13][0] != ele[15][3];
    ele[13][1] != ele[13][10];
    ele[13][1] != ele[13][11];
    ele[13][1] != ele[13][12];
    ele[13][1] != ele[13][13];
    ele[13][1] != ele[13][14];
    ele[13][1] != ele[13][15];
    ele[13][1] != ele[13][2];
    ele[13][1] != ele[13][3];
    ele[13][1] != ele[13][4];
    ele[13][1] != ele[13][5];
    ele[13][1] != ele[13][6];
    ele[13][1] != ele[13][7];
    ele[13][1] != ele[13][8];
    ele[13][1] != ele[13][9];
    ele[13][1] != ele[14][0];
    ele[13][1] != ele[14][1];
    ele[13][1] != ele[14][2];
    ele[13][1] != ele[14][3];
    ele[13][1] != ele[15][0];
    ele[13][1] != ele[15][1];
    ele[13][1] != ele[15][2];
    ele[13][1] != ele[15][3];
    ele[13][10] != ele[13][11];
    ele[13][10] != ele[13][12];
    ele[13][10] != ele[13][13];
    ele[13][10] != ele[13][14];
    ele[13][10] != ele[13][15];
    ele[13][10] != ele[14][10];
    ele[13][10] != ele[14][11];
    ele[13][10] != ele[14][8];
    ele[13][10] != ele[14][9];
    ele[13][10] != ele[15][10];
    ele[13][10] != ele[15][11];
    ele[13][10] != ele[15][8];
    ele[13][10] != ele[15][9];
    ele[13][11] != ele[13][12];
    ele[13][11] != ele[13][13];
    ele[13][11] != ele[13][14];
    ele[13][11] != ele[13][15];
    ele[13][11] != ele[14][10];
    ele[13][11] != ele[14][11];
    ele[13][11] != ele[14][8];
    ele[13][11] != ele[14][9];
    ele[13][11] != ele[15][10];
    ele[13][11] != ele[15][11];
    ele[13][11] != ele[15][8];
    ele[13][11] != ele[15][9];
    ele[13][12] != ele[13][13];
    ele[13][12] != ele[13][14];
    ele[13][12] != ele[13][15];
    ele[13][12] != ele[14][12];
    ele[13][12] != ele[14][13];
    ele[13][12] != ele[14][14];
    ele[13][12] != ele[14][15];
    ele[13][12] != ele[15][12];
    ele[13][12] != ele[15][13];
    ele[13][12] != ele[15][14];
    ele[13][12] != ele[15][15];
    ele[13][13] != ele[13][14];
    ele[13][13] != ele[13][15];
    ele[13][13] != ele[14][12];
    ele[13][13] != ele[14][13];
    ele[13][13] != ele[14][14];
    ele[13][13] != ele[14][15];
    ele[13][13] != ele[15][12];
    ele[13][13] != ele[15][13];
    ele[13][13] != ele[15][14];
    ele[13][13] != ele[15][15];
    ele[13][14] != ele[13][15];
    ele[13][14] != ele[14][12];
    ele[13][14] != ele[14][13];
    ele[13][14] != ele[14][14];
    ele[13][14] != ele[14][15];
    ele[13][14] != ele[15][12];
    ele[13][14] != ele[15][13];
    ele[13][14] != ele[15][14];
    ele[13][14] != ele[15][15];
    ele[13][15] != ele[14][12];
    ele[13][15] != ele[14][13];
    ele[13][15] != ele[14][14];
    ele[13][15] != ele[14][15];
    ele[13][15] != ele[15][12];
    ele[13][15] != ele[15][13];
    ele[13][15] != ele[15][14];
    ele[13][15] != ele[15][15];
    ele[13][2] != ele[13][10];
    ele[13][2] != ele[13][11];
    ele[13][2] != ele[13][12];
    ele[13][2] != ele[13][13];
    ele[13][2] != ele[13][14];
    ele[13][2] != ele[13][15];
    ele[13][2] != ele[13][3];
    ele[13][2] != ele[13][4];
    ele[13][2] != ele[13][5];
    ele[13][2] != ele[13][6];
    ele[13][2] != ele[13][7];
    ele[13][2] != ele[13][8];
    ele[13][2] != ele[13][9];
    ele[13][2] != ele[14][0];
    ele[13][2] != ele[14][1];
    ele[13][2] != ele[14][2];
    ele[13][2] != ele[14][3];
    ele[13][2] != ele[15][0];
    ele[13][2] != ele[15][1];
    ele[13][2] != ele[15][2];
    ele[13][2] != ele[15][3];
    ele[13][3] != ele[13][10];
    ele[13][3] != ele[13][11];
    ele[13][3] != ele[13][12];
    ele[13][3] != ele[13][13];
    ele[13][3] != ele[13][14];
    ele[13][3] != ele[13][15];
    ele[13][3] != ele[13][4];
    ele[13][3] != ele[13][5];
    ele[13][3] != ele[13][6];
    ele[13][3] != ele[13][7];
    ele[13][3] != ele[13][8];
    ele[13][3] != ele[13][9];
    ele[13][3] != ele[14][0];
    ele[13][3] != ele[14][1];
    ele[13][3] != ele[14][2];
    ele[13][3] != ele[14][3];
    ele[13][3] != ele[15][0];
    ele[13][3] != ele[15][1];
    ele[13][3] != ele[15][2];
    ele[13][3] != ele[15][3];
    ele[13][4] != ele[13][10];
    ele[13][4] != ele[13][11];
    ele[13][4] != ele[13][12];
    ele[13][4] != ele[13][13];
    ele[13][4] != ele[13][14];
    ele[13][4] != ele[13][15];
    ele[13][4] != ele[13][5];
    ele[13][4] != ele[13][6];
    ele[13][4] != ele[13][7];
    ele[13][4] != ele[13][8];
    ele[13][4] != ele[13][9];
    ele[13][4] != ele[14][4];
    ele[13][4] != ele[14][5];
    ele[13][4] != ele[14][6];
    ele[13][4] != ele[14][7];
    ele[13][4] != ele[15][4];
    ele[13][4] != ele[15][5];
    ele[13][4] != ele[15][6];
    ele[13][4] != ele[15][7];
    ele[13][5] != ele[13][10];
    ele[13][5] != ele[13][11];
    ele[13][5] != ele[13][12];
    ele[13][5] != ele[13][13];
    ele[13][5] != ele[13][14];
    ele[13][5] != ele[13][15];
    ele[13][5] != ele[13][6];
    ele[13][5] != ele[13][7];
    ele[13][5] != ele[13][8];
    ele[13][5] != ele[13][9];
    ele[13][5] != ele[14][4];
    ele[13][5] != ele[14][5];
    ele[13][5] != ele[14][6];
    ele[13][5] != ele[14][7];
    ele[13][5] != ele[15][4];
    ele[13][5] != ele[15][5];
    ele[13][5] != ele[15][6];
    ele[13][5] != ele[15][7];
    ele[13][6] != ele[13][10];
    ele[13][6] != ele[13][11];
    ele[13][6] != ele[13][12];
    ele[13][6] != ele[13][13];
    ele[13][6] != ele[13][14];
    ele[13][6] != ele[13][15];
    ele[13][6] != ele[13][7];
    ele[13][6] != ele[13][8];
    ele[13][6] != ele[13][9];
    ele[13][6] != ele[14][4];
    ele[13][6] != ele[14][5];
    ele[13][6] != ele[14][6];
    ele[13][6] != ele[14][7];
    ele[13][6] != ele[15][4];
    ele[13][6] != ele[15][5];
    ele[13][6] != ele[15][6];
    ele[13][6] != ele[15][7];
    ele[13][7] != ele[13][10];
    ele[13][7] != ele[13][11];
    ele[13][7] != ele[13][12];
    ele[13][7] != ele[13][13];
    ele[13][7] != ele[13][14];
    ele[13][7] != ele[13][15];
    ele[13][7] != ele[13][8];
    ele[13][7] != ele[13][9];
    ele[13][7] != ele[14][4];
    ele[13][7] != ele[14][5];
    ele[13][7] != ele[14][6];
    ele[13][7] != ele[14][7];
    ele[13][7] != ele[15][4];
    ele[13][7] != ele[15][5];
    ele[13][7] != ele[15][6];
    ele[13][7] != ele[15][7];
    ele[13][8] != ele[13][10];
    ele[13][8] != ele[13][11];
    ele[13][8] != ele[13][12];
    ele[13][8] != ele[13][13];
    ele[13][8] != ele[13][14];
    ele[13][8] != ele[13][15];
    ele[13][8] != ele[13][9];
    ele[13][8] != ele[14][10];
    ele[13][8] != ele[14][11];
    ele[13][8] != ele[14][8];
    ele[13][8] != ele[14][9];
    ele[13][8] != ele[15][10];
    ele[13][8] != ele[15][11];
    ele[13][8] != ele[15][8];
    ele[13][8] != ele[15][9];
    ele[13][9] != ele[13][10];
    ele[13][9] != ele[13][11];
    ele[13][9] != ele[13][12];
    ele[13][9] != ele[13][13];
    ele[13][9] != ele[13][14];
    ele[13][9] != ele[13][15];
    ele[13][9] != ele[14][10];
    ele[13][9] != ele[14][11];
    ele[13][9] != ele[14][8];
    ele[13][9] != ele[14][9];
    ele[13][9] != ele[15][10];
    ele[13][9] != ele[15][11];
    ele[13][9] != ele[15][8];
    ele[13][9] != ele[15][9];
    ele[14][0] != ele[14][1];
    ele[14][0] != ele[14][10];
    ele[14][0] != ele[14][11];
    ele[14][0] != ele[14][12];
    ele[14][0] != ele[14][13];
    ele[14][0] != ele[14][14];
    ele[14][0] != ele[14][15];
    ele[14][0] != ele[14][2];
    ele[14][0] != ele[14][3];
    ele[14][0] != ele[14][4];
    ele[14][0] != ele[14][5];
    ele[14][0] != ele[14][6];
    ele[14][0] != ele[14][7];
    ele[14][0] != ele[14][8];
    ele[14][0] != ele[14][9];
    ele[14][0] != ele[15][0];
    ele[14][0] != ele[15][1];
    ele[14][0] != ele[15][2];
    ele[14][0] != ele[15][3];
    ele[14][1] != ele[14][10];
    ele[14][1] != ele[14][11];
    ele[14][1] != ele[14][12];
    ele[14][1] != ele[14][13];
    ele[14][1] != ele[14][14];
    ele[14][1] != ele[14][15];
    ele[14][1] != ele[14][2];
    ele[14][1] != ele[14][3];
    ele[14][1] != ele[14][4];
    ele[14][1] != ele[14][5];
    ele[14][1] != ele[14][6];
    ele[14][1] != ele[14][7];
    ele[14][1] != ele[14][8];
    ele[14][1] != ele[14][9];
    ele[14][1] != ele[15][0];
    ele[14][1] != ele[15][1];
    ele[14][1] != ele[15][2];
    ele[14][1] != ele[15][3];
    ele[14][10] != ele[14][11];
    ele[14][10] != ele[14][12];
    ele[14][10] != ele[14][13];
    ele[14][10] != ele[14][14];
    ele[14][10] != ele[14][15];
    ele[14][10] != ele[15][10];
    ele[14][10] != ele[15][11];
    ele[14][10] != ele[15][8];
    ele[14][10] != ele[15][9];
    ele[14][11] != ele[14][12];
    ele[14][11] != ele[14][13];
    ele[14][11] != ele[14][14];
    ele[14][11] != ele[14][15];
    ele[14][11] != ele[15][10];
    ele[14][11] != ele[15][11];
    ele[14][11] != ele[15][8];
    ele[14][11] != ele[15][9];
    ele[14][12] != ele[14][13];
    ele[14][12] != ele[14][14];
    ele[14][12] != ele[14][15];
    ele[14][12] != ele[15][12];
    ele[14][12] != ele[15][13];
    ele[14][12] != ele[15][14];
    ele[14][12] != ele[15][15];
    ele[14][13] != ele[14][14];
    ele[14][13] != ele[14][15];
    ele[14][13] != ele[15][12];
    ele[14][13] != ele[15][13];
    ele[14][13] != ele[15][14];
    ele[14][13] != ele[15][15];
    ele[14][14] != ele[14][15];
    ele[14][14] != ele[15][12];
    ele[14][14] != ele[15][13];
    ele[14][14] != ele[15][14];
    ele[14][14] != ele[15][15];
    ele[14][15] != ele[15][12];
    ele[14][15] != ele[15][13];
    ele[14][15] != ele[15][14];
    ele[14][15] != ele[15][15];
    ele[14][2] != ele[14][10];
    ele[14][2] != ele[14][11];
    ele[14][2] != ele[14][12];
    ele[14][2] != ele[14][13];
    ele[14][2] != ele[14][14];
    ele[14][2] != ele[14][15];
    ele[14][2] != ele[14][3];
    ele[14][2] != ele[14][4];
    ele[14][2] != ele[14][5];
    ele[14][2] != ele[14][6];
    ele[14][2] != ele[14][7];
    ele[14][2] != ele[14][8];
    ele[14][2] != ele[14][9];
    ele[14][2] != ele[15][0];
    ele[14][2] != ele[15][1];
    ele[14][2] != ele[15][2];
    ele[14][2] != ele[15][3];
    ele[14][3] != ele[14][10];
    ele[14][3] != ele[14][11];
    ele[14][3] != ele[14][12];
    ele[14][3] != ele[14][13];
    ele[14][3] != ele[14][14];
    ele[14][3] != ele[14][15];
    ele[14][3] != ele[14][4];
    ele[14][3] != ele[14][5];
    ele[14][3] != ele[14][6];
    ele[14][3] != ele[14][7];
    ele[14][3] != ele[14][8];
    ele[14][3] != ele[14][9];
    ele[14][3] != ele[15][0];
    ele[14][3] != ele[15][1];
    ele[14][3] != ele[15][2];
    ele[14][3] != ele[15][3];
    ele[14][4] != ele[14][10];
    ele[14][4] != ele[14][11];
    ele[14][4] != ele[14][12];
    ele[14][4] != ele[14][13];
    ele[14][4] != ele[14][14];
    ele[14][4] != ele[14][15];
    ele[14][4] != ele[14][5];
    ele[14][4] != ele[14][6];
    ele[14][4] != ele[14][7];
    ele[14][4] != ele[14][8];
    ele[14][4] != ele[14][9];
    ele[14][4] != ele[15][4];
    ele[14][4] != ele[15][5];
    ele[14][4] != ele[15][6];
    ele[14][4] != ele[15][7];
    ele[14][5] != ele[14][10];
    ele[14][5] != ele[14][11];
    ele[14][5] != ele[14][12];
    ele[14][5] != ele[14][13];
    ele[14][5] != ele[14][14];
    ele[14][5] != ele[14][15];
    ele[14][5] != ele[14][6];
    ele[14][5] != ele[14][7];
    ele[14][5] != ele[14][8];
    ele[14][5] != ele[14][9];
    ele[14][5] != ele[15][4];
    ele[14][5] != ele[15][5];
    ele[14][5] != ele[15][6];
    ele[14][5] != ele[15][7];
    ele[14][6] != ele[14][10];
    ele[14][6] != ele[14][11];
    ele[14][6] != ele[14][12];
    ele[14][6] != ele[14][13];
    ele[14][6] != ele[14][14];
    ele[14][6] != ele[14][15];
    ele[14][6] != ele[14][7];
    ele[14][6] != ele[14][8];
    ele[14][6] != ele[14][9];
    ele[14][6] != ele[15][4];
    ele[14][6] != ele[15][5];
    ele[14][6] != ele[15][6];
    ele[14][6] != ele[15][7];
    ele[14][7] != ele[14][10];
    ele[14][7] != ele[14][11];
    ele[14][7] != ele[14][12];
    ele[14][7] != ele[14][13];
    ele[14][7] != ele[14][14];
    ele[14][7] != ele[14][15];
    ele[14][7] != ele[14][8];
    ele[14][7] != ele[14][9];
    ele[14][7] != ele[15][4];
    ele[14][7] != ele[15][5];
    ele[14][7] != ele[15][6];
    ele[14][7] != ele[15][7];
    ele[14][8] != ele[14][10];
    ele[14][8] != ele[14][11];
    ele[14][8] != ele[14][12];
    ele[14][8] != ele[14][13];
    ele[14][8] != ele[14][14];
    ele[14][8] != ele[14][15];
    ele[14][8] != ele[14][9];
    ele[14][8] != ele[15][10];
    ele[14][8] != ele[15][11];
    ele[14][8] != ele[15][8];
    ele[14][8] != ele[15][9];
    ele[14][9] != ele[14][10];
    ele[14][9] != ele[14][11];
    ele[14][9] != ele[14][12];
    ele[14][9] != ele[14][13];
    ele[14][9] != ele[14][14];
    ele[14][9] != ele[14][15];
    ele[14][9] != ele[15][10];
    ele[14][9] != ele[15][11];
    ele[14][9] != ele[15][8];
    ele[14][9] != ele[15][9];
    ele[15][0] != ele[15][1];
    ele[15][0] != ele[15][10];
    ele[15][0] != ele[15][11];
    ele[15][0] != ele[15][12];
    ele[15][0] != ele[15][13];
    ele[15][0] != ele[15][14];
    ele[15][0] != ele[15][15];
    ele[15][0] != ele[15][2];
    ele[15][0] != ele[15][3];
    ele[15][0] != ele[15][4];
    ele[15][0] != ele[15][5];
    ele[15][0] != ele[15][6];
    ele[15][0] != ele[15][7];
    ele[15][0] != ele[15][8];
    ele[15][0] != ele[15][9];
    ele[15][1] != ele[15][10];
    ele[15][1] != ele[15][11];
    ele[15][1] != ele[15][12];
    ele[15][1] != ele[15][13];
    ele[15][1] != ele[15][14];
    ele[15][1] != ele[15][15];
    ele[15][1] != ele[15][2];
    ele[15][1] != ele[15][3];
    ele[15][1] != ele[15][4];
    ele[15][1] != ele[15][5];
    ele[15][1] != ele[15][6];
    ele[15][1] != ele[15][7];
    ele[15][1] != ele[15][8];
    ele[15][1] != ele[15][9];
    ele[15][10] != ele[15][11];
    ele[15][10] != ele[15][12];
    ele[15][10] != ele[15][13];
    ele[15][10] != ele[15][14];
    ele[15][10] != ele[15][15];
    ele[15][11] != ele[15][12];
    ele[15][11] != ele[15][13];
    ele[15][11] != ele[15][14];
    ele[15][11] != ele[15][15];
    ele[15][12] != ele[15][13];
    ele[15][12] != ele[15][14];
    ele[15][12] != ele[15][15];
    ele[15][13] != ele[15][14];
    ele[15][13] != ele[15][15];
    ele[15][14] != ele[15][15];
    ele[15][2] != ele[15][10];
    ele[15][2] != ele[15][11];
    ele[15][2] != ele[15][12];
    ele[15][2] != ele[15][13];
    ele[15][2] != ele[15][14];
    ele[15][2] != ele[15][15];
    ele[15][2] != ele[15][3];
    ele[15][2] != ele[15][4];
    ele[15][2] != ele[15][5];
    ele[15][2] != ele[15][6];
    ele[15][2] != ele[15][7];
    ele[15][2] != ele[15][8];
    ele[15][2] != ele[15][9];
    ele[15][3] != ele[15][10];
    ele[15][3] != ele[15][11];
    ele[15][3] != ele[15][12];
    ele[15][3] != ele[15][13];
    ele[15][3] != ele[15][14];
    ele[15][3] != ele[15][15];
    ele[15][3] != ele[15][4];
    ele[15][3] != ele[15][5];
    ele[15][3] != ele[15][6];
    ele[15][3] != ele[15][7];
    ele[15][3] != ele[15][8];
    ele[15][3] != ele[15][9];
    ele[15][4] != ele[15][10];
    ele[15][4] != ele[15][11];
    ele[15][4] != ele[15][12];
    ele[15][4] != ele[15][13];
    ele[15][4] != ele[15][14];
    ele[15][4] != ele[15][15];
    ele[15][4] != ele[15][5];
    ele[15][4] != ele[15][6];
    ele[15][4] != ele[15][7];
    ele[15][4] != ele[15][8];
    ele[15][4] != ele[15][9];
    ele[15][5] != ele[15][10];
    ele[15][5] != ele[15][11];
    ele[15][5] != ele[15][12];
    ele[15][5] != ele[15][13];
    ele[15][5] != ele[15][14];
    ele[15][5] != ele[15][15];
    ele[15][5] != ele[15][6];
    ele[15][5] != ele[15][7];
    ele[15][5] != ele[15][8];
    ele[15][5] != ele[15][9];
    ele[15][6] != ele[15][10];
    ele[15][6] != ele[15][11];
    ele[15][6] != ele[15][12];
    ele[15][6] != ele[15][13];
    ele[15][6] != ele[15][14];
    ele[15][6] != ele[15][15];
    ele[15][6] != ele[15][7];
    ele[15][6] != ele[15][8];
    ele[15][6] != ele[15][9];
    ele[15][7] != ele[15][10];
    ele[15][7] != ele[15][11];
    ele[15][7] != ele[15][12];
    ele[15][7] != ele[15][13];
    ele[15][7] != ele[15][14];
    ele[15][7] != ele[15][15];
    ele[15][7] != ele[15][8];
    ele[15][7] != ele[15][9];
    ele[15][8] != ele[15][10];
    ele[15][8] != ele[15][11];
    ele[15][8] != ele[15][12];
    ele[15][8] != ele[15][13];
    ele[15][8] != ele[15][14];
    ele[15][8] != ele[15][15];
    ele[15][8] != ele[15][9];
    ele[15][9] != ele[15][10];
    ele[15][9] != ele[15][11];
    ele[15][9] != ele[15][12];
    ele[15][9] != ele[15][13];
    ele[15][9] != ele[15][14];
    ele[15][9] != ele[15][15];
    ele[2][0] != ele[10][0];
    ele[2][0] != ele[11][0];
    ele[2][0] != ele[12][0];
    ele[2][0] != ele[13][0];
    ele[2][0] != ele[14][0];
    ele[2][0] != ele[15][0];
    ele[2][0] != ele[2][1];
    ele[2][0] != ele[2][10];
    ele[2][0] != ele[2][11];
    ele[2][0] != ele[2][12];
    ele[2][0] != ele[2][13];
    ele[2][0] != ele[2][14];
    ele[2][0] != ele[2][15];
    ele[2][0] != ele[2][2];
    ele[2][0] != ele[2][3];
    ele[2][0] != ele[2][4];
    ele[2][0] != ele[2][5];
    ele[2][0] != ele[2][6];
    ele[2][0] != ele[2][7];
    ele[2][0] != ele[2][8];
    ele[2][0] != ele[2][9];
    ele[2][0] != ele[3][0];
    ele[2][0] != ele[3][1];
    ele[2][0] != ele[3][2];
    ele[2][0] != ele[3][3];
    ele[2][0] != ele[4][0];
    ele[2][0] != ele[5][0];
    ele[2][0] != ele[6][0];
    ele[2][0] != ele[7][0];
    ele[2][0] != ele[8][0];
    ele[2][0] != ele[9][0];
    ele[2][1] != ele[10][1];
    ele[2][1] != ele[11][1];
    ele[2][1] != ele[12][1];
    ele[2][1] != ele[13][1];
    ele[2][1] != ele[14][1];
    ele[2][1] != ele[15][1];
    ele[2][1] != ele[2][10];
    ele[2][1] != ele[2][11];
    ele[2][1] != ele[2][12];
    ele[2][1] != ele[2][13];
    ele[2][1] != ele[2][14];
    ele[2][1] != ele[2][15];
    ele[2][1] != ele[2][2];
    ele[2][1] != ele[2][3];
    ele[2][1] != ele[2][4];
    ele[2][1] != ele[2][5];
    ele[2][1] != ele[2][6];
    ele[2][1] != ele[2][7];
    ele[2][1] != ele[2][8];
    ele[2][1] != ele[2][9];
    ele[2][1] != ele[3][0];
    ele[2][1] != ele[3][1];
    ele[2][1] != ele[3][2];
    ele[2][1] != ele[3][3];
    ele[2][1] != ele[4][1];
    ele[2][1] != ele[5][1];
    ele[2][1] != ele[6][1];
    ele[2][1] != ele[7][1];
    ele[2][1] != ele[8][1];
    ele[2][1] != ele[9][1];
    ele[2][10] != ele[10][10];
    ele[2][10] != ele[11][10];
    ele[2][10] != ele[12][10];
    ele[2][10] != ele[13][10];
    ele[2][10] != ele[14][10];
    ele[2][10] != ele[15][10];
    ele[2][10] != ele[2][11];
    ele[2][10] != ele[2][12];
    ele[2][10] != ele[2][13];
    ele[2][10] != ele[2][14];
    ele[2][10] != ele[2][15];
    ele[2][10] != ele[3][10];
    ele[2][10] != ele[3][11];
    ele[2][10] != ele[3][8];
    ele[2][10] != ele[3][9];
    ele[2][10] != ele[4][10];
    ele[2][10] != ele[5][10];
    ele[2][10] != ele[6][10];
    ele[2][10] != ele[7][10];
    ele[2][10] != ele[8][10];
    ele[2][10] != ele[9][10];
    ele[2][11] != ele[10][11];
    ele[2][11] != ele[11][11];
    ele[2][11] != ele[12][11];
    ele[2][11] != ele[13][11];
    ele[2][11] != ele[14][11];
    ele[2][11] != ele[15][11];
    ele[2][11] != ele[2][12];
    ele[2][11] != ele[2][13];
    ele[2][11] != ele[2][14];
    ele[2][11] != ele[2][15];
    ele[2][11] != ele[3][10];
    ele[2][11] != ele[3][11];
    ele[2][11] != ele[3][8];
    ele[2][11] != ele[3][9];
    ele[2][11] != ele[4][11];
    ele[2][11] != ele[5][11];
    ele[2][11] != ele[6][11];
    ele[2][11] != ele[7][11];
    ele[2][11] != ele[8][11];
    ele[2][11] != ele[9][11];
    ele[2][12] != ele[10][12];
    ele[2][12] != ele[11][12];
    ele[2][12] != ele[12][12];
    ele[2][12] != ele[13][12];
    ele[2][12] != ele[14][12];
    ele[2][12] != ele[15][12];
    ele[2][12] != ele[2][13];
    ele[2][12] != ele[2][14];
    ele[2][12] != ele[2][15];
    ele[2][12] != ele[3][12];
    ele[2][12] != ele[3][13];
    ele[2][12] != ele[3][14];
    ele[2][12] != ele[3][15];
    ele[2][12] != ele[4][12];
    ele[2][12] != ele[5][12];
    ele[2][12] != ele[6][12];
    ele[2][12] != ele[7][12];
    ele[2][12] != ele[8][12];
    ele[2][12] != ele[9][12];
    ele[2][13] != ele[10][13];
    ele[2][13] != ele[11][13];
    ele[2][13] != ele[12][13];
    ele[2][13] != ele[13][13];
    ele[2][13] != ele[14][13];
    ele[2][13] != ele[15][13];
    ele[2][13] != ele[2][14];
    ele[2][13] != ele[2][15];
    ele[2][13] != ele[3][12];
    ele[2][13] != ele[3][13];
    ele[2][13] != ele[3][14];
    ele[2][13] != ele[3][15];
    ele[2][13] != ele[4][13];
    ele[2][13] != ele[5][13];
    ele[2][13] != ele[6][13];
    ele[2][13] != ele[7][13];
    ele[2][13] != ele[8][13];
    ele[2][13] != ele[9][13];
    ele[2][14] != ele[10][14];
    ele[2][14] != ele[11][14];
    ele[2][14] != ele[12][14];
    ele[2][14] != ele[13][14];
    ele[2][14] != ele[14][14];
    ele[2][14] != ele[15][14];
    ele[2][14] != ele[2][15];
    ele[2][14] != ele[3][12];
    ele[2][14] != ele[3][13];
    ele[2][14] != ele[3][14];
    ele[2][14] != ele[3][15];
    ele[2][14] != ele[4][14];
    ele[2][14] != ele[5][14];
    ele[2][14] != ele[6][14];
    ele[2][14] != ele[7][14];
    ele[2][14] != ele[8][14];
    ele[2][14] != ele[9][14];
    ele[2][15] != ele[10][15];
    ele[2][15] != ele[11][15];
    ele[2][15] != ele[12][15];
    ele[2][15] != ele[13][15];
    ele[2][15] != ele[14][15];
    ele[2][15] != ele[15][15];
    ele[2][15] != ele[3][12];
    ele[2][15] != ele[3][13];
    ele[2][15] != ele[3][14];
    ele[2][15] != ele[3][15];
    ele[2][15] != ele[4][15];
    ele[2][15] != ele[5][15];
    ele[2][15] != ele[6][15];
    ele[2][15] != ele[7][15];
    ele[2][15] != ele[8][15];
    ele[2][15] != ele[9][15];
    ele[2][2] != ele[10][2];
    ele[2][2] != ele[11][2];
    ele[2][2] != ele[12][2];
    ele[2][2] != ele[13][2];
    ele[2][2] != ele[14][2];
    ele[2][2] != ele[15][2];
    ele[2][2] != ele[2][10];
    ele[2][2] != ele[2][11];
    ele[2][2] != ele[2][12];
    ele[2][2] != ele[2][13];
    ele[2][2] != ele[2][14];
    ele[2][2] != ele[2][15];
    ele[2][2] != ele[2][3];
    ele[2][2] != ele[2][4];
    ele[2][2] != ele[2][5];
    ele[2][2] != ele[2][6];
    ele[2][2] != ele[2][7];
    ele[2][2] != ele[2][8];
    ele[2][2] != ele[2][9];
    ele[2][2] != ele[3][0];
    ele[2][2] != ele[3][1];
    ele[2][2] != ele[3][2];
    ele[2][2] != ele[3][3];
    ele[2][2] != ele[4][2];
    ele[2][2] != ele[5][2];
    ele[2][2] != ele[6][2];
    ele[2][2] != ele[7][2];
    ele[2][2] != ele[8][2];
    ele[2][2] != ele[9][2];
    ele[2][3] != ele[10][3];
    ele[2][3] != ele[11][3];
    ele[2][3] != ele[12][3];
    ele[2][3] != ele[13][3];
    ele[2][3] != ele[14][3];
    ele[2][3] != ele[15][3];
    ele[2][3] != ele[2][10];
    ele[2][3] != ele[2][11];
    ele[2][3] != ele[2][12];
    ele[2][3] != ele[2][13];
    ele[2][3] != ele[2][14];
    ele[2][3] != ele[2][15];
    ele[2][3] != ele[2][4];
    ele[2][3] != ele[2][5];
    ele[2][3] != ele[2][6];
    ele[2][3] != ele[2][7];
    ele[2][3] != ele[2][8];
    ele[2][3] != ele[2][9];
    ele[2][3] != ele[3][0];
    ele[2][3] != ele[3][1];
    ele[2][3] != ele[3][2];
    ele[2][3] != ele[3][3];
    ele[2][3] != ele[4][3];
    ele[2][3] != ele[5][3];
    ele[2][3] != ele[6][3];
    ele[2][3] != ele[7][3];
    ele[2][3] != ele[8][3];
    ele[2][3] != ele[9][3];
    ele[2][4] != ele[10][4];
    ele[2][4] != ele[11][4];
    ele[2][4] != ele[12][4];
    ele[2][4] != ele[13][4];
    ele[2][4] != ele[14][4];
    ele[2][4] != ele[15][4];
    ele[2][4] != ele[2][10];
    ele[2][4] != ele[2][11];
    ele[2][4] != ele[2][12];
    ele[2][4] != ele[2][13];
    ele[2][4] != ele[2][14];
    ele[2][4] != ele[2][15];
    ele[2][4] != ele[2][5];
    ele[2][4] != ele[2][6];
    ele[2][4] != ele[2][7];
    ele[2][4] != ele[2][8];
    ele[2][4] != ele[2][9];
    ele[2][4] != ele[3][4];
    ele[2][4] != ele[3][5];
    ele[2][4] != ele[3][6];
    ele[2][4] != ele[3][7];
    ele[2][4] != ele[4][4];
    ele[2][4] != ele[5][4];
    ele[2][4] != ele[6][4];
    ele[2][4] != ele[7][4];
    ele[2][4] != ele[8][4];
    ele[2][4] != ele[9][4];
    ele[2][5] != ele[10][5];
    ele[2][5] != ele[11][5];
    ele[2][5] != ele[12][5];
    ele[2][5] != ele[13][5];
    ele[2][5] != ele[14][5];
    ele[2][5] != ele[15][5];
    ele[2][5] != ele[2][10];
    ele[2][5] != ele[2][11];
    ele[2][5] != ele[2][12];
    ele[2][5] != ele[2][13];
    ele[2][5] != ele[2][14];
    ele[2][5] != ele[2][15];
    ele[2][5] != ele[2][6];
    ele[2][5] != ele[2][7];
    ele[2][5] != ele[2][8];
    ele[2][5] != ele[2][9];
    ele[2][5] != ele[3][4];
    ele[2][5] != ele[3][5];
    ele[2][5] != ele[3][6];
    ele[2][5] != ele[3][7];
    ele[2][5] != ele[4][5];
    ele[2][5] != ele[5][5];
    ele[2][5] != ele[6][5];
    ele[2][5] != ele[7][5];
    ele[2][5] != ele[8][5];
    ele[2][5] != ele[9][5];
    ele[2][6] != ele[10][6];
    ele[2][6] != ele[11][6];
    ele[2][6] != ele[12][6];
    ele[2][6] != ele[13][6];
    ele[2][6] != ele[14][6];
    ele[2][6] != ele[15][6];
    ele[2][6] != ele[2][10];
    ele[2][6] != ele[2][11];
    ele[2][6] != ele[2][12];
    ele[2][6] != ele[2][13];
    ele[2][6] != ele[2][14];
    ele[2][6] != ele[2][15];
    ele[2][6] != ele[2][7];
    ele[2][6] != ele[2][8];
    ele[2][6] != ele[2][9];
    ele[2][6] != ele[3][4];
    ele[2][6] != ele[3][5];
    ele[2][6] != ele[3][6];
    ele[2][6] != ele[3][7];
    ele[2][6] != ele[4][6];
    ele[2][6] != ele[5][6];
    ele[2][6] != ele[6][6];
    ele[2][6] != ele[7][6];
    ele[2][6] != ele[8][6];
    ele[2][6] != ele[9][6];
    ele[2][7] != ele[10][7];
    ele[2][7] != ele[11][7];
    ele[2][7] != ele[12][7];
    ele[2][7] != ele[13][7];
    ele[2][7] != ele[14][7];
    ele[2][7] != ele[15][7];
    ele[2][7] != ele[2][10];
    ele[2][7] != ele[2][11];
    ele[2][7] != ele[2][12];
    ele[2][7] != ele[2][13];
    ele[2][7] != ele[2][14];
    ele[2][7] != ele[2][15];
    ele[2][7] != ele[2][8];
    ele[2][7] != ele[2][9];
    ele[2][7] != ele[3][4];
    ele[2][7] != ele[3][5];
    ele[2][7] != ele[3][6];
    ele[2][7] != ele[3][7];
    ele[2][7] != ele[4][7];
    ele[2][7] != ele[5][7];
    ele[2][7] != ele[6][7];
    ele[2][7] != ele[7][7];
    ele[2][7] != ele[8][7];
    ele[2][7] != ele[9][7];
    ele[2][8] != ele[10][8];
    ele[2][8] != ele[11][8];
    ele[2][8] != ele[12][8];
    ele[2][8] != ele[13][8];
    ele[2][8] != ele[14][8];
    ele[2][8] != ele[15][8];
    ele[2][8] != ele[2][10];
    ele[2][8] != ele[2][11];
    ele[2][8] != ele[2][12];
    ele[2][8] != ele[2][13];
    ele[2][8] != ele[2][14];
    ele[2][8] != ele[2][15];
    ele[2][8] != ele[2][9];
    ele[2][8] != ele[3][10];
    ele[2][8] != ele[3][11];
    ele[2][8] != ele[3][8];
    ele[2][8] != ele[3][9];
    ele[2][8] != ele[4][8];
    ele[2][8] != ele[5][8];
    ele[2][8] != ele[6][8];
    ele[2][8] != ele[7][8];
    ele[2][8] != ele[8][8];
    ele[2][8] != ele[9][8];
    ele[2][9] != ele[10][9];
    ele[2][9] != ele[11][9];
    ele[2][9] != ele[12][9];
    ele[2][9] != ele[13][9];
    ele[2][9] != ele[14][9];
    ele[2][9] != ele[15][9];
    ele[2][9] != ele[2][10];
    ele[2][9] != ele[2][11];
    ele[2][9] != ele[2][12];
    ele[2][9] != ele[2][13];
    ele[2][9] != ele[2][14];
    ele[2][9] != ele[2][15];
    ele[2][9] != ele[3][10];
    ele[2][9] != ele[3][11];
    ele[2][9] != ele[3][8];
    ele[2][9] != ele[3][9];
    ele[2][9] != ele[4][9];
    ele[2][9] != ele[5][9];
    ele[2][9] != ele[6][9];
    ele[2][9] != ele[7][9];
    ele[2][9] != ele[8][9];
    ele[2][9] != ele[9][9];
    ele[3][0] != ele[10][0];
    ele[3][0] != ele[11][0];
    ele[3][0] != ele[12][0];
    ele[3][0] != ele[13][0];
    ele[3][0] != ele[14][0];
    ele[3][0] != ele[15][0];
    ele[3][0] != ele[3][1];
    ele[3][0] != ele[3][10];
    ele[3][0] != ele[3][11];
    ele[3][0] != ele[3][12];
    ele[3][0] != ele[3][13];
    ele[3][0] != ele[3][14];
    ele[3][0] != ele[3][15];
    ele[3][0] != ele[3][2];
    ele[3][0] != ele[3][3];
    ele[3][0] != ele[3][4];
    ele[3][0] != ele[3][5];
    ele[3][0] != ele[3][6];
    ele[3][0] != ele[3][7];
    ele[3][0] != ele[3][8];
    ele[3][0] != ele[3][9];
    ele[3][0] != ele[4][0];
    ele[3][0] != ele[5][0];
    ele[3][0] != ele[6][0];
    ele[3][0] != ele[7][0];
    ele[3][0] != ele[8][0];
    ele[3][0] != ele[9][0];
    ele[3][1] != ele[10][1];
    ele[3][1] != ele[11][1];
    ele[3][1] != ele[12][1];
    ele[3][1] != ele[13][1];
    ele[3][1] != ele[14][1];
    ele[3][1] != ele[15][1];
    ele[3][1] != ele[3][10];
    ele[3][1] != ele[3][11];
    ele[3][1] != ele[3][12];
    ele[3][1] != ele[3][13];
    ele[3][1] != ele[3][14];
    ele[3][1] != ele[3][15];
    ele[3][1] != ele[3][2];
    ele[3][1] != ele[3][3];
    ele[3][1] != ele[3][4];
    ele[3][1] != ele[3][5];
    ele[3][1] != ele[3][6];
    ele[3][1] != ele[3][7];
    ele[3][1] != ele[3][8];
    ele[3][1] != ele[3][9];
    ele[3][1] != ele[4][1];
    ele[3][1] != ele[5][1];
    ele[3][1] != ele[6][1];
    ele[3][1] != ele[7][1];
    ele[3][1] != ele[8][1];
    ele[3][1] != ele[9][1];
    ele[3][10] != ele[10][10];
    ele[3][10] != ele[11][10];
    ele[3][10] != ele[12][10];
    ele[3][10] != ele[13][10];
    ele[3][10] != ele[14][10];
    ele[3][10] != ele[15][10];
    ele[3][10] != ele[3][11];
    ele[3][10] != ele[3][12];
    ele[3][10] != ele[3][13];
    ele[3][10] != ele[3][14];
    ele[3][10] != ele[3][15];
    ele[3][10] != ele[4][10];
    ele[3][10] != ele[5][10];
    ele[3][10] != ele[6][10];
    ele[3][10] != ele[7][10];
    ele[3][10] != ele[8][10];
    ele[3][10] != ele[9][10];
    ele[3][11] != ele[10][11];
    ele[3][11] != ele[11][11];
    ele[3][11] != ele[12][11];
    ele[3][11] != ele[13][11];
    ele[3][11] != ele[14][11];
    ele[3][11] != ele[15][11];
    ele[3][11] != ele[3][12];
    ele[3][11] != ele[3][13];
    ele[3][11] != ele[3][14];
    ele[3][11] != ele[3][15];
    ele[3][11] != ele[4][11];
    ele[3][11] != ele[5][11];
    ele[3][11] != ele[6][11];
    ele[3][11] != ele[7][11];
    ele[3][11] != ele[8][11];
    ele[3][11] != ele[9][11];
    ele[3][12] != ele[10][12];
    ele[3][12] != ele[11][12];
    ele[3][12] != ele[12][12];
    ele[3][12] != ele[13][12];
    ele[3][12] != ele[14][12];
    ele[3][12] != ele[15][12];
    ele[3][12] != ele[3][13];
    ele[3][12] != ele[3][14];
    ele[3][12] != ele[3][15];
    ele[3][12] != ele[4][12];
    ele[3][12] != ele[5][12];
    ele[3][12] != ele[6][12];
    ele[3][12] != ele[7][12];
    ele[3][12] != ele[8][12];
    ele[3][12] != ele[9][12];
    ele[3][13] != ele[10][13];
    ele[3][13] != ele[11][13];
    ele[3][13] != ele[12][13];
    ele[3][13] != ele[13][13];
    ele[3][13] != ele[14][13];
    ele[3][13] != ele[15][13];
    ele[3][13] != ele[3][14];
    ele[3][13] != ele[3][15];
    ele[3][13] != ele[4][13];
    ele[3][13] != ele[5][13];
    ele[3][13] != ele[6][13];
    ele[3][13] != ele[7][13];
    ele[3][13] != ele[8][13];
    ele[3][13] != ele[9][13];
    ele[3][14] != ele[10][14];
    ele[3][14] != ele[11][14];
    ele[3][14] != ele[12][14];
    ele[3][14] != ele[13][14];
    ele[3][14] != ele[14][14];
    ele[3][14] != ele[15][14];
    ele[3][14] != ele[3][15];
    ele[3][14] != ele[4][14];
    ele[3][14] != ele[5][14];
    ele[3][14] != ele[6][14];
    ele[3][14] != ele[7][14];
    ele[3][14] != ele[8][14];
    ele[3][14] != ele[9][14];
    ele[3][15] != ele[10][15];
    ele[3][15] != ele[11][15];
    ele[3][15] != ele[12][15];
    ele[3][15] != ele[13][15];
    ele[3][15] != ele[14][15];
    ele[3][15] != ele[15][15];
    ele[3][15] != ele[4][15];
    ele[3][15] != ele[5][15];
    ele[3][15] != ele[6][15];
    ele[3][15] != ele[7][15];
    ele[3][15] != ele[8][15];
    ele[3][15] != ele[9][15];
    ele[3][2] != ele[10][2];
    ele[3][2] != ele[11][2];
    ele[3][2] != ele[12][2];
    ele[3][2] != ele[13][2];
    ele[3][2] != ele[14][2];
    ele[3][2] != ele[15][2];
    ele[3][2] != ele[3][10];
    ele[3][2] != ele[3][11];
    ele[3][2] != ele[3][12];
    ele[3][2] != ele[3][13];
    ele[3][2] != ele[3][14];
    ele[3][2] != ele[3][15];
    ele[3][2] != ele[3][3];
    ele[3][2] != ele[3][4];
    ele[3][2] != ele[3][5];
    ele[3][2] != ele[3][6];
    ele[3][2] != ele[3][7];
    ele[3][2] != ele[3][8];
    ele[3][2] != ele[3][9];
    ele[3][2] != ele[4][2];
    ele[3][2] != ele[5][2];
    ele[3][2] != ele[6][2];
    ele[3][2] != ele[7][2];
    ele[3][2] != ele[8][2];
    ele[3][2] != ele[9][2];
    ele[3][3] != ele[10][3];
    ele[3][3] != ele[11][3];
    ele[3][3] != ele[12][3];
    ele[3][3] != ele[13][3];
    ele[3][3] != ele[14][3];
    ele[3][3] != ele[15][3];
    ele[3][3] != ele[3][10];
    ele[3][3] != ele[3][11];
    ele[3][3] != ele[3][12];
    ele[3][3] != ele[3][13];
    ele[3][3] != ele[3][14];
    ele[3][3] != ele[3][15];
    ele[3][3] != ele[3][4];
    ele[3][3] != ele[3][5];
    ele[3][3] != ele[3][6];
    ele[3][3] != ele[3][7];
    ele[3][3] != ele[3][8];
    ele[3][3] != ele[3][9];
    ele[3][3] != ele[4][3];
    ele[3][3] != ele[5][3];
    ele[3][3] != ele[6][3];
    ele[3][3] != ele[7][3];
    ele[3][3] != ele[8][3];
    ele[3][3] != ele[9][3];
    ele[3][4] != ele[10][4];
    ele[3][4] != ele[11][4];
    ele[3][4] != ele[12][4];
    ele[3][4] != ele[13][4];
    ele[3][4] != ele[14][4];
    ele[3][4] != ele[15][4];
    ele[3][4] != ele[3][10];
    ele[3][4] != ele[3][11];
    ele[3][4] != ele[3][12];
    ele[3][4] != ele[3][13];
    ele[3][4] != ele[3][14];
    ele[3][4] != ele[3][15];
    ele[3][4] != ele[3][5];
    ele[3][4] != ele[3][6];
    ele[3][4] != ele[3][7];
    ele[3][4] != ele[3][8];
    ele[3][4] != ele[3][9];
    ele[3][4] != ele[4][4];
    ele[3][4] != ele[5][4];
    ele[3][4] != ele[6][4];
    ele[3][4] != ele[7][4];
    ele[3][4] != ele[8][4];
    ele[3][4] != ele[9][4];
    ele[3][5] != ele[10][5];
    ele[3][5] != ele[11][5];
    ele[3][5] != ele[12][5];
    ele[3][5] != ele[13][5];
    ele[3][5] != ele[14][5];
    ele[3][5] != ele[15][5];
    ele[3][5] != ele[3][10];
    ele[3][5] != ele[3][11];
    ele[3][5] != ele[3][12];
    ele[3][5] != ele[3][13];
    ele[3][5] != ele[3][14];
    ele[3][5] != ele[3][15];
    ele[3][5] != ele[3][6];
    ele[3][5] != ele[3][7];
    ele[3][5] != ele[3][8];
    ele[3][5] != ele[3][9];
    ele[3][5] != ele[4][5];
    ele[3][5] != ele[5][5];
    ele[3][5] != ele[6][5];
    ele[3][5] != ele[7][5];
    ele[3][5] != ele[8][5];
    ele[3][5] != ele[9][5];
    ele[3][6] != ele[10][6];
    ele[3][6] != ele[11][6];
    ele[3][6] != ele[12][6];
    ele[3][6] != ele[13][6];
    ele[3][6] != ele[14][6];
    ele[3][6] != ele[15][6];
    ele[3][6] != ele[3][10];
    ele[3][6] != ele[3][11];
    ele[3][6] != ele[3][12];
    ele[3][6] != ele[3][13];
    ele[3][6] != ele[3][14];
    ele[3][6] != ele[3][15];
    ele[3][6] != ele[3][7];
    ele[3][6] != ele[3][8];
    ele[3][6] != ele[3][9];
    ele[3][6] != ele[4][6];
    ele[3][6] != ele[5][6];
    ele[3][6] != ele[6][6];
    ele[3][6] != ele[7][6];
    ele[3][6] != ele[8][6];
    ele[3][6] != ele[9][6];
    ele[3][7] != ele[10][7];
    ele[3][7] != ele[11][7];
    ele[3][7] != ele[12][7];
    ele[3][7] != ele[13][7];
    ele[3][7] != ele[14][7];
    ele[3][7] != ele[15][7];
    ele[3][7] != ele[3][10];
    ele[3][7] != ele[3][11];
    ele[3][7] != ele[3][12];
    ele[3][7] != ele[3][13];
    ele[3][7] != ele[3][14];
    ele[3][7] != ele[3][15];
    ele[3][7] != ele[3][8];
    ele[3][7] != ele[3][9];
    ele[3][7] != ele[4][7];
    ele[3][7] != ele[5][7];
    ele[3][7] != ele[6][7];
    ele[3][7] != ele[7][7];
    ele[3][7] != ele[8][7];
    ele[3][7] != ele[9][7];
    ele[3][8] != ele[10][8];
    ele[3][8] != ele[11][8];
    ele[3][8] != ele[12][8];
    ele[3][8] != ele[13][8];
    ele[3][8] != ele[14][8];
    ele[3][8] != ele[15][8];
    ele[3][8] != ele[3][10];
    ele[3][8] != ele[3][11];
    ele[3][8] != ele[3][12];
    ele[3][8] != ele[3][13];
    ele[3][8] != ele[3][14];
    ele[3][8] != ele[3][15];
    ele[3][8] != ele[3][9];
    ele[3][8] != ele[4][8];
    ele[3][8] != ele[5][8];
    ele[3][8] != ele[6][8];
    ele[3][8] != ele[7][8];
    ele[3][8] != ele[8][8];
    ele[3][8] != ele[9][8];
    ele[3][9] != ele[10][9];
    ele[3][9] != ele[11][9];
    ele[3][9] != ele[12][9];
    ele[3][9] != ele[13][9];
    ele[3][9] != ele[14][9];
    ele[3][9] != ele[15][9];
    ele[3][9] != ele[3][10];
    ele[3][9] != ele[3][11];
    ele[3][9] != ele[3][12];
    ele[3][9] != ele[3][13];
    ele[3][9] != ele[3][14];
    ele[3][9] != ele[3][15];
    ele[3][9] != ele[4][9];
    ele[3][9] != ele[5][9];
    ele[3][9] != ele[6][9];
    ele[3][9] != ele[7][9];
    ele[3][9] != ele[8][9];
    ele[3][9] != ele[9][9];
    ele[4][0] != ele[10][0];
    ele[4][0] != ele[11][0];
    ele[4][0] != ele[12][0];
    ele[4][0] != ele[13][0];
    ele[4][0] != ele[14][0];
    ele[4][0] != ele[15][0];
    ele[4][0] != ele[4][1];
    ele[4][0] != ele[4][10];
    ele[4][0] != ele[4][11];
    ele[4][0] != ele[4][12];
    ele[4][0] != ele[4][13];
    ele[4][0] != ele[4][14];
    ele[4][0] != ele[4][15];
    ele[4][0] != ele[4][2];
    ele[4][0] != ele[4][3];
    ele[4][0] != ele[4][4];
    ele[4][0] != ele[4][5];
    ele[4][0] != ele[4][6];
    ele[4][0] != ele[4][7];
    ele[4][0] != ele[4][8];
    ele[4][0] != ele[4][9];
    ele[4][0] != ele[5][0];
    ele[4][0] != ele[5][1];
    ele[4][0] != ele[5][2];
    ele[4][0] != ele[5][3];
    ele[4][0] != ele[6][0];
    ele[4][0] != ele[6][1];
    ele[4][0] != ele[6][2];
    ele[4][0] != ele[6][3];
    ele[4][0] != ele[7][0];
    ele[4][0] != ele[7][1];
    ele[4][0] != ele[7][2];
    ele[4][0] != ele[7][3];
    ele[4][0] != ele[8][0];
    ele[4][0] != ele[9][0];
    ele[4][1] != ele[10][1];
    ele[4][1] != ele[11][1];
    ele[4][1] != ele[12][1];
    ele[4][1] != ele[13][1];
    ele[4][1] != ele[14][1];
    ele[4][1] != ele[15][1];
    ele[4][1] != ele[4][10];
    ele[4][1] != ele[4][11];
    ele[4][1] != ele[4][12];
    ele[4][1] != ele[4][13];
    ele[4][1] != ele[4][14];
    ele[4][1] != ele[4][15];
    ele[4][1] != ele[4][2];
    ele[4][1] != ele[4][3];
    ele[4][1] != ele[4][4];
    ele[4][1] != ele[4][5];
    ele[4][1] != ele[4][6];
    ele[4][1] != ele[4][7];
    ele[4][1] != ele[4][8];
    ele[4][1] != ele[4][9];
    ele[4][1] != ele[5][0];
    ele[4][1] != ele[5][1];
    ele[4][1] != ele[5][2];
    ele[4][1] != ele[5][3];
    ele[4][1] != ele[6][0];
    ele[4][1] != ele[6][1];
    ele[4][1] != ele[6][2];
    ele[4][1] != ele[6][3];
    ele[4][1] != ele[7][0];
    ele[4][1] != ele[7][1];
    ele[4][1] != ele[7][2];
    ele[4][1] != ele[7][3];
    ele[4][1] != ele[8][1];
    ele[4][1] != ele[9][1];
    ele[4][10] != ele[10][10];
    ele[4][10] != ele[11][10];
    ele[4][10] != ele[12][10];
    ele[4][10] != ele[13][10];
    ele[4][10] != ele[14][10];
    ele[4][10] != ele[15][10];
    ele[4][10] != ele[4][11];
    ele[4][10] != ele[4][12];
    ele[4][10] != ele[4][13];
    ele[4][10] != ele[4][14];
    ele[4][10] != ele[4][15];
    ele[4][10] != ele[5][10];
    ele[4][10] != ele[5][11];
    ele[4][10] != ele[5][8];
    ele[4][10] != ele[5][9];
    ele[4][10] != ele[6][10];
    ele[4][10] != ele[6][11];
    ele[4][10] != ele[6][8];
    ele[4][10] != ele[6][9];
    ele[4][10] != ele[7][10];
    ele[4][10] != ele[7][11];
    ele[4][10] != ele[7][8];
    ele[4][10] != ele[7][9];
    ele[4][10] != ele[8][10];
    ele[4][10] != ele[9][10];
    ele[4][11] != ele[10][11];
    ele[4][11] != ele[11][11];
    ele[4][11] != ele[12][11];
    ele[4][11] != ele[13][11];
    ele[4][11] != ele[14][11];
    ele[4][11] != ele[15][11];
    ele[4][11] != ele[4][12];
    ele[4][11] != ele[4][13];
    ele[4][11] != ele[4][14];
    ele[4][11] != ele[4][15];
    ele[4][11] != ele[5][10];
    ele[4][11] != ele[5][11];
    ele[4][11] != ele[5][8];
    ele[4][11] != ele[5][9];
    ele[4][11] != ele[6][10];
    ele[4][11] != ele[6][11];
    ele[4][11] != ele[6][8];
    ele[4][11] != ele[6][9];
    ele[4][11] != ele[7][10];
    ele[4][11] != ele[7][11];
    ele[4][11] != ele[7][8];
    ele[4][11] != ele[7][9];
    ele[4][11] != ele[8][11];
    ele[4][11] != ele[9][11];
    ele[4][12] != ele[10][12];
    ele[4][12] != ele[11][12];
    ele[4][12] != ele[12][12];
    ele[4][12] != ele[13][12];
    ele[4][12] != ele[14][12];
    ele[4][12] != ele[15][12];
    ele[4][12] != ele[4][13];
    ele[4][12] != ele[4][14];
    ele[4][12] != ele[4][15];
    ele[4][12] != ele[5][12];
    ele[4][12] != ele[5][13];
    ele[4][12] != ele[5][14];
    ele[4][12] != ele[5][15];
    ele[4][12] != ele[6][12];
    ele[4][12] != ele[6][13];
    ele[4][12] != ele[6][14];
    ele[4][12] != ele[6][15];
    ele[4][12] != ele[7][12];
    ele[4][12] != ele[7][13];
    ele[4][12] != ele[7][14];
    ele[4][12] != ele[7][15];
    ele[4][12] != ele[8][12];
    ele[4][12] != ele[9][12];
    ele[4][13] != ele[10][13];
    ele[4][13] != ele[11][13];
    ele[4][13] != ele[12][13];
    ele[4][13] != ele[13][13];
    ele[4][13] != ele[14][13];
    ele[4][13] != ele[15][13];
    ele[4][13] != ele[4][14];
    ele[4][13] != ele[4][15];
    ele[4][13] != ele[5][12];
    ele[4][13] != ele[5][13];
    ele[4][13] != ele[5][14];
    ele[4][13] != ele[5][15];
    ele[4][13] != ele[6][12];
    ele[4][13] != ele[6][13];
    ele[4][13] != ele[6][14];
    ele[4][13] != ele[6][15];
    ele[4][13] != ele[7][12];
    ele[4][13] != ele[7][13];
    ele[4][13] != ele[7][14];
    ele[4][13] != ele[7][15];
    ele[4][13] != ele[8][13];
    ele[4][13] != ele[9][13];
    ele[4][14] != ele[10][14];
    ele[4][14] != ele[11][14];
    ele[4][14] != ele[12][14];
    ele[4][14] != ele[13][14];
    ele[4][14] != ele[14][14];
    ele[4][14] != ele[15][14];
    ele[4][14] != ele[4][15];
    ele[4][14] != ele[5][12];
    ele[4][14] != ele[5][13];
    ele[4][14] != ele[5][14];
    ele[4][14] != ele[5][15];
    ele[4][14] != ele[6][12];
    ele[4][14] != ele[6][13];
    ele[4][14] != ele[6][14];
    ele[4][14] != ele[6][15];
    ele[4][14] != ele[7][12];
    ele[4][14] != ele[7][13];
    ele[4][14] != ele[7][14];
    ele[4][14] != ele[7][15];
    ele[4][14] != ele[8][14];
    ele[4][14] != ele[9][14];
    ele[4][15] != ele[10][15];
    ele[4][15] != ele[11][15];
    ele[4][15] != ele[12][15];
    ele[4][15] != ele[13][15];
    ele[4][15] != ele[14][15];
    ele[4][15] != ele[15][15];
    ele[4][15] != ele[5][12];
    ele[4][15] != ele[5][13];
    ele[4][15] != ele[5][14];
    ele[4][15] != ele[5][15];
    ele[4][15] != ele[6][12];
    ele[4][15] != ele[6][13];
    ele[4][15] != ele[6][14];
    ele[4][15] != ele[6][15];
    ele[4][15] != ele[7][12];
    ele[4][15] != ele[7][13];
    ele[4][15] != ele[7][14];
    ele[4][15] != ele[7][15];
    ele[4][15] != ele[8][15];
    ele[4][15] != ele[9][15];
    ele[4][2] != ele[10][2];
    ele[4][2] != ele[11][2];
    ele[4][2] != ele[12][2];
    ele[4][2] != ele[13][2];
    ele[4][2] != ele[14][2];
    ele[4][2] != ele[15][2];
    ele[4][2] != ele[4][10];
    ele[4][2] != ele[4][11];
    ele[4][2] != ele[4][12];
    ele[4][2] != ele[4][13];
    ele[4][2] != ele[4][14];
    ele[4][2] != ele[4][15];
    ele[4][2] != ele[4][3];
    ele[4][2] != ele[4][4];
    ele[4][2] != ele[4][5];
    ele[4][2] != ele[4][6];
    ele[4][2] != ele[4][7];
    ele[4][2] != ele[4][8];
    ele[4][2] != ele[4][9];
    ele[4][2] != ele[5][0];
    ele[4][2] != ele[5][1];
    ele[4][2] != ele[5][2];
    ele[4][2] != ele[5][3];
    ele[4][2] != ele[6][0];
    ele[4][2] != ele[6][1];
    ele[4][2] != ele[6][2];
    ele[4][2] != ele[6][3];
    ele[4][2] != ele[7][0];
    ele[4][2] != ele[7][1];
    ele[4][2] != ele[7][2];
    ele[4][2] != ele[7][3];
    ele[4][2] != ele[8][2];
    ele[4][2] != ele[9][2];
    ele[4][3] != ele[10][3];
    ele[4][3] != ele[11][3];
    ele[4][3] != ele[12][3];
    ele[4][3] != ele[13][3];
    ele[4][3] != ele[14][3];
    ele[4][3] != ele[15][3];
    ele[4][3] != ele[4][10];
    ele[4][3] != ele[4][11];
    ele[4][3] != ele[4][12];
    ele[4][3] != ele[4][13];
    ele[4][3] != ele[4][14];
    ele[4][3] != ele[4][15];
    ele[4][3] != ele[4][4];
    ele[4][3] != ele[4][5];
    ele[4][3] != ele[4][6];
    ele[4][3] != ele[4][7];
    ele[4][3] != ele[4][8];
    ele[4][3] != ele[4][9];
    ele[4][3] != ele[5][0];
    ele[4][3] != ele[5][1];
    ele[4][3] != ele[5][2];
    ele[4][3] != ele[5][3];
    ele[4][3] != ele[6][0];
    ele[4][3] != ele[6][1];
    ele[4][3] != ele[6][2];
    ele[4][3] != ele[6][3];
    ele[4][3] != ele[7][0];
    ele[4][3] != ele[7][1];
    ele[4][3] != ele[7][2];
    ele[4][3] != ele[7][3];
    ele[4][3] != ele[8][3];
    ele[4][3] != ele[9][3];
    ele[4][4] != ele[10][4];
    ele[4][4] != ele[11][4];
    ele[4][4] != ele[12][4];
    ele[4][4] != ele[13][4];
    ele[4][4] != ele[14][4];
    ele[4][4] != ele[15][4];
    ele[4][4] != ele[4][10];
    ele[4][4] != ele[4][11];
    ele[4][4] != ele[4][12];
    ele[4][4] != ele[4][13];
    ele[4][4] != ele[4][14];
    ele[4][4] != ele[4][15];
    ele[4][4] != ele[4][5];
    ele[4][4] != ele[4][6];
    ele[4][4] != ele[4][7];
    ele[4][4] != ele[4][8];
    ele[4][4] != ele[4][9];
    ele[4][4] != ele[5][4];
    ele[4][4] != ele[5][5];
    ele[4][4] != ele[5][6];
    ele[4][4] != ele[5][7];
    ele[4][4] != ele[6][4];
    ele[4][4] != ele[6][5];
    ele[4][4] != ele[6][6];
    ele[4][4] != ele[6][7];
    ele[4][4] != ele[7][4];
    ele[4][4] != ele[7][5];
    ele[4][4] != ele[7][6];
    ele[4][4] != ele[7][7];
    ele[4][4] != ele[8][4];
    ele[4][4] != ele[9][4];
    ele[4][5] != ele[10][5];
    ele[4][5] != ele[11][5];
    ele[4][5] != ele[12][5];
    ele[4][5] != ele[13][5];
    ele[4][5] != ele[14][5];
    ele[4][5] != ele[15][5];
    ele[4][5] != ele[4][10];
    ele[4][5] != ele[4][11];
    ele[4][5] != ele[4][12];
    ele[4][5] != ele[4][13];
    ele[4][5] != ele[4][14];
    ele[4][5] != ele[4][15];
    ele[4][5] != ele[4][6];
    ele[4][5] != ele[4][7];
    ele[4][5] != ele[4][8];
    ele[4][5] != ele[4][9];
    ele[4][5] != ele[5][4];
    ele[4][5] != ele[5][5];
    ele[4][5] != ele[5][6];
    ele[4][5] != ele[5][7];
    ele[4][5] != ele[6][4];
    ele[4][5] != ele[6][5];
    ele[4][5] != ele[6][6];
    ele[4][5] != ele[6][7];
    ele[4][5] != ele[7][4];
    ele[4][5] != ele[7][5];
    ele[4][5] != ele[7][6];
    ele[4][5] != ele[7][7];
    ele[4][5] != ele[8][5];
    ele[4][5] != ele[9][5];
    ele[4][6] != ele[10][6];
    ele[4][6] != ele[11][6];
    ele[4][6] != ele[12][6];
    ele[4][6] != ele[13][6];
    ele[4][6] != ele[14][6];
    ele[4][6] != ele[15][6];
    ele[4][6] != ele[4][10];
    ele[4][6] != ele[4][11];
    ele[4][6] != ele[4][12];
    ele[4][6] != ele[4][13];
    ele[4][6] != ele[4][14];
    ele[4][6] != ele[4][15];
    ele[4][6] != ele[4][7];
    ele[4][6] != ele[4][8];
    ele[4][6] != ele[4][9];
    ele[4][6] != ele[5][4];
    ele[4][6] != ele[5][5];
    ele[4][6] != ele[5][6];
    ele[4][6] != ele[5][7];
    ele[4][6] != ele[6][4];
    ele[4][6] != ele[6][5];
    ele[4][6] != ele[6][6];
    ele[4][6] != ele[6][7];
    ele[4][6] != ele[7][4];
    ele[4][6] != ele[7][5];
    ele[4][6] != ele[7][6];
    ele[4][6] != ele[7][7];
    ele[4][6] != ele[8][6];
    ele[4][6] != ele[9][6];
    ele[4][7] != ele[10][7];
    ele[4][7] != ele[11][7];
    ele[4][7] != ele[12][7];
    ele[4][7] != ele[13][7];
    ele[4][7] != ele[14][7];
    ele[4][7] != ele[15][7];
    ele[4][7] != ele[4][10];
    ele[4][7] != ele[4][11];
    ele[4][7] != ele[4][12];
    ele[4][7] != ele[4][13];
    ele[4][7] != ele[4][14];
    ele[4][7] != ele[4][15];
    ele[4][7] != ele[4][8];
    ele[4][7] != ele[4][9];
    ele[4][7] != ele[5][4];
    ele[4][7] != ele[5][5];
    ele[4][7] != ele[5][6];
    ele[4][7] != ele[5][7];
    ele[4][7] != ele[6][4];
    ele[4][7] != ele[6][5];
    ele[4][7] != ele[6][6];
    ele[4][7] != ele[6][7];
    ele[4][7] != ele[7][4];
    ele[4][7] != ele[7][5];
    ele[4][7] != ele[7][6];
    ele[4][7] != ele[7][7];
    ele[4][7] != ele[8][7];
    ele[4][7] != ele[9][7];
    ele[4][8] != ele[10][8];
    ele[4][8] != ele[11][8];
    ele[4][8] != ele[12][8];
    ele[4][8] != ele[13][8];
    ele[4][8] != ele[14][8];
    ele[4][8] != ele[15][8];
    ele[4][8] != ele[4][10];
    ele[4][8] != ele[4][11];
    ele[4][8] != ele[4][12];
    ele[4][8] != ele[4][13];
    ele[4][8] != ele[4][14];
    ele[4][8] != ele[4][15];
    ele[4][8] != ele[4][9];
    ele[4][8] != ele[5][10];
    ele[4][8] != ele[5][11];
    ele[4][8] != ele[5][8];
    ele[4][8] != ele[5][9];
    ele[4][8] != ele[6][10];
    ele[4][8] != ele[6][11];
    ele[4][8] != ele[6][8];
    ele[4][8] != ele[6][9];
    ele[4][8] != ele[7][10];
    ele[4][8] != ele[7][11];
    ele[4][8] != ele[7][8];
    ele[4][8] != ele[7][9];
    ele[4][8] != ele[8][8];
    ele[4][8] != ele[9][8];
    ele[4][9] != ele[10][9];
    ele[4][9] != ele[11][9];
    ele[4][9] != ele[12][9];
    ele[4][9] != ele[13][9];
    ele[4][9] != ele[14][9];
    ele[4][9] != ele[15][9];
    ele[4][9] != ele[4][10];
    ele[4][9] != ele[4][11];
    ele[4][9] != ele[4][12];
    ele[4][9] != ele[4][13];
    ele[4][9] != ele[4][14];
    ele[4][9] != ele[4][15];
    ele[4][9] != ele[5][10];
    ele[4][9] != ele[5][11];
    ele[4][9] != ele[5][8];
    ele[4][9] != ele[5][9];
    ele[4][9] != ele[6][10];
    ele[4][9] != ele[6][11];
    ele[4][9] != ele[6][8];
    ele[4][9] != ele[6][9];
    ele[4][9] != ele[7][10];
    ele[4][9] != ele[7][11];
    ele[4][9] != ele[7][8];
    ele[4][9] != ele[7][9];
    ele[4][9] != ele[8][9];
    ele[4][9] != ele[9][9];
    ele[5][0] != ele[10][0];
    ele[5][0] != ele[11][0];
    ele[5][0] != ele[12][0];
    ele[5][0] != ele[13][0];
    ele[5][0] != ele[14][0];
    ele[5][0] != ele[15][0];
    ele[5][0] != ele[5][1];
    ele[5][0] != ele[5][10];
    ele[5][0] != ele[5][11];
    ele[5][0] != ele[5][12];
    ele[5][0] != ele[5][13];
    ele[5][0] != ele[5][14];
    ele[5][0] != ele[5][15];
    ele[5][0] != ele[5][2];
    ele[5][0] != ele[5][3];
    ele[5][0] != ele[5][4];
    ele[5][0] != ele[5][5];
    ele[5][0] != ele[5][6];
    ele[5][0] != ele[5][7];
    ele[5][0] != ele[5][8];
    ele[5][0] != ele[5][9];
    ele[5][0] != ele[6][0];
    ele[5][0] != ele[6][1];
    ele[5][0] != ele[6][2];
    ele[5][0] != ele[6][3];
    ele[5][0] != ele[7][0];
    ele[5][0] != ele[7][1];
    ele[5][0] != ele[7][2];
    ele[5][0] != ele[7][3];
    ele[5][0] != ele[8][0];
    ele[5][0] != ele[9][0];
    ele[5][1] != ele[10][1];
    ele[5][1] != ele[11][1];
    ele[5][1] != ele[12][1];
    ele[5][1] != ele[13][1];
    ele[5][1] != ele[14][1];
    ele[5][1] != ele[15][1];
    ele[5][1] != ele[5][10];
    ele[5][1] != ele[5][11];
    ele[5][1] != ele[5][12];
    ele[5][1] != ele[5][13];
    ele[5][1] != ele[5][14];
    ele[5][1] != ele[5][15];
    ele[5][1] != ele[5][2];
    ele[5][1] != ele[5][3];
    ele[5][1] != ele[5][4];
    ele[5][1] != ele[5][5];
    ele[5][1] != ele[5][6];
    ele[5][1] != ele[5][7];
    ele[5][1] != ele[5][8];
    ele[5][1] != ele[5][9];
    ele[5][1] != ele[6][0];
    ele[5][1] != ele[6][1];
    ele[5][1] != ele[6][2];
    ele[5][1] != ele[6][3];
    ele[5][1] != ele[7][0];
    ele[5][1] != ele[7][1];
    ele[5][1] != ele[7][2];
    ele[5][1] != ele[7][3];
    ele[5][1] != ele[8][1];
    ele[5][1] != ele[9][1];
    ele[5][10] != ele[10][10];
    ele[5][10] != ele[11][10];
    ele[5][10] != ele[12][10];
    ele[5][10] != ele[13][10];
    ele[5][10] != ele[14][10];
    ele[5][10] != ele[15][10];
    ele[5][10] != ele[5][11];
    ele[5][10] != ele[5][12];
    ele[5][10] != ele[5][13];
    ele[5][10] != ele[5][14];
    ele[5][10] != ele[5][15];
    ele[5][10] != ele[6][10];
    ele[5][10] != ele[6][11];
    ele[5][10] != ele[6][8];
    ele[5][10] != ele[6][9];
    ele[5][10] != ele[7][10];
    ele[5][10] != ele[7][11];
    ele[5][10] != ele[7][8];
    ele[5][10] != ele[7][9];
    ele[5][10] != ele[8][10];
    ele[5][10] != ele[9][10];
    ele[5][11] != ele[10][11];
    ele[5][11] != ele[11][11];
    ele[5][11] != ele[12][11];
    ele[5][11] != ele[13][11];
    ele[5][11] != ele[14][11];
    ele[5][11] != ele[15][11];
    ele[5][11] != ele[5][12];
    ele[5][11] != ele[5][13];
    ele[5][11] != ele[5][14];
    ele[5][11] != ele[5][15];
    ele[5][11] != ele[6][10];
    ele[5][11] != ele[6][11];
    ele[5][11] != ele[6][8];
    ele[5][11] != ele[6][9];
    ele[5][11] != ele[7][10];
    ele[5][11] != ele[7][11];
    ele[5][11] != ele[7][8];
    ele[5][11] != ele[7][9];
    ele[5][11] != ele[8][11];
    ele[5][11] != ele[9][11];
    ele[5][12] != ele[10][12];
    ele[5][12] != ele[11][12];
    ele[5][12] != ele[12][12];
    ele[5][12] != ele[13][12];
    ele[5][12] != ele[14][12];
    ele[5][12] != ele[15][12];
    ele[5][12] != ele[5][13];
    ele[5][12] != ele[5][14];
    ele[5][12] != ele[5][15];
    ele[5][12] != ele[6][12];
    ele[5][12] != ele[6][13];
    ele[5][12] != ele[6][14];
    ele[5][12] != ele[6][15];
    ele[5][12] != ele[7][12];
    ele[5][12] != ele[7][13];
    ele[5][12] != ele[7][14];
    ele[5][12] != ele[7][15];
    ele[5][12] != ele[8][12];
    ele[5][12] != ele[9][12];
    ele[5][13] != ele[10][13];
    ele[5][13] != ele[11][13];
    ele[5][13] != ele[12][13];
    ele[5][13] != ele[13][13];
    ele[5][13] != ele[14][13];
    ele[5][13] != ele[15][13];
    ele[5][13] != ele[5][14];
    ele[5][13] != ele[5][15];
    ele[5][13] != ele[6][12];
    ele[5][13] != ele[6][13];
    ele[5][13] != ele[6][14];
    ele[5][13] != ele[6][15];
    ele[5][13] != ele[7][12];
    ele[5][13] != ele[7][13];
    ele[5][13] != ele[7][14];
    ele[5][13] != ele[7][15];
    ele[5][13] != ele[8][13];
    ele[5][13] != ele[9][13];
    ele[5][14] != ele[10][14];
    ele[5][14] != ele[11][14];
    ele[5][14] != ele[12][14];
    ele[5][14] != ele[13][14];
    ele[5][14] != ele[14][14];
    ele[5][14] != ele[15][14];
    ele[5][14] != ele[5][15];
    ele[5][14] != ele[6][12];
    ele[5][14] != ele[6][13];
    ele[5][14] != ele[6][14];
    ele[5][14] != ele[6][15];
    ele[5][14] != ele[7][12];
    ele[5][14] != ele[7][13];
    ele[5][14] != ele[7][14];
    ele[5][14] != ele[7][15];
    ele[5][14] != ele[8][14];
    ele[5][14] != ele[9][14];
    ele[5][15] != ele[10][15];
    ele[5][15] != ele[11][15];
    ele[5][15] != ele[12][15];
    ele[5][15] != ele[13][15];
    ele[5][15] != ele[14][15];
    ele[5][15] != ele[15][15];
    ele[5][15] != ele[6][12];
    ele[5][15] != ele[6][13];
    ele[5][15] != ele[6][14];
    ele[5][15] != ele[6][15];
    ele[5][15] != ele[7][12];
    ele[5][15] != ele[7][13];
    ele[5][15] != ele[7][14];
    ele[5][15] != ele[7][15];
    ele[5][15] != ele[8][15];
    ele[5][15] != ele[9][15];
    ele[5][2] != ele[10][2];
    ele[5][2] != ele[11][2];
    ele[5][2] != ele[12][2];
    ele[5][2] != ele[13][2];
    ele[5][2] != ele[14][2];
    ele[5][2] != ele[15][2];
    ele[5][2] != ele[5][10];
    ele[5][2] != ele[5][11];
    ele[5][2] != ele[5][12];
    ele[5][2] != ele[5][13];
    ele[5][2] != ele[5][14];
    ele[5][2] != ele[5][15];
    ele[5][2] != ele[5][3];
    ele[5][2] != ele[5][4];
    ele[5][2] != ele[5][5];
    ele[5][2] != ele[5][6];
    ele[5][2] != ele[5][7];
    ele[5][2] != ele[5][8];
    ele[5][2] != ele[5][9];
    ele[5][2] != ele[6][0];
    ele[5][2] != ele[6][1];
    ele[5][2] != ele[6][2];
    ele[5][2] != ele[6][3];
    ele[5][2] != ele[7][0];
    ele[5][2] != ele[7][1];
    ele[5][2] != ele[7][2];
    ele[5][2] != ele[7][3];
    ele[5][2] != ele[8][2];
    ele[5][2] != ele[9][2];
    ele[5][3] != ele[10][3];
    ele[5][3] != ele[11][3];
    ele[5][3] != ele[12][3];
    ele[5][3] != ele[13][3];
    ele[5][3] != ele[14][3];
    ele[5][3] != ele[15][3];
    ele[5][3] != ele[5][10];
    ele[5][3] != ele[5][11];
    ele[5][3] != ele[5][12];
    ele[5][3] != ele[5][13];
    ele[5][3] != ele[5][14];
    ele[5][3] != ele[5][15];
    ele[5][3] != ele[5][4];
    ele[5][3] != ele[5][5];
    ele[5][3] != ele[5][6];
    ele[5][3] != ele[5][7];
    ele[5][3] != ele[5][8];
    ele[5][3] != ele[5][9];
    ele[5][3] != ele[6][0];
    ele[5][3] != ele[6][1];
    ele[5][3] != ele[6][2];
    ele[5][3] != ele[6][3];
    ele[5][3] != ele[7][0];
    ele[5][3] != ele[7][1];
    ele[5][3] != ele[7][2];
    ele[5][3] != ele[7][3];
    ele[5][3] != ele[8][3];
    ele[5][3] != ele[9][3];
    ele[5][4] != ele[10][4];
    ele[5][4] != ele[11][4];
    ele[5][4] != ele[12][4];
    ele[5][4] != ele[13][4];
    ele[5][4] != ele[14][4];
    ele[5][4] != ele[15][4];
    ele[5][4] != ele[5][10];
    ele[5][4] != ele[5][11];
    ele[5][4] != ele[5][12];
    ele[5][4] != ele[5][13];
    ele[5][4] != ele[5][14];
    ele[5][4] != ele[5][15];
    ele[5][4] != ele[5][5];
    ele[5][4] != ele[5][6];
    ele[5][4] != ele[5][7];
    ele[5][4] != ele[5][8];
    ele[5][4] != ele[5][9];
    ele[5][4] != ele[6][4];
    ele[5][4] != ele[6][5];
    ele[5][4] != ele[6][6];
    ele[5][4] != ele[6][7];
    ele[5][4] != ele[7][4];
    ele[5][4] != ele[7][5];
    ele[5][4] != ele[7][6];
    ele[5][4] != ele[7][7];
    ele[5][4] != ele[8][4];
    ele[5][4] != ele[9][4];
    ele[5][5] != ele[10][5];
    ele[5][5] != ele[11][5];
    ele[5][5] != ele[12][5];
    ele[5][5] != ele[13][5];
    ele[5][5] != ele[14][5];
    ele[5][5] != ele[15][5];
    ele[5][5] != ele[5][10];
    ele[5][5] != ele[5][11];
    ele[5][5] != ele[5][12];
    ele[5][5] != ele[5][13];
    ele[5][5] != ele[5][14];
    ele[5][5] != ele[5][15];
    ele[5][5] != ele[5][6];
    ele[5][5] != ele[5][7];
    ele[5][5] != ele[5][8];
    ele[5][5] != ele[5][9];
    ele[5][5] != ele[6][4];
    ele[5][5] != ele[6][5];
    ele[5][5] != ele[6][6];
    ele[5][5] != ele[6][7];
    ele[5][5] != ele[7][4];
    ele[5][5] != ele[7][5];
    ele[5][5] != ele[7][6];
    ele[5][5] != ele[7][7];
    ele[5][5] != ele[8][5];
    ele[5][5] != ele[9][5];
    ele[5][6] != ele[10][6];
    ele[5][6] != ele[11][6];
    ele[5][6] != ele[12][6];
    ele[5][6] != ele[13][6];
    ele[5][6] != ele[14][6];
    ele[5][6] != ele[15][6];
    ele[5][6] != ele[5][10];
    ele[5][6] != ele[5][11];
    ele[5][6] != ele[5][12];
    ele[5][6] != ele[5][13];
    ele[5][6] != ele[5][14];
    ele[5][6] != ele[5][15];
    ele[5][6] != ele[5][7];
    ele[5][6] != ele[5][8];
    ele[5][6] != ele[5][9];
    ele[5][6] != ele[6][4];
    ele[5][6] != ele[6][5];
    ele[5][6] != ele[6][6];
    ele[5][6] != ele[6][7];
    ele[5][6] != ele[7][4];
    ele[5][6] != ele[7][5];
    ele[5][6] != ele[7][6];
    ele[5][6] != ele[7][7];
    ele[5][6] != ele[8][6];
    ele[5][6] != ele[9][6];
    ele[5][7] != ele[10][7];
    ele[5][7] != ele[11][7];
    ele[5][7] != ele[12][7];
    ele[5][7] != ele[13][7];
    ele[5][7] != ele[14][7];
    ele[5][7] != ele[15][7];
    ele[5][7] != ele[5][10];
    ele[5][7] != ele[5][11];
    ele[5][7] != ele[5][12];
    ele[5][7] != ele[5][13];
    ele[5][7] != ele[5][14];
    ele[5][7] != ele[5][15];
    ele[5][7] != ele[5][8];
    ele[5][7] != ele[5][9];
    ele[5][7] != ele[6][4];
    ele[5][7] != ele[6][5];
    ele[5][7] != ele[6][6];
    ele[5][7] != ele[6][7];
    ele[5][7] != ele[7][4];
    ele[5][7] != ele[7][5];
    ele[5][7] != ele[7][6];
    ele[5][7] != ele[7][7];
    ele[5][7] != ele[8][7];
    ele[5][7] != ele[9][7];
    ele[5][8] != ele[10][8];
    ele[5][8] != ele[11][8];
    ele[5][8] != ele[12][8];
    ele[5][8] != ele[13][8];
    ele[5][8] != ele[14][8];
    ele[5][8] != ele[15][8];
    ele[5][8] != ele[5][10];
    ele[5][8] != ele[5][11];
    ele[5][8] != ele[5][12];
    ele[5][8] != ele[5][13];
    ele[5][8] != ele[5][14];
    ele[5][8] != ele[5][15];
    ele[5][8] != ele[5][9];
    ele[5][8] != ele[6][10];
    ele[5][8] != ele[6][11];
    ele[5][8] != ele[6][8];
    ele[5][8] != ele[6][9];
    ele[5][8] != ele[7][10];
    ele[5][8] != ele[7][11];
    ele[5][8] != ele[7][8];
    ele[5][8] != ele[7][9];
    ele[5][8] != ele[8][8];
    ele[5][8] != ele[9][8];
    ele[5][9] != ele[10][9];
    ele[5][9] != ele[11][9];
    ele[5][9] != ele[12][9];
    ele[5][9] != ele[13][9];
    ele[5][9] != ele[14][9];
    ele[5][9] != ele[15][9];
    ele[5][9] != ele[5][10];
    ele[5][9] != ele[5][11];
    ele[5][9] != ele[5][12];
    ele[5][9] != ele[5][13];
    ele[5][9] != ele[5][14];
    ele[5][9] != ele[5][15];
    ele[5][9] != ele[6][10];
    ele[5][9] != ele[6][11];
    ele[5][9] != ele[6][8];
    ele[5][9] != ele[6][9];
    ele[5][9] != ele[7][10];
    ele[5][9] != ele[7][11];
    ele[5][9] != ele[7][8];
    ele[5][9] != ele[7][9];
    ele[5][9] != ele[8][9];
    ele[5][9] != ele[9][9];
    ele[6][0] != ele[10][0];
    ele[6][0] != ele[11][0];
    ele[6][0] != ele[12][0];
    ele[6][0] != ele[13][0];
    ele[6][0] != ele[14][0];
    ele[6][0] != ele[15][0];
    ele[6][0] != ele[6][1];
    ele[6][0] != ele[6][10];
    ele[6][0] != ele[6][11];
    ele[6][0] != ele[6][12];
    ele[6][0] != ele[6][13];
    ele[6][0] != ele[6][14];
    ele[6][0] != ele[6][15];
    ele[6][0] != ele[6][2];
    ele[6][0] != ele[6][3];
    ele[6][0] != ele[6][4];
    ele[6][0] != ele[6][5];
    ele[6][0] != ele[6][6];
    ele[6][0] != ele[6][7];
    ele[6][0] != ele[6][8];
    ele[6][0] != ele[6][9];
    ele[6][0] != ele[7][0];
    ele[6][0] != ele[7][1];
    ele[6][0] != ele[7][2];
    ele[6][0] != ele[7][3];
    ele[6][0] != ele[8][0];
    ele[6][0] != ele[9][0];
    ele[6][1] != ele[10][1];
    ele[6][1] != ele[11][1];
    ele[6][1] != ele[12][1];
    ele[6][1] != ele[13][1];
    ele[6][1] != ele[14][1];
    ele[6][1] != ele[15][1];
    ele[6][1] != ele[6][10];
    ele[6][1] != ele[6][11];
    ele[6][1] != ele[6][12];
    ele[6][1] != ele[6][13];
    ele[6][1] != ele[6][14];
    ele[6][1] != ele[6][15];
    ele[6][1] != ele[6][2];
    ele[6][1] != ele[6][3];
    ele[6][1] != ele[6][4];
    ele[6][1] != ele[6][5];
    ele[6][1] != ele[6][6];
    ele[6][1] != ele[6][7];
    ele[6][1] != ele[6][8];
    ele[6][1] != ele[6][9];
    ele[6][1] != ele[7][0];
    ele[6][1] != ele[7][1];
    ele[6][1] != ele[7][2];
    ele[6][1] != ele[7][3];
    ele[6][1] != ele[8][1];
    ele[6][1] != ele[9][1];
    ele[6][10] != ele[10][10];
    ele[6][10] != ele[11][10];
    ele[6][10] != ele[12][10];
    ele[6][10] != ele[13][10];
    ele[6][10] != ele[14][10];
    ele[6][10] != ele[15][10];
    ele[6][10] != ele[6][11];
    ele[6][10] != ele[6][12];
    ele[6][10] != ele[6][13];
    ele[6][10] != ele[6][14];
    ele[6][10] != ele[6][15];
    ele[6][10] != ele[7][10];
    ele[6][10] != ele[7][11];
    ele[6][10] != ele[7][8];
    ele[6][10] != ele[7][9];
    ele[6][10] != ele[8][10];
    ele[6][10] != ele[9][10];
    ele[6][11] != ele[10][11];
    ele[6][11] != ele[11][11];
    ele[6][11] != ele[12][11];
    ele[6][11] != ele[13][11];
    ele[6][11] != ele[14][11];
    ele[6][11] != ele[15][11];
    ele[6][11] != ele[6][12];
    ele[6][11] != ele[6][13];
    ele[6][11] != ele[6][14];
    ele[6][11] != ele[6][15];
    ele[6][11] != ele[7][10];
    ele[6][11] != ele[7][11];
    ele[6][11] != ele[7][8];
    ele[6][11] != ele[7][9];
    ele[6][11] != ele[8][11];
    ele[6][11] != ele[9][11];
    ele[6][12] != ele[10][12];
    ele[6][12] != ele[11][12];
    ele[6][12] != ele[12][12];
    ele[6][12] != ele[13][12];
    ele[6][12] != ele[14][12];
    ele[6][12] != ele[15][12];
    ele[6][12] != ele[6][13];
    ele[6][12] != ele[6][14];
    ele[6][12] != ele[6][15];
    ele[6][12] != ele[7][12];
    ele[6][12] != ele[7][13];
    ele[6][12] != ele[7][14];
    ele[6][12] != ele[7][15];
    ele[6][12] != ele[8][12];
    ele[6][12] != ele[9][12];
    ele[6][13] != ele[10][13];
    ele[6][13] != ele[11][13];
    ele[6][13] != ele[12][13];
    ele[6][13] != ele[13][13];
    ele[6][13] != ele[14][13];
    ele[6][13] != ele[15][13];
    ele[6][13] != ele[6][14];
    ele[6][13] != ele[6][15];
    ele[6][13] != ele[7][12];
    ele[6][13] != ele[7][13];
    ele[6][13] != ele[7][14];
    ele[6][13] != ele[7][15];
    ele[6][13] != ele[8][13];
    ele[6][13] != ele[9][13];
    ele[6][14] != ele[10][14];
    ele[6][14] != ele[11][14];
    ele[6][14] != ele[12][14];
    ele[6][14] != ele[13][14];
    ele[6][14] != ele[14][14];
    ele[6][14] != ele[15][14];
    ele[6][14] != ele[6][15];
    ele[6][14] != ele[7][12];
    ele[6][14] != ele[7][13];
    ele[6][14] != ele[7][14];
    ele[6][14] != ele[7][15];
    ele[6][14] != ele[8][14];
    ele[6][14] != ele[9][14];
    ele[6][15] != ele[10][15];
    ele[6][15] != ele[11][15];
    ele[6][15] != ele[12][15];
    ele[6][15] != ele[13][15];
    ele[6][15] != ele[14][15];
    ele[6][15] != ele[15][15];
    ele[6][15] != ele[7][12];
    ele[6][15] != ele[7][13];
    ele[6][15] != ele[7][14];
    ele[6][15] != ele[7][15];
    ele[6][15] != ele[8][15];
    ele[6][15] != ele[9][15];
    ele[6][2] != ele[10][2];
    ele[6][2] != ele[11][2];
    ele[6][2] != ele[12][2];
    ele[6][2] != ele[13][2];
    ele[6][2] != ele[14][2];
    ele[6][2] != ele[15][2];
    ele[6][2] != ele[6][10];
    ele[6][2] != ele[6][11];
    ele[6][2] != ele[6][12];
    ele[6][2] != ele[6][13];
    ele[6][2] != ele[6][14];
    ele[6][2] != ele[6][15];
    ele[6][2] != ele[6][3];
    ele[6][2] != ele[6][4];
    ele[6][2] != ele[6][5];
    ele[6][2] != ele[6][6];
    ele[6][2] != ele[6][7];
    ele[6][2] != ele[6][8];
    ele[6][2] != ele[6][9];
    ele[6][2] != ele[7][0];
    ele[6][2] != ele[7][1];
    ele[6][2] != ele[7][2];
    ele[6][2] != ele[7][3];
    ele[6][2] != ele[8][2];
    ele[6][2] != ele[9][2];
    ele[6][3] != ele[10][3];
    ele[6][3] != ele[11][3];
    ele[6][3] != ele[12][3];
    ele[6][3] != ele[13][3];
    ele[6][3] != ele[14][3];
    ele[6][3] != ele[15][3];
    ele[6][3] != ele[6][10];
    ele[6][3] != ele[6][11];
    ele[6][3] != ele[6][12];
    ele[6][3] != ele[6][13];
    ele[6][3] != ele[6][14];
    ele[6][3] != ele[6][15];
    ele[6][3] != ele[6][4];
    ele[6][3] != ele[6][5];
    ele[6][3] != ele[6][6];
    ele[6][3] != ele[6][7];
    ele[6][3] != ele[6][8];
    ele[6][3] != ele[6][9];
    ele[6][3] != ele[7][0];
    ele[6][3] != ele[7][1];
    ele[6][3] != ele[7][2];
    ele[6][3] != ele[7][3];
    ele[6][3] != ele[8][3];
    ele[6][3] != ele[9][3];
    ele[6][4] != ele[10][4];
    ele[6][4] != ele[11][4];
    ele[6][4] != ele[12][4];
    ele[6][4] != ele[13][4];
    ele[6][4] != ele[14][4];
    ele[6][4] != ele[15][4];
    ele[6][4] != ele[6][10];
    ele[6][4] != ele[6][11];
    ele[6][4] != ele[6][12];
    ele[6][4] != ele[6][13];
    ele[6][4] != ele[6][14];
    ele[6][4] != ele[6][15];
    ele[6][4] != ele[6][5];
    ele[6][4] != ele[6][6];
    ele[6][4] != ele[6][7];
    ele[6][4] != ele[6][8];
    ele[6][4] != ele[6][9];
    ele[6][4] != ele[7][4];
    ele[6][4] != ele[7][5];
    ele[6][4] != ele[7][6];
    ele[6][4] != ele[7][7];
    ele[6][4] != ele[8][4];
    ele[6][4] != ele[9][4];
    ele[6][5] != ele[10][5];
    ele[6][5] != ele[11][5];
    ele[6][5] != ele[12][5];
    ele[6][5] != ele[13][5];
    ele[6][5] != ele[14][5];
    ele[6][5] != ele[15][5];
    ele[6][5] != ele[6][10];
    ele[6][5] != ele[6][11];
    ele[6][5] != ele[6][12];
    ele[6][5] != ele[6][13];
    ele[6][5] != ele[6][14];
    ele[6][5] != ele[6][15];
    ele[6][5] != ele[6][6];
    ele[6][5] != ele[6][7];
    ele[6][5] != ele[6][8];
    ele[6][5] != ele[6][9];
    ele[6][5] != ele[7][4];
    ele[6][5] != ele[7][5];
    ele[6][5] != ele[7][6];
    ele[6][5] != ele[7][7];
    ele[6][5] != ele[8][5];
    ele[6][5] != ele[9][5];
    ele[6][6] != ele[10][6];
    ele[6][6] != ele[11][6];
    ele[6][6] != ele[12][6];
    ele[6][6] != ele[13][6];
    ele[6][6] != ele[14][6];
    ele[6][6] != ele[15][6];
    ele[6][6] != ele[6][10];
    ele[6][6] != ele[6][11];
    ele[6][6] != ele[6][12];
    ele[6][6] != ele[6][13];
    ele[6][6] != ele[6][14];
    ele[6][6] != ele[6][15];
    ele[6][6] != ele[6][7];
    ele[6][6] != ele[6][8];
    ele[6][6] != ele[6][9];
    ele[6][6] != ele[7][4];
    ele[6][6] != ele[7][5];
    ele[6][6] != ele[7][6];
    ele[6][6] != ele[7][7];
    ele[6][6] != ele[8][6];
    ele[6][6] != ele[9][6];
    ele[6][7] != ele[10][7];
    ele[6][7] != ele[11][7];
    ele[6][7] != ele[12][7];
    ele[6][7] != ele[13][7];
    ele[6][7] != ele[14][7];
    ele[6][7] != ele[15][7];
    ele[6][7] != ele[6][10];
    ele[6][7] != ele[6][11];
    ele[6][7] != ele[6][12];
    ele[6][7] != ele[6][13];
    ele[6][7] != ele[6][14];
    ele[6][7] != ele[6][15];
    ele[6][7] != ele[6][8];
    ele[6][7] != ele[6][9];
    ele[6][7] != ele[7][4];
    ele[6][7] != ele[7][5];
    ele[6][7] != ele[7][6];
    ele[6][7] != ele[7][7];
    ele[6][7] != ele[8][7];
    ele[6][7] != ele[9][7];
    ele[6][8] != ele[10][8];
    ele[6][8] != ele[11][8];
    ele[6][8] != ele[12][8];
    ele[6][8] != ele[13][8];
    ele[6][8] != ele[14][8];
    ele[6][8] != ele[15][8];
    ele[6][8] != ele[6][10];
    ele[6][8] != ele[6][11];
    ele[6][8] != ele[6][12];
    ele[6][8] != ele[6][13];
    ele[6][8] != ele[6][14];
    ele[6][8] != ele[6][15];
    ele[6][8] != ele[6][9];
    ele[6][8] != ele[7][10];
    ele[6][8] != ele[7][11];
    ele[6][8] != ele[7][8];
    ele[6][8] != ele[7][9];
    ele[6][8] != ele[8][8];
    ele[6][8] != ele[9][8];
    ele[6][9] != ele[10][9];
    ele[6][9] != ele[11][9];
    ele[6][9] != ele[12][9];
    ele[6][9] != ele[13][9];
    ele[6][9] != ele[14][9];
    ele[6][9] != ele[15][9];
    ele[6][9] != ele[6][10];
    ele[6][9] != ele[6][11];
    ele[6][9] != ele[6][12];
    ele[6][9] != ele[6][13];
    ele[6][9] != ele[6][14];
    ele[6][9] != ele[6][15];
    ele[6][9] != ele[7][10];
    ele[6][9] != ele[7][11];
    ele[6][9] != ele[7][8];
    ele[6][9] != ele[7][9];
    ele[6][9] != ele[8][9];
    ele[6][9] != ele[9][9];
    ele[7][0] != ele[10][0];
    ele[7][0] != ele[11][0];
    ele[7][0] != ele[12][0];
    ele[7][0] != ele[13][0];
    ele[7][0] != ele[14][0];
    ele[7][0] != ele[15][0];
    ele[7][0] != ele[7][1];
    ele[7][0] != ele[7][10];
    ele[7][0] != ele[7][11];
    ele[7][0] != ele[7][12];
    ele[7][0] != ele[7][13];
    ele[7][0] != ele[7][14];
    ele[7][0] != ele[7][15];
    ele[7][0] != ele[7][2];
    ele[7][0] != ele[7][3];
    ele[7][0] != ele[7][4];
    ele[7][0] != ele[7][5];
    ele[7][0] != ele[7][6];
    ele[7][0] != ele[7][7];
    ele[7][0] != ele[7][8];
    ele[7][0] != ele[7][9];
    ele[7][0] != ele[8][0];
    ele[7][0] != ele[9][0];
    ele[7][1] != ele[10][1];
    ele[7][1] != ele[11][1];
    ele[7][1] != ele[12][1];
    ele[7][1] != ele[13][1];
    ele[7][1] != ele[14][1];
    ele[7][1] != ele[15][1];
    ele[7][1] != ele[7][10];
    ele[7][1] != ele[7][11];
    ele[7][1] != ele[7][12];
    ele[7][1] != ele[7][13];
    ele[7][1] != ele[7][14];
    ele[7][1] != ele[7][15];
    ele[7][1] != ele[7][2];
    ele[7][1] != ele[7][3];
    ele[7][1] != ele[7][4];
    ele[7][1] != ele[7][5];
    ele[7][1] != ele[7][6];
    ele[7][1] != ele[7][7];
    ele[7][1] != ele[7][8];
    ele[7][1] != ele[7][9];
    ele[7][1] != ele[8][1];
    ele[7][1] != ele[9][1];
    ele[7][10] != ele[10][10];
    ele[7][10] != ele[11][10];
    ele[7][10] != ele[12][10];
    ele[7][10] != ele[13][10];
    ele[7][10] != ele[14][10];
    ele[7][10] != ele[15][10];
    ele[7][10] != ele[7][11];
    ele[7][10] != ele[7][12];
    ele[7][10] != ele[7][13];
    ele[7][10] != ele[7][14];
    ele[7][10] != ele[7][15];
    ele[7][10] != ele[8][10];
    ele[7][10] != ele[9][10];
    ele[7][11] != ele[10][11];
    ele[7][11] != ele[11][11];
    ele[7][11] != ele[12][11];
    ele[7][11] != ele[13][11];
    ele[7][11] != ele[14][11];
    ele[7][11] != ele[15][11];
    ele[7][11] != ele[7][12];
    ele[7][11] != ele[7][13];
    ele[7][11] != ele[7][14];
    ele[7][11] != ele[7][15];
    ele[7][11] != ele[8][11];
    ele[7][11] != ele[9][11];
    ele[7][12] != ele[10][12];
    ele[7][12] != ele[11][12];
    ele[7][12] != ele[12][12];
    ele[7][12] != ele[13][12];
    ele[7][12] != ele[14][12];
    ele[7][12] != ele[15][12];
    ele[7][12] != ele[7][13];
    ele[7][12] != ele[7][14];
    ele[7][12] != ele[7][15];
    ele[7][12] != ele[8][12];
    ele[7][12] != ele[9][12];
    ele[7][13] != ele[10][13];
    ele[7][13] != ele[11][13];
    ele[7][13] != ele[12][13];
    ele[7][13] != ele[13][13];
    ele[7][13] != ele[14][13];
    ele[7][13] != ele[15][13];
    ele[7][13] != ele[7][14];
    ele[7][13] != ele[7][15];
    ele[7][13] != ele[8][13];
    ele[7][13] != ele[9][13];
    ele[7][14] != ele[10][14];
    ele[7][14] != ele[11][14];
    ele[7][14] != ele[12][14];
    ele[7][14] != ele[13][14];
    ele[7][14] != ele[14][14];
    ele[7][14] != ele[15][14];
    ele[7][14] != ele[7][15];
    ele[7][14] != ele[8][14];
    ele[7][14] != ele[9][14];
    ele[7][15] != ele[10][15];
    ele[7][15] != ele[11][15];
    ele[7][15] != ele[12][15];
    ele[7][15] != ele[13][15];
    ele[7][15] != ele[14][15];
    ele[7][15] != ele[15][15];
    ele[7][15] != ele[8][15];
    ele[7][15] != ele[9][15];
    ele[7][2] != ele[10][2];
    ele[7][2] != ele[11][2];
    ele[7][2] != ele[12][2];
    ele[7][2] != ele[13][2];
    ele[7][2] != ele[14][2];
    ele[7][2] != ele[15][2];
    ele[7][2] != ele[7][10];
    ele[7][2] != ele[7][11];
    ele[7][2] != ele[7][12];
    ele[7][2] != ele[7][13];
    ele[7][2] != ele[7][14];
    ele[7][2] != ele[7][15];
    ele[7][2] != ele[7][3];
    ele[7][2] != ele[7][4];
    ele[7][2] != ele[7][5];
    ele[7][2] != ele[7][6];
    ele[7][2] != ele[7][7];
    ele[7][2] != ele[7][8];
    ele[7][2] != ele[7][9];
    ele[7][2] != ele[8][2];
    ele[7][2] != ele[9][2];
    ele[7][3] != ele[10][3];
    ele[7][3] != ele[11][3];
    ele[7][3] != ele[12][3];
    ele[7][3] != ele[13][3];
    ele[7][3] != ele[14][3];
    ele[7][3] != ele[15][3];
    ele[7][3] != ele[7][10];
    ele[7][3] != ele[7][11];
    ele[7][3] != ele[7][12];
    ele[7][3] != ele[7][13];
    ele[7][3] != ele[7][14];
    ele[7][3] != ele[7][15];
    ele[7][3] != ele[7][4];
    ele[7][3] != ele[7][5];
    ele[7][3] != ele[7][6];
    ele[7][3] != ele[7][7];
    ele[7][3] != ele[7][8];
    ele[7][3] != ele[7][9];
    ele[7][3] != ele[8][3];
    ele[7][3] != ele[9][3];
    ele[7][4] != ele[10][4];
    ele[7][4] != ele[11][4];
    ele[7][4] != ele[12][4];
    ele[7][4] != ele[13][4];
    ele[7][4] != ele[14][4];
    ele[7][4] != ele[15][4];
    ele[7][4] != ele[7][10];
    ele[7][4] != ele[7][11];
    ele[7][4] != ele[7][12];
    ele[7][4] != ele[7][13];
    ele[7][4] != ele[7][14];
    ele[7][4] != ele[7][15];
    ele[7][4] != ele[7][5];
    ele[7][4] != ele[7][6];
    ele[7][4] != ele[7][7];
    ele[7][4] != ele[7][8];
    ele[7][4] != ele[7][9];
    ele[7][4] != ele[8][4];
    ele[7][4] != ele[9][4];
    ele[7][5] != ele[10][5];
    ele[7][5] != ele[11][5];
    ele[7][5] != ele[12][5];
    ele[7][5] != ele[13][5];
    ele[7][5] != ele[14][5];
    ele[7][5] != ele[15][5];
    ele[7][5] != ele[7][10];
    ele[7][5] != ele[7][11];
    ele[7][5] != ele[7][12];
    ele[7][5] != ele[7][13];
    ele[7][5] != ele[7][14];
    ele[7][5] != ele[7][15];
    ele[7][5] != ele[7][6];
    ele[7][5] != ele[7][7];
    ele[7][5] != ele[7][8];
    ele[7][5] != ele[7][9];
    ele[7][5] != ele[8][5];
    ele[7][5] != ele[9][5];
    ele[7][6] != ele[10][6];
    ele[7][6] != ele[11][6];
    ele[7][6] != ele[12][6];
    ele[7][6] != ele[13][6];
    ele[7][6] != ele[14][6];
    ele[7][6] != ele[15][6];
    ele[7][6] != ele[7][10];
    ele[7][6] != ele[7][11];
    ele[7][6] != ele[7][12];
    ele[7][6] != ele[7][13];
    ele[7][6] != ele[7][14];
    ele[7][6] != ele[7][15];
    ele[7][6] != ele[7][7];
    ele[7][6] != ele[7][8];
    ele[7][6] != ele[7][9];
    ele[7][6] != ele[8][6];
    ele[7][6] != ele[9][6];
    ele[7][7] != ele[10][7];
    ele[7][7] != ele[11][7];
    ele[7][7] != ele[12][7];
    ele[7][7] != ele[13][7];
    ele[7][7] != ele[14][7];
    ele[7][7] != ele[15][7];
    ele[7][7] != ele[7][10];
    ele[7][7] != ele[7][11];
    ele[7][7] != ele[7][12];
    ele[7][7] != ele[7][13];
    ele[7][7] != ele[7][14];
    ele[7][7] != ele[7][15];
    ele[7][7] != ele[7][8];
    ele[7][7] != ele[7][9];
    ele[7][7] != ele[8][7];
    ele[7][7] != ele[9][7];
    ele[7][8] != ele[10][8];
    ele[7][8] != ele[11][8];
    ele[7][8] != ele[12][8];
    ele[7][8] != ele[13][8];
    ele[7][8] != ele[14][8];
    ele[7][8] != ele[15][8];
    ele[7][8] != ele[7][10];
    ele[7][8] != ele[7][11];
    ele[7][8] != ele[7][12];
    ele[7][8] != ele[7][13];
    ele[7][8] != ele[7][14];
    ele[7][8] != ele[7][15];
    ele[7][8] != ele[7][9];
    ele[7][8] != ele[8][8];
    ele[7][8] != ele[9][8];
    ele[7][9] != ele[10][9];
    ele[7][9] != ele[11][9];
    ele[7][9] != ele[12][9];
    ele[7][9] != ele[13][9];
    ele[7][9] != ele[14][9];
    ele[7][9] != ele[15][9];
    ele[7][9] != ele[7][10];
    ele[7][9] != ele[7][11];
    ele[7][9] != ele[7][12];
    ele[7][9] != ele[7][13];
    ele[7][9] != ele[7][14];
    ele[7][9] != ele[7][15];
    ele[7][9] != ele[8][9];
    ele[7][9] != ele[9][9];
    ele[8][0] != ele[10][0];
    ele[8][0] != ele[10][1];
    ele[8][0] != ele[10][2];
    ele[8][0] != ele[10][3];
    ele[8][0] != ele[11][0];
    ele[8][0] != ele[11][1];
    ele[8][0] != ele[11][2];
    ele[8][0] != ele[11][3];
    ele[8][0] != ele[12][0];
    ele[8][0] != ele[13][0];
    ele[8][0] != ele[14][0];
    ele[8][0] != ele[15][0];
    ele[8][0] != ele[8][1];
    ele[8][0] != ele[8][10];
    ele[8][0] != ele[8][11];
    ele[8][0] != ele[8][12];
    ele[8][0] != ele[8][13];
    ele[8][0] != ele[8][14];
    ele[8][0] != ele[8][15];
    ele[8][0] != ele[8][2];
    ele[8][0] != ele[8][3];
    ele[8][0] != ele[8][4];
    ele[8][0] != ele[8][5];
    ele[8][0] != ele[8][6];
    ele[8][0] != ele[8][7];
    ele[8][0] != ele[8][8];
    ele[8][0] != ele[8][9];
    ele[8][0] != ele[9][0];
    ele[8][0] != ele[9][1];
    ele[8][0] != ele[9][2];
    ele[8][0] != ele[9][3];
    ele[8][1] != ele[10][0];
    ele[8][1] != ele[10][1];
    ele[8][1] != ele[10][2];
    ele[8][1] != ele[10][3];
    ele[8][1] != ele[11][0];
    ele[8][1] != ele[11][1];
    ele[8][1] != ele[11][2];
    ele[8][1] != ele[11][3];
    ele[8][1] != ele[12][1];
    ele[8][1] != ele[13][1];
    ele[8][1] != ele[14][1];
    ele[8][1] != ele[15][1];
    ele[8][1] != ele[8][10];
    ele[8][1] != ele[8][11];
    ele[8][1] != ele[8][12];
    ele[8][1] != ele[8][13];
    ele[8][1] != ele[8][14];
    ele[8][1] != ele[8][15];
    ele[8][1] != ele[8][2];
    ele[8][1] != ele[8][3];
    ele[8][1] != ele[8][4];
    ele[8][1] != ele[8][5];
    ele[8][1] != ele[8][6];
    ele[8][1] != ele[8][7];
    ele[8][1] != ele[8][8];
    ele[8][1] != ele[8][9];
    ele[8][1] != ele[9][0];
    ele[8][1] != ele[9][1];
    ele[8][1] != ele[9][2];
    ele[8][1] != ele[9][3];
    ele[8][10] != ele[10][10];
    ele[8][10] != ele[10][11];
    ele[8][10] != ele[10][8];
    ele[8][10] != ele[10][9];
    ele[8][10] != ele[11][10];
    ele[8][10] != ele[11][11];
    ele[8][10] != ele[11][8];
    ele[8][10] != ele[11][9];
    ele[8][10] != ele[12][10];
    ele[8][10] != ele[13][10];
    ele[8][10] != ele[14][10];
    ele[8][10] != ele[15][10];
    ele[8][10] != ele[8][11];
    ele[8][10] != ele[8][12];
    ele[8][10] != ele[8][13];
    ele[8][10] != ele[8][14];
    ele[8][10] != ele[8][15];
    ele[8][10] != ele[9][10];
    ele[8][10] != ele[9][11];
    ele[8][10] != ele[9][8];
    ele[8][10] != ele[9][9];
    ele[8][11] != ele[10][10];
    ele[8][11] != ele[10][11];
    ele[8][11] != ele[10][8];
    ele[8][11] != ele[10][9];
    ele[8][11] != ele[11][10];
    ele[8][11] != ele[11][11];
    ele[8][11] != ele[11][8];
    ele[8][11] != ele[11][9];
    ele[8][11] != ele[12][11];
    ele[8][11] != ele[13][11];
    ele[8][11] != ele[14][11];
    ele[8][11] != ele[15][11];
    ele[8][11] != ele[8][12];
    ele[8][11] != ele[8][13];
    ele[8][11] != ele[8][14];
    ele[8][11] != ele[8][15];
    ele[8][11] != ele[9][10];
    ele[8][11] != ele[9][11];
    ele[8][11] != ele[9][8];
    ele[8][11] != ele[9][9];
    ele[8][12] != ele[10][12];
    ele[8][12] != ele[10][13];
    ele[8][12] != ele[10][14];
    ele[8][12] != ele[10][15];
    ele[8][12] != ele[11][12];
    ele[8][12] != ele[11][13];
    ele[8][12] != ele[11][14];
    ele[8][12] != ele[11][15];
    ele[8][12] != ele[12][12];
    ele[8][12] != ele[13][12];
    ele[8][12] != ele[14][12];
    ele[8][12] != ele[15][12];
    ele[8][12] != ele[8][13];
    ele[8][12] != ele[8][14];
    ele[8][12] != ele[8][15];
    ele[8][12] != ele[9][12];
    ele[8][12] != ele[9][13];
    ele[8][12] != ele[9][14];
    ele[8][12] != ele[9][15];
    ele[8][13] != ele[10][12];
    ele[8][13] != ele[10][13];
    ele[8][13] != ele[10][14];
    ele[8][13] != ele[10][15];
    ele[8][13] != ele[11][12];
    ele[8][13] != ele[11][13];
    ele[8][13] != ele[11][14];
    ele[8][13] != ele[11][15];
    ele[8][13] != ele[12][13];
    ele[8][13] != ele[13][13];
    ele[8][13] != ele[14][13];
    ele[8][13] != ele[15][13];
    ele[8][13] != ele[8][14];
    ele[8][13] != ele[8][15];
    ele[8][13] != ele[9][12];
    ele[8][13] != ele[9][13];
    ele[8][13] != ele[9][14];
    ele[8][13] != ele[9][15];
    ele[8][14] != ele[10][12];
    ele[8][14] != ele[10][13];
    ele[8][14] != ele[10][14];
    ele[8][14] != ele[10][15];
    ele[8][14] != ele[11][12];
    ele[8][14] != ele[11][13];
    ele[8][14] != ele[11][14];
    ele[8][14] != ele[11][15];
    ele[8][14] != ele[12][14];
    ele[8][14] != ele[13][14];
    ele[8][14] != ele[14][14];
    ele[8][14] != ele[15][14];
    ele[8][14] != ele[8][15];
    ele[8][14] != ele[9][12];
    ele[8][14] != ele[9][13];
    ele[8][14] != ele[9][14];
    ele[8][14] != ele[9][15];
    ele[8][15] != ele[10][12];
    ele[8][15] != ele[10][13];
    ele[8][15] != ele[10][14];
    ele[8][15] != ele[10][15];
    ele[8][15] != ele[11][12];
    ele[8][15] != ele[11][13];
    ele[8][15] != ele[11][14];
    ele[8][15] != ele[11][15];
    ele[8][15] != ele[12][15];
    ele[8][15] != ele[13][15];
    ele[8][15] != ele[14][15];
    ele[8][15] != ele[15][15];
    ele[8][15] != ele[9][12];
    ele[8][15] != ele[9][13];
    ele[8][15] != ele[9][14];
    ele[8][15] != ele[9][15];
    ele[8][2] != ele[10][0];
    ele[8][2] != ele[10][1];
    ele[8][2] != ele[10][2];
    ele[8][2] != ele[10][3];
    ele[8][2] != ele[11][0];
    ele[8][2] != ele[11][1];
    ele[8][2] != ele[11][2];
    ele[8][2] != ele[11][3];
    ele[8][2] != ele[12][2];
    ele[8][2] != ele[13][2];
    ele[8][2] != ele[14][2];
    ele[8][2] != ele[15][2];
    ele[8][2] != ele[8][10];
    ele[8][2] != ele[8][11];
    ele[8][2] != ele[8][12];
    ele[8][2] != ele[8][13];
    ele[8][2] != ele[8][14];
    ele[8][2] != ele[8][15];
    ele[8][2] != ele[8][3];
    ele[8][2] != ele[8][4];
    ele[8][2] != ele[8][5];
    ele[8][2] != ele[8][6];
    ele[8][2] != ele[8][7];
    ele[8][2] != ele[8][8];
    ele[8][2] != ele[8][9];
    ele[8][2] != ele[9][0];
    ele[8][2] != ele[9][1];
    ele[8][2] != ele[9][2];
    ele[8][2] != ele[9][3];
    ele[8][3] != ele[10][0];
    ele[8][3] != ele[10][1];
    ele[8][3] != ele[10][2];
    ele[8][3] != ele[10][3];
    ele[8][3] != ele[11][0];
    ele[8][3] != ele[11][1];
    ele[8][3] != ele[11][2];
    ele[8][3] != ele[11][3];
    ele[8][3] != ele[12][3];
    ele[8][3] != ele[13][3];
    ele[8][3] != ele[14][3];
    ele[8][3] != ele[15][3];
    ele[8][3] != ele[8][10];
    ele[8][3] != ele[8][11];
    ele[8][3] != ele[8][12];
    ele[8][3] != ele[8][13];
    ele[8][3] != ele[8][14];
    ele[8][3] != ele[8][15];
    ele[8][3] != ele[8][4];
    ele[8][3] != ele[8][5];
    ele[8][3] != ele[8][6];
    ele[8][3] != ele[8][7];
    ele[8][3] != ele[8][8];
    ele[8][3] != ele[8][9];
    ele[8][3] != ele[9][0];
    ele[8][3] != ele[9][1];
    ele[8][3] != ele[9][2];
    ele[8][3] != ele[9][3];
    ele[8][4] != ele[10][4];
    ele[8][4] != ele[10][5];
    ele[8][4] != ele[10][6];
    ele[8][4] != ele[10][7];
    ele[8][4] != ele[11][4];
    ele[8][4] != ele[11][5];
    ele[8][4] != ele[11][6];
    ele[8][4] != ele[11][7];
    ele[8][4] != ele[12][4];
    ele[8][4] != ele[13][4];
    ele[8][4] != ele[14][4];
    ele[8][4] != ele[15][4];
    ele[8][4] != ele[8][10];
    ele[8][4] != ele[8][11];
    ele[8][4] != ele[8][12];
    ele[8][4] != ele[8][13];
    ele[8][4] != ele[8][14];
    ele[8][4] != ele[8][15];
    ele[8][4] != ele[8][5];
    ele[8][4] != ele[8][6];
    ele[8][4] != ele[8][7];
    ele[8][4] != ele[8][8];
    ele[8][4] != ele[8][9];
    ele[8][4] != ele[9][4];
    ele[8][4] != ele[9][5];
    ele[8][4] != ele[9][6];
    ele[8][4] != ele[9][7];
    ele[8][5] != ele[10][4];
    ele[8][5] != ele[10][5];
    ele[8][5] != ele[10][6];
    ele[8][5] != ele[10][7];
    ele[8][5] != ele[11][4];
    ele[8][5] != ele[11][5];
    ele[8][5] != ele[11][6];
    ele[8][5] != ele[11][7];
    ele[8][5] != ele[12][5];
    ele[8][5] != ele[13][5];
    ele[8][5] != ele[14][5];
    ele[8][5] != ele[15][5];
    ele[8][5] != ele[8][10];
    ele[8][5] != ele[8][11];
    ele[8][5] != ele[8][12];
    ele[8][5] != ele[8][13];
    ele[8][5] != ele[8][14];
    ele[8][5] != ele[8][15];
    ele[8][5] != ele[8][6];
    ele[8][5] != ele[8][7];
    ele[8][5] != ele[8][8];
    ele[8][5] != ele[8][9];
    ele[8][5] != ele[9][4];
    ele[8][5] != ele[9][5];
    ele[8][5] != ele[9][6];
    ele[8][5] != ele[9][7];
    ele[8][6] != ele[10][4];
    ele[8][6] != ele[10][5];
    ele[8][6] != ele[10][6];
    ele[8][6] != ele[10][7];
    ele[8][6] != ele[11][4];
    ele[8][6] != ele[11][5];
    ele[8][6] != ele[11][6];
    ele[8][6] != ele[11][7];
    ele[8][6] != ele[12][6];
    ele[8][6] != ele[13][6];
    ele[8][6] != ele[14][6];
    ele[8][6] != ele[15][6];
    ele[8][6] != ele[8][10];
    ele[8][6] != ele[8][11];
    ele[8][6] != ele[8][12];
    ele[8][6] != ele[8][13];
    ele[8][6] != ele[8][14];
    ele[8][6] != ele[8][15];
    ele[8][6] != ele[8][7];
    ele[8][6] != ele[8][8];
    ele[8][6] != ele[8][9];
    ele[8][6] != ele[9][4];
    ele[8][6] != ele[9][5];
    ele[8][6] != ele[9][6];
    ele[8][6] != ele[9][7];
    ele[8][7] != ele[10][4];
    ele[8][7] != ele[10][5];
    ele[8][7] != ele[10][6];
    ele[8][7] != ele[10][7];
    ele[8][7] != ele[11][4];
    ele[8][7] != ele[11][5];
    ele[8][7] != ele[11][6];
    ele[8][7] != ele[11][7];
    ele[8][7] != ele[12][7];
    ele[8][7] != ele[13][7];
    ele[8][7] != ele[14][7];
    ele[8][7] != ele[15][7];
    ele[8][7] != ele[8][10];
    ele[8][7] != ele[8][11];
    ele[8][7] != ele[8][12];
    ele[8][7] != ele[8][13];
    ele[8][7] != ele[8][14];
    ele[8][7] != ele[8][15];
    ele[8][7] != ele[8][8];
    ele[8][7] != ele[8][9];
    ele[8][7] != ele[9][4];
    ele[8][7] != ele[9][5];
    ele[8][7] != ele[9][6];
    ele[8][7] != ele[9][7];
    ele[8][8] != ele[10][10];
    ele[8][8] != ele[10][11];
    ele[8][8] != ele[10][8];
    ele[8][8] != ele[10][9];
    ele[8][8] != ele[11][10];
    ele[8][8] != ele[11][11];
    ele[8][8] != ele[11][8];
    ele[8][8] != ele[11][9];
    ele[8][8] != ele[12][8];
    ele[8][8] != ele[13][8];
    ele[8][8] != ele[14][8];
    ele[8][8] != ele[15][8];
    ele[8][8] != ele[8][10];
    ele[8][8] != ele[8][11];
    ele[8][8] != ele[8][12];
    ele[8][8] != ele[8][13];
    ele[8][8] != ele[8][14];
    ele[8][8] != ele[8][15];
    ele[8][8] != ele[8][9];
    ele[8][8] != ele[9][10];
    ele[8][8] != ele[9][11];
    ele[8][8] != ele[9][8];
    ele[8][8] != ele[9][9];
    ele[8][9] != ele[10][10];
    ele[8][9] != ele[10][11];
    ele[8][9] != ele[10][8];
    ele[8][9] != ele[10][9];
    ele[8][9] != ele[11][10];
    ele[8][9] != ele[11][11];
    ele[8][9] != ele[11][8];
    ele[8][9] != ele[11][9];
    ele[8][9] != ele[12][9];
    ele[8][9] != ele[13][9];
    ele[8][9] != ele[14][9];
    ele[8][9] != ele[15][9];
    ele[8][9] != ele[8][10];
    ele[8][9] != ele[8][11];
    ele[8][9] != ele[8][12];
    ele[8][9] != ele[8][13];
    ele[8][9] != ele[8][14];
    ele[8][9] != ele[8][15];
    ele[8][9] != ele[9][10];
    ele[8][9] != ele[9][11];
    ele[8][9] != ele[9][8];
    ele[8][9] != ele[9][9];
    ele[9][0] != ele[10][0];
    ele[9][0] != ele[10][1];
    ele[9][0] != ele[10][2];
    ele[9][0] != ele[10][3];
    ele[9][0] != ele[11][0];
    ele[9][0] != ele[11][1];
    ele[9][0] != ele[11][2];
    ele[9][0] != ele[11][3];
    ele[9][0] != ele[12][0];
    ele[9][0] != ele[13][0];
    ele[9][0] != ele[14][0];
    ele[9][0] != ele[15][0];
    ele[9][0] != ele[9][1];
    ele[9][0] != ele[9][10];
    ele[9][0] != ele[9][11];
    ele[9][0] != ele[9][12];
    ele[9][0] != ele[9][13];
    ele[9][0] != ele[9][14];
    ele[9][0] != ele[9][15];
    ele[9][0] != ele[9][2];
    ele[9][0] != ele[9][3];
    ele[9][0] != ele[9][4];
    ele[9][0] != ele[9][5];
    ele[9][0] != ele[9][6];
    ele[9][0] != ele[9][7];
    ele[9][0] != ele[9][8];
    ele[9][0] != ele[9][9];
    ele[9][1] != ele[10][0];
    ele[9][1] != ele[10][1];
    ele[9][1] != ele[10][2];
    ele[9][1] != ele[10][3];
    ele[9][1] != ele[11][0];
    ele[9][1] != ele[11][1];
    ele[9][1] != ele[11][2];
    ele[9][1] != ele[11][3];
    ele[9][1] != ele[12][1];
    ele[9][1] != ele[13][1];
    ele[9][1] != ele[14][1];
    ele[9][1] != ele[15][1];
    ele[9][1] != ele[9][10];
    ele[9][1] != ele[9][11];
    ele[9][1] != ele[9][12];
    ele[9][1] != ele[9][13];
    ele[9][1] != ele[9][14];
    ele[9][1] != ele[9][15];
    ele[9][1] != ele[9][2];
    ele[9][1] != ele[9][3];
    ele[9][1] != ele[9][4];
    ele[9][1] != ele[9][5];
    ele[9][1] != ele[9][6];
    ele[9][1] != ele[9][7];
    ele[9][1] != ele[9][8];
    ele[9][1] != ele[9][9];
    ele[9][10] != ele[10][10];
    ele[9][10] != ele[10][11];
    ele[9][10] != ele[10][8];
    ele[9][10] != ele[10][9];
    ele[9][10] != ele[11][10];
    ele[9][10] != ele[11][11];
    ele[9][10] != ele[11][8];
    ele[9][10] != ele[11][9];
    ele[9][10] != ele[12][10];
    ele[9][10] != ele[13][10];
    ele[9][10] != ele[14][10];
    ele[9][10] != ele[15][10];
    ele[9][10] != ele[9][11];
    ele[9][10] != ele[9][12];
    ele[9][10] != ele[9][13];
    ele[9][10] != ele[9][14];
    ele[9][10] != ele[9][15];
    ele[9][11] != ele[10][10];
    ele[9][11] != ele[10][11];
    ele[9][11] != ele[10][8];
    ele[9][11] != ele[10][9];
    ele[9][11] != ele[11][10];
    ele[9][11] != ele[11][11];
    ele[9][11] != ele[11][8];
    ele[9][11] != ele[11][9];
    ele[9][11] != ele[12][11];
    ele[9][11] != ele[13][11];
    ele[9][11] != ele[14][11];
    ele[9][11] != ele[15][11];
    ele[9][11] != ele[9][12];
    ele[9][11] != ele[9][13];
    ele[9][11] != ele[9][14];
    ele[9][11] != ele[9][15];
    ele[9][12] != ele[10][12];
    ele[9][12] != ele[10][13];
    ele[9][12] != ele[10][14];
    ele[9][12] != ele[10][15];
    ele[9][12] != ele[11][12];
    ele[9][12] != ele[11][13];
    ele[9][12] != ele[11][14];
    ele[9][12] != ele[11][15];
    ele[9][12] != ele[12][12];
    ele[9][12] != ele[13][12];
    ele[9][12] != ele[14][12];
    ele[9][12] != ele[15][12];
    ele[9][12] != ele[9][13];
    ele[9][12] != ele[9][14];
    ele[9][12] != ele[9][15];
    ele[9][13] != ele[10][12];
    ele[9][13] != ele[10][13];
    ele[9][13] != ele[10][14];
    ele[9][13] != ele[10][15];
    ele[9][13] != ele[11][12];
    ele[9][13] != ele[11][13];
    ele[9][13] != ele[11][14];
    ele[9][13] != ele[11][15];
    ele[9][13] != ele[12][13];
    ele[9][13] != ele[13][13];
    ele[9][13] != ele[14][13];
    ele[9][13] != ele[15][13];
    ele[9][13] != ele[9][14];
    ele[9][13] != ele[9][15];
    ele[9][14] != ele[10][12];
    ele[9][14] != ele[10][13];
    ele[9][14] != ele[10][14];
    ele[9][14] != ele[10][15];
    ele[9][14] != ele[11][12];
    ele[9][14] != ele[11][13];
    ele[9][14] != ele[11][14];
    ele[9][14] != ele[11][15];
    ele[9][14] != ele[12][14];
    ele[9][14] != ele[13][14];
    ele[9][14] != ele[14][14];
    ele[9][14] != ele[15][14];
    ele[9][14] != ele[9][15];
    ele[9][15] != ele[10][12];
    ele[9][15] != ele[10][13];
    ele[9][15] != ele[10][14];
    ele[9][15] != ele[10][15];
    ele[9][15] != ele[11][12];
    ele[9][15] != ele[11][13];
    ele[9][15] != ele[11][14];
    ele[9][15] != ele[11][15];
    ele[9][15] != ele[12][15];
    ele[9][15] != ele[13][15];
    ele[9][15] != ele[14][15];
    ele[9][15] != ele[15][15];
    ele[9][2] != ele[10][0];
    ele[9][2] != ele[10][1];
    ele[9][2] != ele[10][2];
    ele[9][2] != ele[10][3];
    ele[9][2] != ele[11][0];
    ele[9][2] != ele[11][1];
    ele[9][2] != ele[11][2];
    ele[9][2] != ele[11][3];
    ele[9][2] != ele[12][2];
    ele[9][2] != ele[13][2];
    ele[9][2] != ele[14][2];
    ele[9][2] != ele[15][2];
    ele[9][2] != ele[9][10];
    ele[9][2] != ele[9][11];
    ele[9][2] != ele[9][12];
    ele[9][2] != ele[9][13];
    ele[9][2] != ele[9][14];
    ele[9][2] != ele[9][15];
    ele[9][2] != ele[9][3];
    ele[9][2] != ele[9][4];
    ele[9][2] != ele[9][5];
    ele[9][2] != ele[9][6];
    ele[9][2] != ele[9][7];
    ele[9][2] != ele[9][8];
    ele[9][2] != ele[9][9];
    ele[9][3] != ele[10][0];
    ele[9][3] != ele[10][1];
    ele[9][3] != ele[10][2];
    ele[9][3] != ele[10][3];
    ele[9][3] != ele[11][0];
    ele[9][3] != ele[11][1];
    ele[9][3] != ele[11][2];
    ele[9][3] != ele[11][3];
    ele[9][3] != ele[12][3];
    ele[9][3] != ele[13][3];
    ele[9][3] != ele[14][3];
    ele[9][3] != ele[15][3];
    ele[9][3] != ele[9][10];
    ele[9][3] != ele[9][11];
    ele[9][3] != ele[9][12];
    ele[9][3] != ele[9][13];
    ele[9][3] != ele[9][14];
    ele[9][3] != ele[9][15];
    ele[9][3] != ele[9][4];
    ele[9][3] != ele[9][5];
    ele[9][3] != ele[9][6];
    ele[9][3] != ele[9][7];
    ele[9][3] != ele[9][8];
    ele[9][3] != ele[9][9];
    ele[9][4] != ele[10][4];
    ele[9][4] != ele[10][5];
    ele[9][4] != ele[10][6];
    ele[9][4] != ele[10][7];
    ele[9][4] != ele[11][4];
    ele[9][4] != ele[11][5];
    ele[9][4] != ele[11][6];
    ele[9][4] != ele[11][7];
    ele[9][4] != ele[12][4];
    ele[9][4] != ele[13][4];
    ele[9][4] != ele[14][4];
    ele[9][4] != ele[15][4];
    ele[9][4] != ele[9][10];
    ele[9][4] != ele[9][11];
    ele[9][4] != ele[9][12];
    ele[9][4] != ele[9][13];
    ele[9][4] != ele[9][14];
    ele[9][4] != ele[9][15];
    ele[9][4] != ele[9][5];
    ele[9][4] != ele[9][6];
    ele[9][4] != ele[9][7];
    ele[9][4] != ele[9][8];
    ele[9][4] != ele[9][9];
    ele[9][5] != ele[10][4];
    ele[9][5] != ele[10][5];
    ele[9][5] != ele[10][6];
    ele[9][5] != ele[10][7];
    ele[9][5] != ele[11][4];
    ele[9][5] != ele[11][5];
    ele[9][5] != ele[11][6];
    ele[9][5] != ele[11][7];
    ele[9][5] != ele[12][5];
    ele[9][5] != ele[13][5];
    ele[9][5] != ele[14][5];
    ele[9][5] != ele[15][5];
    ele[9][5] != ele[9][10];
    ele[9][5] != ele[9][11];
    ele[9][5] != ele[9][12];
    ele[9][5] != ele[9][13];
    ele[9][5] != ele[9][14];
    ele[9][5] != ele[9][15];
    ele[9][5] != ele[9][6];
    ele[9][5] != ele[9][7];
    ele[9][5] != ele[9][8];
    ele[9][5] != ele[9][9];
    ele[9][6] != ele[10][4];
    ele[9][6] != ele[10][5];
    ele[9][6] != ele[10][6];
    ele[9][6] != ele[10][7];
    ele[9][6] != ele[11][4];
    ele[9][6] != ele[11][5];
    ele[9][6] != ele[11][6];
    ele[9][6] != ele[11][7];
    ele[9][6] != ele[12][6];
    ele[9][6] != ele[13][6];
    ele[9][6] != ele[14][6];
    ele[9][6] != ele[15][6];
    ele[9][6] != ele[9][10];
    ele[9][6] != ele[9][11];
    ele[9][6] != ele[9][12];
    ele[9][6] != ele[9][13];
    ele[9][6] != ele[9][14];
    ele[9][6] != ele[9][15];
    ele[9][6] != ele[9][7];
    ele[9][6] != ele[9][8];
    ele[9][6] != ele[9][9];
    ele[9][7] != ele[10][4];
    ele[9][7] != ele[10][5];
    ele[9][7] != ele[10][6];
    ele[9][7] != ele[10][7];
    ele[9][7] != ele[11][4];
    ele[9][7] != ele[11][5];
    ele[9][7] != ele[11][6];
    ele[9][7] != ele[11][7];
    ele[9][7] != ele[12][7];
    ele[9][7] != ele[13][7];
    ele[9][7] != ele[14][7];
    ele[9][7] != ele[15][7];
    ele[9][7] != ele[9][10];
    ele[9][7] != ele[9][11];
    ele[9][7] != ele[9][12];
    ele[9][7] != ele[9][13];
    ele[9][7] != ele[9][14];
    ele[9][7] != ele[9][15];
    ele[9][7] != ele[9][8];
    ele[9][7] != ele[9][9];
    ele[9][8] != ele[10][10];
    ele[9][8] != ele[10][11];
    ele[9][8] != ele[10][8];
    ele[9][8] != ele[10][9];
    ele[9][8] != ele[11][10];
    ele[9][8] != ele[11][11];
    ele[9][8] != ele[11][8];
    ele[9][8] != ele[11][9];
    ele[9][8] != ele[12][8];
    ele[9][8] != ele[13][8];
    ele[9][8] != ele[14][8];
    ele[9][8] != ele[15][8];
    ele[9][8] != ele[9][10];
    ele[9][8] != ele[9][11];
    ele[9][8] != ele[9][12];
    ele[9][8] != ele[9][13];
    ele[9][8] != ele[9][14];
    ele[9][8] != ele[9][15];
    ele[9][8] != ele[9][9];
    ele[9][9] != ele[10][10];
    ele[9][9] != ele[10][11];
    ele[9][9] != ele[10][8];
    ele[9][9] != ele[10][9];
    ele[9][9] != ele[11][10];
    ele[9][9] != ele[11][11];
    ele[9][9] != ele[11][8];
    ele[9][9] != ele[11][9];
    ele[9][9] != ele[12][9];
    ele[9][9] != ele[13][9];
    ele[9][9] != ele[14][9];
    ele[9][9] != ele[15][9];
    ele[9][9] != ele[9][10];
    ele[9][9] != ele[9][11];
    ele[9][9] != ele[9][12];
    ele[9][9] != ele[9][13];
    ele[9][9] != ele[9][14];
    ele[9][9] != ele[9][15];
  // NUMBER OF CONSTRAINTS: 4992
  }
  function new ();
    if (! this.randomize ()) begin
      $display ("ERROR: Randomization failed...!!!");
    end
  endfunction: new
  function show ();
    $display (ele[0][0], ele[0][1], ele[0][2], ele[0][3], ele[0][4], ele[0][5], ele[0][6], ele[0][7], ele[0][8], ele[0][9], ele[0][10], ele[0][11], ele[0][12], ele[0][13], ele[0][14], ele[0][15]);
    $display (ele[1][0], ele[1][1], ele[1][2], ele[1][3], ele[1][4], ele[1][5], ele[1][6], ele[1][7], ele[1][8], ele[1][9], ele[1][10], ele[1][11], ele[1][12], ele[1][13], ele[1][14], ele[1][15]);
    $display (ele[2][0], ele[2][1], ele[2][2], ele[2][3], ele[2][4], ele[2][5], ele[2][6], ele[2][7], ele[2][8], ele[2][9], ele[2][10], ele[2][11], ele[2][12], ele[2][13], ele[2][14], ele[2][15]);
    $display (ele[3][0], ele[3][1], ele[3][2], ele[3][3], ele[3][4], ele[3][5], ele[3][6], ele[3][7], ele[3][8], ele[3][9], ele[3][10], ele[3][11], ele[3][12], ele[3][13], ele[3][14], ele[3][15]);
    $display (ele[4][0], ele[4][1], ele[4][2], ele[4][3], ele[4][4], ele[4][5], ele[4][6], ele[4][7], ele[4][8], ele[4][9], ele[4][10], ele[4][11], ele[4][12], ele[4][13], ele[4][14], ele[4][15]);
    $display (ele[5][0], ele[5][1], ele[5][2], ele[5][3], ele[5][4], ele[5][5], ele[5][6], ele[5][7], ele[5][8], ele[5][9], ele[5][10], ele[5][11], ele[5][12], ele[5][13], ele[5][14], ele[5][15]);
    $display (ele[6][0], ele[6][1], ele[6][2], ele[6][3], ele[6][4], ele[6][5], ele[6][6], ele[6][7], ele[6][8], ele[6][9], ele[6][10], ele[6][11], ele[6][12], ele[6][13], ele[6][14], ele[6][15]);
    $display (ele[7][0], ele[7][1], ele[7][2], ele[7][3], ele[7][4], ele[7][5], ele[7][6], ele[7][7], ele[7][8], ele[7][9], ele[7][10], ele[7][11], ele[7][12], ele[7][13], ele[7][14], ele[7][15]);
    $display (ele[8][0], ele[8][1], ele[8][2], ele[8][3], ele[8][4], ele[8][5], ele[8][6], ele[8][7], ele[8][8], ele[8][9], ele[8][10], ele[8][11], ele[8][12], ele[8][13], ele[8][14], ele[8][15]);
    $display (ele[9][0], ele[9][1], ele[9][2], ele[9][3], ele[9][4], ele[9][5], ele[9][6], ele[9][7], ele[9][8], ele[9][9], ele[9][10], ele[9][11], ele[9][12], ele[9][13], ele[9][14], ele[9][15]);
    $display (ele[10][0], ele[10][1], ele[10][2], ele[10][3], ele[10][4], ele[10][5], ele[10][6], ele[10][7], ele[10][8], ele[10][9], ele[10][10], ele[10][11], ele[10][12], ele[10][13], ele[10][14], ele[10][15]);
    $display (ele[11][0], ele[11][1], ele[11][2], ele[11][3], ele[11][4], ele[11][5], ele[11][6], ele[11][7], ele[11][8], ele[11][9], ele[11][10], ele[11][11], ele[11][12], ele[11][13], ele[11][14], ele[11][15]);
    $display (ele[12][0], ele[12][1], ele[12][2], ele[12][3], ele[12][4], ele[12][5], ele[12][6], ele[12][7], ele[12][8], ele[12][9], ele[12][10], ele[12][11], ele[12][12], ele[12][13], ele[12][14], ele[12][15]);
    $display (ele[13][0], ele[13][1], ele[13][2], ele[13][3], ele[13][4], ele[13][5], ele[13][6], ele[13][7], ele[13][8], ele[13][9], ele[13][10], ele[13][11], ele[13][12], ele[13][13], ele[13][14], ele[13][15]);
    $display (ele[14][0], ele[14][1], ele[14][2], ele[14][3], ele[14][4], ele[14][5], ele[14][6], ele[14][7], ele[14][8], ele[14][9], ele[14][10], ele[14][11], ele[14][12], ele[14][13], ele[14][14], ele[14][15]);
    $display (ele[15][0], ele[15][1], ele[15][2], ele[15][3], ele[15][4], ele[15][5], ele[15][6], ele[15][7], ele[15][8], ele[15][9], ele[15][10], ele[15][11], ele[15][12], ele[15][13], ele[15][14], ele[15][15]);
  endfunction: show
endclass: board
