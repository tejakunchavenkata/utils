class board;
  typedef enum {
    AAA=1,
    AAB=2,
    AAC=3,
    AAD=4,
    AAE=5,
    AAF=6,
    AAG=7,
    AAH=8,
    AAI=9,
    AAJ=10,
    AAK=11,
    AAL=12,
    AAM=13,
    AAN=14,
    AAO=15,
    AAP=16,
    AAQ=17,
    AAR=18,
    AAS=19,
    AAT=20,
    AAU=21,
    AAV=22,
    AAW=23,
    AAX=24,
    AAY=25,
    AAZ=26,
    ABA=27,
    ABB=28,
    ABC=29,
    ABD=30,
    ABE=31,
    ABF=32,
    ABG=33,
    ABH=34,
    ABI=35,
    ABJ
  } elements;
  rand elements ele[36][36];
  constraint all {
    ele[0][0] != ele[0][1];
    ele[0][0] != ele[0][10];
    ele[0][0] != ele[0][11];
    ele[0][0] != ele[0][12];
    ele[0][0] != ele[0][13];
    ele[0][0] != ele[0][14];
    ele[0][0] != ele[0][15];
    ele[0][0] != ele[0][16];
    ele[0][0] != ele[0][17];
    ele[0][0] != ele[0][18];
    ele[0][0] != ele[0][19];
    ele[0][0] != ele[0][2];
    ele[0][0] != ele[0][20];
    ele[0][0] != ele[0][21];
    ele[0][0] != ele[0][22];
    ele[0][0] != ele[0][23];
    ele[0][0] != ele[0][24];
    ele[0][0] != ele[0][25];
    ele[0][0] != ele[0][26];
    ele[0][0] != ele[0][27];
    ele[0][0] != ele[0][28];
    ele[0][0] != ele[0][29];
    ele[0][0] != ele[0][3];
    ele[0][0] != ele[0][30];
    ele[0][0] != ele[0][31];
    ele[0][0] != ele[0][32];
    ele[0][0] != ele[0][33];
    ele[0][0] != ele[0][34];
    ele[0][0] != ele[0][35];
    ele[0][0] != ele[0][4];
    ele[0][0] != ele[0][5];
    ele[0][0] != ele[0][6];
    ele[0][0] != ele[0][7];
    ele[0][0] != ele[0][8];
    ele[0][0] != ele[0][9];
    ele[0][0] != ele[1][0];
    ele[0][0] != ele[1][1];
    ele[0][0] != ele[1][2];
    ele[0][0] != ele[1][3];
    ele[0][0] != ele[1][4];
    ele[0][0] != ele[1][5];
    ele[0][0] != ele[10][0];
    ele[0][0] != ele[11][0];
    ele[0][0] != ele[12][0];
    ele[0][0] != ele[13][0];
    ele[0][0] != ele[14][0];
    ele[0][0] != ele[15][0];
    ele[0][0] != ele[16][0];
    ele[0][0] != ele[17][0];
    ele[0][0] != ele[18][0];
    ele[0][0] != ele[19][0];
    ele[0][0] != ele[2][0];
    ele[0][0] != ele[2][1];
    ele[0][0] != ele[2][2];
    ele[0][0] != ele[2][3];
    ele[0][0] != ele[2][4];
    ele[0][0] != ele[2][5];
    ele[0][0] != ele[20][0];
    ele[0][0] != ele[21][0];
    ele[0][0] != ele[22][0];
    ele[0][0] != ele[23][0];
    ele[0][0] != ele[24][0];
    ele[0][0] != ele[25][0];
    ele[0][0] != ele[26][0];
    ele[0][0] != ele[27][0];
    ele[0][0] != ele[28][0];
    ele[0][0] != ele[29][0];
    ele[0][0] != ele[3][0];
    ele[0][0] != ele[3][1];
    ele[0][0] != ele[3][2];
    ele[0][0] != ele[3][3];
    ele[0][0] != ele[3][4];
    ele[0][0] != ele[3][5];
    ele[0][0] != ele[30][0];
    ele[0][0] != ele[31][0];
    ele[0][0] != ele[32][0];
    ele[0][0] != ele[33][0];
    ele[0][0] != ele[34][0];
    ele[0][0] != ele[35][0];
    ele[0][0] != ele[4][0];
    ele[0][0] != ele[4][1];
    ele[0][0] != ele[4][2];
    ele[0][0] != ele[4][3];
    ele[0][0] != ele[4][4];
    ele[0][0] != ele[4][5];
    ele[0][0] != ele[5][0];
    ele[0][0] != ele[5][1];
    ele[0][0] != ele[5][2];
    ele[0][0] != ele[5][3];
    ele[0][0] != ele[5][4];
    ele[0][0] != ele[5][5];
    ele[0][0] != ele[6][0];
    ele[0][0] != ele[7][0];
    ele[0][0] != ele[8][0];
    ele[0][0] != ele[9][0];
    ele[0][1] != ele[0][10];
    ele[0][1] != ele[0][11];
    ele[0][1] != ele[0][12];
    ele[0][1] != ele[0][13];
    ele[0][1] != ele[0][14];
    ele[0][1] != ele[0][15];
    ele[0][1] != ele[0][16];
    ele[0][1] != ele[0][17];
    ele[0][1] != ele[0][18];
    ele[0][1] != ele[0][19];
    ele[0][1] != ele[0][2];
    ele[0][1] != ele[0][20];
    ele[0][1] != ele[0][21];
    ele[0][1] != ele[0][22];
    ele[0][1] != ele[0][23];
    ele[0][1] != ele[0][24];
    ele[0][1] != ele[0][25];
    ele[0][1] != ele[0][26];
    ele[0][1] != ele[0][27];
    ele[0][1] != ele[0][28];
    ele[0][1] != ele[0][29];
    ele[0][1] != ele[0][3];
    ele[0][1] != ele[0][30];
    ele[0][1] != ele[0][31];
    ele[0][1] != ele[0][32];
    ele[0][1] != ele[0][33];
    ele[0][1] != ele[0][34];
    ele[0][1] != ele[0][35];
    ele[0][1] != ele[0][4];
    ele[0][1] != ele[0][5];
    ele[0][1] != ele[0][6];
    ele[0][1] != ele[0][7];
    ele[0][1] != ele[0][8];
    ele[0][1] != ele[0][9];
    ele[0][1] != ele[1][0];
    ele[0][1] != ele[1][1];
    ele[0][1] != ele[1][2];
    ele[0][1] != ele[1][3];
    ele[0][1] != ele[1][4];
    ele[0][1] != ele[1][5];
    ele[0][1] != ele[10][1];
    ele[0][1] != ele[11][1];
    ele[0][1] != ele[12][1];
    ele[0][1] != ele[13][1];
    ele[0][1] != ele[14][1];
    ele[0][1] != ele[15][1];
    ele[0][1] != ele[16][1];
    ele[0][1] != ele[17][1];
    ele[0][1] != ele[18][1];
    ele[0][1] != ele[19][1];
    ele[0][1] != ele[2][0];
    ele[0][1] != ele[2][1];
    ele[0][1] != ele[2][2];
    ele[0][1] != ele[2][3];
    ele[0][1] != ele[2][4];
    ele[0][1] != ele[2][5];
    ele[0][1] != ele[20][1];
    ele[0][1] != ele[21][1];
    ele[0][1] != ele[22][1];
    ele[0][1] != ele[23][1];
    ele[0][1] != ele[24][1];
    ele[0][1] != ele[25][1];
    ele[0][1] != ele[26][1];
    ele[0][1] != ele[27][1];
    ele[0][1] != ele[28][1];
    ele[0][1] != ele[29][1];
    ele[0][1] != ele[3][0];
    ele[0][1] != ele[3][1];
    ele[0][1] != ele[3][2];
    ele[0][1] != ele[3][3];
    ele[0][1] != ele[3][4];
    ele[0][1] != ele[3][5];
    ele[0][1] != ele[30][1];
    ele[0][1] != ele[31][1];
    ele[0][1] != ele[32][1];
    ele[0][1] != ele[33][1];
    ele[0][1] != ele[34][1];
    ele[0][1] != ele[35][1];
    ele[0][1] != ele[4][0];
    ele[0][1] != ele[4][1];
    ele[0][1] != ele[4][2];
    ele[0][1] != ele[4][3];
    ele[0][1] != ele[4][4];
    ele[0][1] != ele[4][5];
    ele[0][1] != ele[5][0];
    ele[0][1] != ele[5][1];
    ele[0][1] != ele[5][2];
    ele[0][1] != ele[5][3];
    ele[0][1] != ele[5][4];
    ele[0][1] != ele[5][5];
    ele[0][1] != ele[6][1];
    ele[0][1] != ele[7][1];
    ele[0][1] != ele[8][1];
    ele[0][1] != ele[9][1];
    ele[0][10] != ele[0][11];
    ele[0][10] != ele[0][12];
    ele[0][10] != ele[0][13];
    ele[0][10] != ele[0][14];
    ele[0][10] != ele[0][15];
    ele[0][10] != ele[0][16];
    ele[0][10] != ele[0][17];
    ele[0][10] != ele[0][18];
    ele[0][10] != ele[0][19];
    ele[0][10] != ele[0][20];
    ele[0][10] != ele[0][21];
    ele[0][10] != ele[0][22];
    ele[0][10] != ele[0][23];
    ele[0][10] != ele[0][24];
    ele[0][10] != ele[0][25];
    ele[0][10] != ele[0][26];
    ele[0][10] != ele[0][27];
    ele[0][10] != ele[0][28];
    ele[0][10] != ele[0][29];
    ele[0][10] != ele[0][30];
    ele[0][10] != ele[0][31];
    ele[0][10] != ele[0][32];
    ele[0][10] != ele[0][33];
    ele[0][10] != ele[0][34];
    ele[0][10] != ele[0][35];
    ele[0][10] != ele[1][10];
    ele[0][10] != ele[1][11];
    ele[0][10] != ele[1][6];
    ele[0][10] != ele[1][7];
    ele[0][10] != ele[1][8];
    ele[0][10] != ele[1][9];
    ele[0][10] != ele[10][10];
    ele[0][10] != ele[11][10];
    ele[0][10] != ele[12][10];
    ele[0][10] != ele[13][10];
    ele[0][10] != ele[14][10];
    ele[0][10] != ele[15][10];
    ele[0][10] != ele[16][10];
    ele[0][10] != ele[17][10];
    ele[0][10] != ele[18][10];
    ele[0][10] != ele[19][10];
    ele[0][10] != ele[2][10];
    ele[0][10] != ele[2][11];
    ele[0][10] != ele[2][6];
    ele[0][10] != ele[2][7];
    ele[0][10] != ele[2][8];
    ele[0][10] != ele[2][9];
    ele[0][10] != ele[20][10];
    ele[0][10] != ele[21][10];
    ele[0][10] != ele[22][10];
    ele[0][10] != ele[23][10];
    ele[0][10] != ele[24][10];
    ele[0][10] != ele[25][10];
    ele[0][10] != ele[26][10];
    ele[0][10] != ele[27][10];
    ele[0][10] != ele[28][10];
    ele[0][10] != ele[29][10];
    ele[0][10] != ele[3][10];
    ele[0][10] != ele[3][11];
    ele[0][10] != ele[3][6];
    ele[0][10] != ele[3][7];
    ele[0][10] != ele[3][8];
    ele[0][10] != ele[3][9];
    ele[0][10] != ele[30][10];
    ele[0][10] != ele[31][10];
    ele[0][10] != ele[32][10];
    ele[0][10] != ele[33][10];
    ele[0][10] != ele[34][10];
    ele[0][10] != ele[35][10];
    ele[0][10] != ele[4][10];
    ele[0][10] != ele[4][11];
    ele[0][10] != ele[4][6];
    ele[0][10] != ele[4][7];
    ele[0][10] != ele[4][8];
    ele[0][10] != ele[4][9];
    ele[0][10] != ele[5][10];
    ele[0][10] != ele[5][11];
    ele[0][10] != ele[5][6];
    ele[0][10] != ele[5][7];
    ele[0][10] != ele[5][8];
    ele[0][10] != ele[5][9];
    ele[0][10] != ele[6][10];
    ele[0][10] != ele[7][10];
    ele[0][10] != ele[8][10];
    ele[0][10] != ele[9][10];
    ele[0][11] != ele[0][12];
    ele[0][11] != ele[0][13];
    ele[0][11] != ele[0][14];
    ele[0][11] != ele[0][15];
    ele[0][11] != ele[0][16];
    ele[0][11] != ele[0][17];
    ele[0][11] != ele[0][18];
    ele[0][11] != ele[0][19];
    ele[0][11] != ele[0][20];
    ele[0][11] != ele[0][21];
    ele[0][11] != ele[0][22];
    ele[0][11] != ele[0][23];
    ele[0][11] != ele[0][24];
    ele[0][11] != ele[0][25];
    ele[0][11] != ele[0][26];
    ele[0][11] != ele[0][27];
    ele[0][11] != ele[0][28];
    ele[0][11] != ele[0][29];
    ele[0][11] != ele[0][30];
    ele[0][11] != ele[0][31];
    ele[0][11] != ele[0][32];
    ele[0][11] != ele[0][33];
    ele[0][11] != ele[0][34];
    ele[0][11] != ele[0][35];
    ele[0][11] != ele[1][10];
    ele[0][11] != ele[1][11];
    ele[0][11] != ele[1][6];
    ele[0][11] != ele[1][7];
    ele[0][11] != ele[1][8];
    ele[0][11] != ele[1][9];
    ele[0][11] != ele[10][11];
    ele[0][11] != ele[11][11];
    ele[0][11] != ele[12][11];
    ele[0][11] != ele[13][11];
    ele[0][11] != ele[14][11];
    ele[0][11] != ele[15][11];
    ele[0][11] != ele[16][11];
    ele[0][11] != ele[17][11];
    ele[0][11] != ele[18][11];
    ele[0][11] != ele[19][11];
    ele[0][11] != ele[2][10];
    ele[0][11] != ele[2][11];
    ele[0][11] != ele[2][6];
    ele[0][11] != ele[2][7];
    ele[0][11] != ele[2][8];
    ele[0][11] != ele[2][9];
    ele[0][11] != ele[20][11];
    ele[0][11] != ele[21][11];
    ele[0][11] != ele[22][11];
    ele[0][11] != ele[23][11];
    ele[0][11] != ele[24][11];
    ele[0][11] != ele[25][11];
    ele[0][11] != ele[26][11];
    ele[0][11] != ele[27][11];
    ele[0][11] != ele[28][11];
    ele[0][11] != ele[29][11];
    ele[0][11] != ele[3][10];
    ele[0][11] != ele[3][11];
    ele[0][11] != ele[3][6];
    ele[0][11] != ele[3][7];
    ele[0][11] != ele[3][8];
    ele[0][11] != ele[3][9];
    ele[0][11] != ele[30][11];
    ele[0][11] != ele[31][11];
    ele[0][11] != ele[32][11];
    ele[0][11] != ele[33][11];
    ele[0][11] != ele[34][11];
    ele[0][11] != ele[35][11];
    ele[0][11] != ele[4][10];
    ele[0][11] != ele[4][11];
    ele[0][11] != ele[4][6];
    ele[0][11] != ele[4][7];
    ele[0][11] != ele[4][8];
    ele[0][11] != ele[4][9];
    ele[0][11] != ele[5][10];
    ele[0][11] != ele[5][11];
    ele[0][11] != ele[5][6];
    ele[0][11] != ele[5][7];
    ele[0][11] != ele[5][8];
    ele[0][11] != ele[5][9];
    ele[0][11] != ele[6][11];
    ele[0][11] != ele[7][11];
    ele[0][11] != ele[8][11];
    ele[0][11] != ele[9][11];
    ele[0][12] != ele[0][13];
    ele[0][12] != ele[0][14];
    ele[0][12] != ele[0][15];
    ele[0][12] != ele[0][16];
    ele[0][12] != ele[0][17];
    ele[0][12] != ele[0][18];
    ele[0][12] != ele[0][19];
    ele[0][12] != ele[0][20];
    ele[0][12] != ele[0][21];
    ele[0][12] != ele[0][22];
    ele[0][12] != ele[0][23];
    ele[0][12] != ele[0][24];
    ele[0][12] != ele[0][25];
    ele[0][12] != ele[0][26];
    ele[0][12] != ele[0][27];
    ele[0][12] != ele[0][28];
    ele[0][12] != ele[0][29];
    ele[0][12] != ele[0][30];
    ele[0][12] != ele[0][31];
    ele[0][12] != ele[0][32];
    ele[0][12] != ele[0][33];
    ele[0][12] != ele[0][34];
    ele[0][12] != ele[0][35];
    ele[0][12] != ele[1][12];
    ele[0][12] != ele[1][13];
    ele[0][12] != ele[1][14];
    ele[0][12] != ele[1][15];
    ele[0][12] != ele[1][16];
    ele[0][12] != ele[1][17];
    ele[0][12] != ele[10][12];
    ele[0][12] != ele[11][12];
    ele[0][12] != ele[12][12];
    ele[0][12] != ele[13][12];
    ele[0][12] != ele[14][12];
    ele[0][12] != ele[15][12];
    ele[0][12] != ele[16][12];
    ele[0][12] != ele[17][12];
    ele[0][12] != ele[18][12];
    ele[0][12] != ele[19][12];
    ele[0][12] != ele[2][12];
    ele[0][12] != ele[2][13];
    ele[0][12] != ele[2][14];
    ele[0][12] != ele[2][15];
    ele[0][12] != ele[2][16];
    ele[0][12] != ele[2][17];
    ele[0][12] != ele[20][12];
    ele[0][12] != ele[21][12];
    ele[0][12] != ele[22][12];
    ele[0][12] != ele[23][12];
    ele[0][12] != ele[24][12];
    ele[0][12] != ele[25][12];
    ele[0][12] != ele[26][12];
    ele[0][12] != ele[27][12];
    ele[0][12] != ele[28][12];
    ele[0][12] != ele[29][12];
    ele[0][12] != ele[3][12];
    ele[0][12] != ele[3][13];
    ele[0][12] != ele[3][14];
    ele[0][12] != ele[3][15];
    ele[0][12] != ele[3][16];
    ele[0][12] != ele[3][17];
    ele[0][12] != ele[30][12];
    ele[0][12] != ele[31][12];
    ele[0][12] != ele[32][12];
    ele[0][12] != ele[33][12];
    ele[0][12] != ele[34][12];
    ele[0][12] != ele[35][12];
    ele[0][12] != ele[4][12];
    ele[0][12] != ele[4][13];
    ele[0][12] != ele[4][14];
    ele[0][12] != ele[4][15];
    ele[0][12] != ele[4][16];
    ele[0][12] != ele[4][17];
    ele[0][12] != ele[5][12];
    ele[0][12] != ele[5][13];
    ele[0][12] != ele[5][14];
    ele[0][12] != ele[5][15];
    ele[0][12] != ele[5][16];
    ele[0][12] != ele[5][17];
    ele[0][12] != ele[6][12];
    ele[0][12] != ele[7][12];
    ele[0][12] != ele[8][12];
    ele[0][12] != ele[9][12];
    ele[0][13] != ele[0][14];
    ele[0][13] != ele[0][15];
    ele[0][13] != ele[0][16];
    ele[0][13] != ele[0][17];
    ele[0][13] != ele[0][18];
    ele[0][13] != ele[0][19];
    ele[0][13] != ele[0][20];
    ele[0][13] != ele[0][21];
    ele[0][13] != ele[0][22];
    ele[0][13] != ele[0][23];
    ele[0][13] != ele[0][24];
    ele[0][13] != ele[0][25];
    ele[0][13] != ele[0][26];
    ele[0][13] != ele[0][27];
    ele[0][13] != ele[0][28];
    ele[0][13] != ele[0][29];
    ele[0][13] != ele[0][30];
    ele[0][13] != ele[0][31];
    ele[0][13] != ele[0][32];
    ele[0][13] != ele[0][33];
    ele[0][13] != ele[0][34];
    ele[0][13] != ele[0][35];
    ele[0][13] != ele[1][12];
    ele[0][13] != ele[1][13];
    ele[0][13] != ele[1][14];
    ele[0][13] != ele[1][15];
    ele[0][13] != ele[1][16];
    ele[0][13] != ele[1][17];
    ele[0][13] != ele[10][13];
    ele[0][13] != ele[11][13];
    ele[0][13] != ele[12][13];
    ele[0][13] != ele[13][13];
    ele[0][13] != ele[14][13];
    ele[0][13] != ele[15][13];
    ele[0][13] != ele[16][13];
    ele[0][13] != ele[17][13];
    ele[0][13] != ele[18][13];
    ele[0][13] != ele[19][13];
    ele[0][13] != ele[2][12];
    ele[0][13] != ele[2][13];
    ele[0][13] != ele[2][14];
    ele[0][13] != ele[2][15];
    ele[0][13] != ele[2][16];
    ele[0][13] != ele[2][17];
    ele[0][13] != ele[20][13];
    ele[0][13] != ele[21][13];
    ele[0][13] != ele[22][13];
    ele[0][13] != ele[23][13];
    ele[0][13] != ele[24][13];
    ele[0][13] != ele[25][13];
    ele[0][13] != ele[26][13];
    ele[0][13] != ele[27][13];
    ele[0][13] != ele[28][13];
    ele[0][13] != ele[29][13];
    ele[0][13] != ele[3][12];
    ele[0][13] != ele[3][13];
    ele[0][13] != ele[3][14];
    ele[0][13] != ele[3][15];
    ele[0][13] != ele[3][16];
    ele[0][13] != ele[3][17];
    ele[0][13] != ele[30][13];
    ele[0][13] != ele[31][13];
    ele[0][13] != ele[32][13];
    ele[0][13] != ele[33][13];
    ele[0][13] != ele[34][13];
    ele[0][13] != ele[35][13];
    ele[0][13] != ele[4][12];
    ele[0][13] != ele[4][13];
    ele[0][13] != ele[4][14];
    ele[0][13] != ele[4][15];
    ele[0][13] != ele[4][16];
    ele[0][13] != ele[4][17];
    ele[0][13] != ele[5][12];
    ele[0][13] != ele[5][13];
    ele[0][13] != ele[5][14];
    ele[0][13] != ele[5][15];
    ele[0][13] != ele[5][16];
    ele[0][13] != ele[5][17];
    ele[0][13] != ele[6][13];
    ele[0][13] != ele[7][13];
    ele[0][13] != ele[8][13];
    ele[0][13] != ele[9][13];
    ele[0][14] != ele[0][15];
    ele[0][14] != ele[0][16];
    ele[0][14] != ele[0][17];
    ele[0][14] != ele[0][18];
    ele[0][14] != ele[0][19];
    ele[0][14] != ele[0][20];
    ele[0][14] != ele[0][21];
    ele[0][14] != ele[0][22];
    ele[0][14] != ele[0][23];
    ele[0][14] != ele[0][24];
    ele[0][14] != ele[0][25];
    ele[0][14] != ele[0][26];
    ele[0][14] != ele[0][27];
    ele[0][14] != ele[0][28];
    ele[0][14] != ele[0][29];
    ele[0][14] != ele[0][30];
    ele[0][14] != ele[0][31];
    ele[0][14] != ele[0][32];
    ele[0][14] != ele[0][33];
    ele[0][14] != ele[0][34];
    ele[0][14] != ele[0][35];
    ele[0][14] != ele[1][12];
    ele[0][14] != ele[1][13];
    ele[0][14] != ele[1][14];
    ele[0][14] != ele[1][15];
    ele[0][14] != ele[1][16];
    ele[0][14] != ele[1][17];
    ele[0][14] != ele[10][14];
    ele[0][14] != ele[11][14];
    ele[0][14] != ele[12][14];
    ele[0][14] != ele[13][14];
    ele[0][14] != ele[14][14];
    ele[0][14] != ele[15][14];
    ele[0][14] != ele[16][14];
    ele[0][14] != ele[17][14];
    ele[0][14] != ele[18][14];
    ele[0][14] != ele[19][14];
    ele[0][14] != ele[2][12];
    ele[0][14] != ele[2][13];
    ele[0][14] != ele[2][14];
    ele[0][14] != ele[2][15];
    ele[0][14] != ele[2][16];
    ele[0][14] != ele[2][17];
    ele[0][14] != ele[20][14];
    ele[0][14] != ele[21][14];
    ele[0][14] != ele[22][14];
    ele[0][14] != ele[23][14];
    ele[0][14] != ele[24][14];
    ele[0][14] != ele[25][14];
    ele[0][14] != ele[26][14];
    ele[0][14] != ele[27][14];
    ele[0][14] != ele[28][14];
    ele[0][14] != ele[29][14];
    ele[0][14] != ele[3][12];
    ele[0][14] != ele[3][13];
    ele[0][14] != ele[3][14];
    ele[0][14] != ele[3][15];
    ele[0][14] != ele[3][16];
    ele[0][14] != ele[3][17];
    ele[0][14] != ele[30][14];
    ele[0][14] != ele[31][14];
    ele[0][14] != ele[32][14];
    ele[0][14] != ele[33][14];
    ele[0][14] != ele[34][14];
    ele[0][14] != ele[35][14];
    ele[0][14] != ele[4][12];
    ele[0][14] != ele[4][13];
    ele[0][14] != ele[4][14];
    ele[0][14] != ele[4][15];
    ele[0][14] != ele[4][16];
    ele[0][14] != ele[4][17];
    ele[0][14] != ele[5][12];
    ele[0][14] != ele[5][13];
    ele[0][14] != ele[5][14];
    ele[0][14] != ele[5][15];
    ele[0][14] != ele[5][16];
    ele[0][14] != ele[5][17];
    ele[0][14] != ele[6][14];
    ele[0][14] != ele[7][14];
    ele[0][14] != ele[8][14];
    ele[0][14] != ele[9][14];
    ele[0][15] != ele[0][16];
    ele[0][15] != ele[0][17];
    ele[0][15] != ele[0][18];
    ele[0][15] != ele[0][19];
    ele[0][15] != ele[0][20];
    ele[0][15] != ele[0][21];
    ele[0][15] != ele[0][22];
    ele[0][15] != ele[0][23];
    ele[0][15] != ele[0][24];
    ele[0][15] != ele[0][25];
    ele[0][15] != ele[0][26];
    ele[0][15] != ele[0][27];
    ele[0][15] != ele[0][28];
    ele[0][15] != ele[0][29];
    ele[0][15] != ele[0][30];
    ele[0][15] != ele[0][31];
    ele[0][15] != ele[0][32];
    ele[0][15] != ele[0][33];
    ele[0][15] != ele[0][34];
    ele[0][15] != ele[0][35];
    ele[0][15] != ele[1][12];
    ele[0][15] != ele[1][13];
    ele[0][15] != ele[1][14];
    ele[0][15] != ele[1][15];
    ele[0][15] != ele[1][16];
    ele[0][15] != ele[1][17];
    ele[0][15] != ele[10][15];
    ele[0][15] != ele[11][15];
    ele[0][15] != ele[12][15];
    ele[0][15] != ele[13][15];
    ele[0][15] != ele[14][15];
    ele[0][15] != ele[15][15];
    ele[0][15] != ele[16][15];
    ele[0][15] != ele[17][15];
    ele[0][15] != ele[18][15];
    ele[0][15] != ele[19][15];
    ele[0][15] != ele[2][12];
    ele[0][15] != ele[2][13];
    ele[0][15] != ele[2][14];
    ele[0][15] != ele[2][15];
    ele[0][15] != ele[2][16];
    ele[0][15] != ele[2][17];
    ele[0][15] != ele[20][15];
    ele[0][15] != ele[21][15];
    ele[0][15] != ele[22][15];
    ele[0][15] != ele[23][15];
    ele[0][15] != ele[24][15];
    ele[0][15] != ele[25][15];
    ele[0][15] != ele[26][15];
    ele[0][15] != ele[27][15];
    ele[0][15] != ele[28][15];
    ele[0][15] != ele[29][15];
    ele[0][15] != ele[3][12];
    ele[0][15] != ele[3][13];
    ele[0][15] != ele[3][14];
    ele[0][15] != ele[3][15];
    ele[0][15] != ele[3][16];
    ele[0][15] != ele[3][17];
    ele[0][15] != ele[30][15];
    ele[0][15] != ele[31][15];
    ele[0][15] != ele[32][15];
    ele[0][15] != ele[33][15];
    ele[0][15] != ele[34][15];
    ele[0][15] != ele[35][15];
    ele[0][15] != ele[4][12];
    ele[0][15] != ele[4][13];
    ele[0][15] != ele[4][14];
    ele[0][15] != ele[4][15];
    ele[0][15] != ele[4][16];
    ele[0][15] != ele[4][17];
    ele[0][15] != ele[5][12];
    ele[0][15] != ele[5][13];
    ele[0][15] != ele[5][14];
    ele[0][15] != ele[5][15];
    ele[0][15] != ele[5][16];
    ele[0][15] != ele[5][17];
    ele[0][15] != ele[6][15];
    ele[0][15] != ele[7][15];
    ele[0][15] != ele[8][15];
    ele[0][15] != ele[9][15];
    ele[0][16] != ele[0][17];
    ele[0][16] != ele[0][18];
    ele[0][16] != ele[0][19];
    ele[0][16] != ele[0][20];
    ele[0][16] != ele[0][21];
    ele[0][16] != ele[0][22];
    ele[0][16] != ele[0][23];
    ele[0][16] != ele[0][24];
    ele[0][16] != ele[0][25];
    ele[0][16] != ele[0][26];
    ele[0][16] != ele[0][27];
    ele[0][16] != ele[0][28];
    ele[0][16] != ele[0][29];
    ele[0][16] != ele[0][30];
    ele[0][16] != ele[0][31];
    ele[0][16] != ele[0][32];
    ele[0][16] != ele[0][33];
    ele[0][16] != ele[0][34];
    ele[0][16] != ele[0][35];
    ele[0][16] != ele[1][12];
    ele[0][16] != ele[1][13];
    ele[0][16] != ele[1][14];
    ele[0][16] != ele[1][15];
    ele[0][16] != ele[1][16];
    ele[0][16] != ele[1][17];
    ele[0][16] != ele[10][16];
    ele[0][16] != ele[11][16];
    ele[0][16] != ele[12][16];
    ele[0][16] != ele[13][16];
    ele[0][16] != ele[14][16];
    ele[0][16] != ele[15][16];
    ele[0][16] != ele[16][16];
    ele[0][16] != ele[17][16];
    ele[0][16] != ele[18][16];
    ele[0][16] != ele[19][16];
    ele[0][16] != ele[2][12];
    ele[0][16] != ele[2][13];
    ele[0][16] != ele[2][14];
    ele[0][16] != ele[2][15];
    ele[0][16] != ele[2][16];
    ele[0][16] != ele[2][17];
    ele[0][16] != ele[20][16];
    ele[0][16] != ele[21][16];
    ele[0][16] != ele[22][16];
    ele[0][16] != ele[23][16];
    ele[0][16] != ele[24][16];
    ele[0][16] != ele[25][16];
    ele[0][16] != ele[26][16];
    ele[0][16] != ele[27][16];
    ele[0][16] != ele[28][16];
    ele[0][16] != ele[29][16];
    ele[0][16] != ele[3][12];
    ele[0][16] != ele[3][13];
    ele[0][16] != ele[3][14];
    ele[0][16] != ele[3][15];
    ele[0][16] != ele[3][16];
    ele[0][16] != ele[3][17];
    ele[0][16] != ele[30][16];
    ele[0][16] != ele[31][16];
    ele[0][16] != ele[32][16];
    ele[0][16] != ele[33][16];
    ele[0][16] != ele[34][16];
    ele[0][16] != ele[35][16];
    ele[0][16] != ele[4][12];
    ele[0][16] != ele[4][13];
    ele[0][16] != ele[4][14];
    ele[0][16] != ele[4][15];
    ele[0][16] != ele[4][16];
    ele[0][16] != ele[4][17];
    ele[0][16] != ele[5][12];
    ele[0][16] != ele[5][13];
    ele[0][16] != ele[5][14];
    ele[0][16] != ele[5][15];
    ele[0][16] != ele[5][16];
    ele[0][16] != ele[5][17];
    ele[0][16] != ele[6][16];
    ele[0][16] != ele[7][16];
    ele[0][16] != ele[8][16];
    ele[0][16] != ele[9][16];
    ele[0][17] != ele[0][18];
    ele[0][17] != ele[0][19];
    ele[0][17] != ele[0][20];
    ele[0][17] != ele[0][21];
    ele[0][17] != ele[0][22];
    ele[0][17] != ele[0][23];
    ele[0][17] != ele[0][24];
    ele[0][17] != ele[0][25];
    ele[0][17] != ele[0][26];
    ele[0][17] != ele[0][27];
    ele[0][17] != ele[0][28];
    ele[0][17] != ele[0][29];
    ele[0][17] != ele[0][30];
    ele[0][17] != ele[0][31];
    ele[0][17] != ele[0][32];
    ele[0][17] != ele[0][33];
    ele[0][17] != ele[0][34];
    ele[0][17] != ele[0][35];
    ele[0][17] != ele[1][12];
    ele[0][17] != ele[1][13];
    ele[0][17] != ele[1][14];
    ele[0][17] != ele[1][15];
    ele[0][17] != ele[1][16];
    ele[0][17] != ele[1][17];
    ele[0][17] != ele[10][17];
    ele[0][17] != ele[11][17];
    ele[0][17] != ele[12][17];
    ele[0][17] != ele[13][17];
    ele[0][17] != ele[14][17];
    ele[0][17] != ele[15][17];
    ele[0][17] != ele[16][17];
    ele[0][17] != ele[17][17];
    ele[0][17] != ele[18][17];
    ele[0][17] != ele[19][17];
    ele[0][17] != ele[2][12];
    ele[0][17] != ele[2][13];
    ele[0][17] != ele[2][14];
    ele[0][17] != ele[2][15];
    ele[0][17] != ele[2][16];
    ele[0][17] != ele[2][17];
    ele[0][17] != ele[20][17];
    ele[0][17] != ele[21][17];
    ele[0][17] != ele[22][17];
    ele[0][17] != ele[23][17];
    ele[0][17] != ele[24][17];
    ele[0][17] != ele[25][17];
    ele[0][17] != ele[26][17];
    ele[0][17] != ele[27][17];
    ele[0][17] != ele[28][17];
    ele[0][17] != ele[29][17];
    ele[0][17] != ele[3][12];
    ele[0][17] != ele[3][13];
    ele[0][17] != ele[3][14];
    ele[0][17] != ele[3][15];
    ele[0][17] != ele[3][16];
    ele[0][17] != ele[3][17];
    ele[0][17] != ele[30][17];
    ele[0][17] != ele[31][17];
    ele[0][17] != ele[32][17];
    ele[0][17] != ele[33][17];
    ele[0][17] != ele[34][17];
    ele[0][17] != ele[35][17];
    ele[0][17] != ele[4][12];
    ele[0][17] != ele[4][13];
    ele[0][17] != ele[4][14];
    ele[0][17] != ele[4][15];
    ele[0][17] != ele[4][16];
    ele[0][17] != ele[4][17];
    ele[0][17] != ele[5][12];
    ele[0][17] != ele[5][13];
    ele[0][17] != ele[5][14];
    ele[0][17] != ele[5][15];
    ele[0][17] != ele[5][16];
    ele[0][17] != ele[5][17];
    ele[0][17] != ele[6][17];
    ele[0][17] != ele[7][17];
    ele[0][17] != ele[8][17];
    ele[0][17] != ele[9][17];
    ele[0][18] != ele[0][19];
    ele[0][18] != ele[0][20];
    ele[0][18] != ele[0][21];
    ele[0][18] != ele[0][22];
    ele[0][18] != ele[0][23];
    ele[0][18] != ele[0][24];
    ele[0][18] != ele[0][25];
    ele[0][18] != ele[0][26];
    ele[0][18] != ele[0][27];
    ele[0][18] != ele[0][28];
    ele[0][18] != ele[0][29];
    ele[0][18] != ele[0][30];
    ele[0][18] != ele[0][31];
    ele[0][18] != ele[0][32];
    ele[0][18] != ele[0][33];
    ele[0][18] != ele[0][34];
    ele[0][18] != ele[0][35];
    ele[0][18] != ele[1][18];
    ele[0][18] != ele[1][19];
    ele[0][18] != ele[1][20];
    ele[0][18] != ele[1][21];
    ele[0][18] != ele[1][22];
    ele[0][18] != ele[1][23];
    ele[0][18] != ele[10][18];
    ele[0][18] != ele[11][18];
    ele[0][18] != ele[12][18];
    ele[0][18] != ele[13][18];
    ele[0][18] != ele[14][18];
    ele[0][18] != ele[15][18];
    ele[0][18] != ele[16][18];
    ele[0][18] != ele[17][18];
    ele[0][18] != ele[18][18];
    ele[0][18] != ele[19][18];
    ele[0][18] != ele[2][18];
    ele[0][18] != ele[2][19];
    ele[0][18] != ele[2][20];
    ele[0][18] != ele[2][21];
    ele[0][18] != ele[2][22];
    ele[0][18] != ele[2][23];
    ele[0][18] != ele[20][18];
    ele[0][18] != ele[21][18];
    ele[0][18] != ele[22][18];
    ele[0][18] != ele[23][18];
    ele[0][18] != ele[24][18];
    ele[0][18] != ele[25][18];
    ele[0][18] != ele[26][18];
    ele[0][18] != ele[27][18];
    ele[0][18] != ele[28][18];
    ele[0][18] != ele[29][18];
    ele[0][18] != ele[3][18];
    ele[0][18] != ele[3][19];
    ele[0][18] != ele[3][20];
    ele[0][18] != ele[3][21];
    ele[0][18] != ele[3][22];
    ele[0][18] != ele[3][23];
    ele[0][18] != ele[30][18];
    ele[0][18] != ele[31][18];
    ele[0][18] != ele[32][18];
    ele[0][18] != ele[33][18];
    ele[0][18] != ele[34][18];
    ele[0][18] != ele[35][18];
    ele[0][18] != ele[4][18];
    ele[0][18] != ele[4][19];
    ele[0][18] != ele[4][20];
    ele[0][18] != ele[4][21];
    ele[0][18] != ele[4][22];
    ele[0][18] != ele[4][23];
    ele[0][18] != ele[5][18];
    ele[0][18] != ele[5][19];
    ele[0][18] != ele[5][20];
    ele[0][18] != ele[5][21];
    ele[0][18] != ele[5][22];
    ele[0][18] != ele[5][23];
    ele[0][18] != ele[6][18];
    ele[0][18] != ele[7][18];
    ele[0][18] != ele[8][18];
    ele[0][18] != ele[9][18];
    ele[0][19] != ele[0][20];
    ele[0][19] != ele[0][21];
    ele[0][19] != ele[0][22];
    ele[0][19] != ele[0][23];
    ele[0][19] != ele[0][24];
    ele[0][19] != ele[0][25];
    ele[0][19] != ele[0][26];
    ele[0][19] != ele[0][27];
    ele[0][19] != ele[0][28];
    ele[0][19] != ele[0][29];
    ele[0][19] != ele[0][30];
    ele[0][19] != ele[0][31];
    ele[0][19] != ele[0][32];
    ele[0][19] != ele[0][33];
    ele[0][19] != ele[0][34];
    ele[0][19] != ele[0][35];
    ele[0][19] != ele[1][18];
    ele[0][19] != ele[1][19];
    ele[0][19] != ele[1][20];
    ele[0][19] != ele[1][21];
    ele[0][19] != ele[1][22];
    ele[0][19] != ele[1][23];
    ele[0][19] != ele[10][19];
    ele[0][19] != ele[11][19];
    ele[0][19] != ele[12][19];
    ele[0][19] != ele[13][19];
    ele[0][19] != ele[14][19];
    ele[0][19] != ele[15][19];
    ele[0][19] != ele[16][19];
    ele[0][19] != ele[17][19];
    ele[0][19] != ele[18][19];
    ele[0][19] != ele[19][19];
    ele[0][19] != ele[2][18];
    ele[0][19] != ele[2][19];
    ele[0][19] != ele[2][20];
    ele[0][19] != ele[2][21];
    ele[0][19] != ele[2][22];
    ele[0][19] != ele[2][23];
    ele[0][19] != ele[20][19];
    ele[0][19] != ele[21][19];
    ele[0][19] != ele[22][19];
    ele[0][19] != ele[23][19];
    ele[0][19] != ele[24][19];
    ele[0][19] != ele[25][19];
    ele[0][19] != ele[26][19];
    ele[0][19] != ele[27][19];
    ele[0][19] != ele[28][19];
    ele[0][19] != ele[29][19];
    ele[0][19] != ele[3][18];
    ele[0][19] != ele[3][19];
    ele[0][19] != ele[3][20];
    ele[0][19] != ele[3][21];
    ele[0][19] != ele[3][22];
    ele[0][19] != ele[3][23];
    ele[0][19] != ele[30][19];
    ele[0][19] != ele[31][19];
    ele[0][19] != ele[32][19];
    ele[0][19] != ele[33][19];
    ele[0][19] != ele[34][19];
    ele[0][19] != ele[35][19];
    ele[0][19] != ele[4][18];
    ele[0][19] != ele[4][19];
    ele[0][19] != ele[4][20];
    ele[0][19] != ele[4][21];
    ele[0][19] != ele[4][22];
    ele[0][19] != ele[4][23];
    ele[0][19] != ele[5][18];
    ele[0][19] != ele[5][19];
    ele[0][19] != ele[5][20];
    ele[0][19] != ele[5][21];
    ele[0][19] != ele[5][22];
    ele[0][19] != ele[5][23];
    ele[0][19] != ele[6][19];
    ele[0][19] != ele[7][19];
    ele[0][19] != ele[8][19];
    ele[0][19] != ele[9][19];
    ele[0][2] != ele[0][10];
    ele[0][2] != ele[0][11];
    ele[0][2] != ele[0][12];
    ele[0][2] != ele[0][13];
    ele[0][2] != ele[0][14];
    ele[0][2] != ele[0][15];
    ele[0][2] != ele[0][16];
    ele[0][2] != ele[0][17];
    ele[0][2] != ele[0][18];
    ele[0][2] != ele[0][19];
    ele[0][2] != ele[0][20];
    ele[0][2] != ele[0][21];
    ele[0][2] != ele[0][22];
    ele[0][2] != ele[0][23];
    ele[0][2] != ele[0][24];
    ele[0][2] != ele[0][25];
    ele[0][2] != ele[0][26];
    ele[0][2] != ele[0][27];
    ele[0][2] != ele[0][28];
    ele[0][2] != ele[0][29];
    ele[0][2] != ele[0][3];
    ele[0][2] != ele[0][30];
    ele[0][2] != ele[0][31];
    ele[0][2] != ele[0][32];
    ele[0][2] != ele[0][33];
    ele[0][2] != ele[0][34];
    ele[0][2] != ele[0][35];
    ele[0][2] != ele[0][4];
    ele[0][2] != ele[0][5];
    ele[0][2] != ele[0][6];
    ele[0][2] != ele[0][7];
    ele[0][2] != ele[0][8];
    ele[0][2] != ele[0][9];
    ele[0][2] != ele[1][0];
    ele[0][2] != ele[1][1];
    ele[0][2] != ele[1][2];
    ele[0][2] != ele[1][3];
    ele[0][2] != ele[1][4];
    ele[0][2] != ele[1][5];
    ele[0][2] != ele[10][2];
    ele[0][2] != ele[11][2];
    ele[0][2] != ele[12][2];
    ele[0][2] != ele[13][2];
    ele[0][2] != ele[14][2];
    ele[0][2] != ele[15][2];
    ele[0][2] != ele[16][2];
    ele[0][2] != ele[17][2];
    ele[0][2] != ele[18][2];
    ele[0][2] != ele[19][2];
    ele[0][2] != ele[2][0];
    ele[0][2] != ele[2][1];
    ele[0][2] != ele[2][2];
    ele[0][2] != ele[2][3];
    ele[0][2] != ele[2][4];
    ele[0][2] != ele[2][5];
    ele[0][2] != ele[20][2];
    ele[0][2] != ele[21][2];
    ele[0][2] != ele[22][2];
    ele[0][2] != ele[23][2];
    ele[0][2] != ele[24][2];
    ele[0][2] != ele[25][2];
    ele[0][2] != ele[26][2];
    ele[0][2] != ele[27][2];
    ele[0][2] != ele[28][2];
    ele[0][2] != ele[29][2];
    ele[0][2] != ele[3][0];
    ele[0][2] != ele[3][1];
    ele[0][2] != ele[3][2];
    ele[0][2] != ele[3][3];
    ele[0][2] != ele[3][4];
    ele[0][2] != ele[3][5];
    ele[0][2] != ele[30][2];
    ele[0][2] != ele[31][2];
    ele[0][2] != ele[32][2];
    ele[0][2] != ele[33][2];
    ele[0][2] != ele[34][2];
    ele[0][2] != ele[35][2];
    ele[0][2] != ele[4][0];
    ele[0][2] != ele[4][1];
    ele[0][2] != ele[4][2];
    ele[0][2] != ele[4][3];
    ele[0][2] != ele[4][4];
    ele[0][2] != ele[4][5];
    ele[0][2] != ele[5][0];
    ele[0][2] != ele[5][1];
    ele[0][2] != ele[5][2];
    ele[0][2] != ele[5][3];
    ele[0][2] != ele[5][4];
    ele[0][2] != ele[5][5];
    ele[0][2] != ele[6][2];
    ele[0][2] != ele[7][2];
    ele[0][2] != ele[8][2];
    ele[0][2] != ele[9][2];
    ele[0][20] != ele[0][21];
    ele[0][20] != ele[0][22];
    ele[0][20] != ele[0][23];
    ele[0][20] != ele[0][24];
    ele[0][20] != ele[0][25];
    ele[0][20] != ele[0][26];
    ele[0][20] != ele[0][27];
    ele[0][20] != ele[0][28];
    ele[0][20] != ele[0][29];
    ele[0][20] != ele[0][30];
    ele[0][20] != ele[0][31];
    ele[0][20] != ele[0][32];
    ele[0][20] != ele[0][33];
    ele[0][20] != ele[0][34];
    ele[0][20] != ele[0][35];
    ele[0][20] != ele[1][18];
    ele[0][20] != ele[1][19];
    ele[0][20] != ele[1][20];
    ele[0][20] != ele[1][21];
    ele[0][20] != ele[1][22];
    ele[0][20] != ele[1][23];
    ele[0][20] != ele[10][20];
    ele[0][20] != ele[11][20];
    ele[0][20] != ele[12][20];
    ele[0][20] != ele[13][20];
    ele[0][20] != ele[14][20];
    ele[0][20] != ele[15][20];
    ele[0][20] != ele[16][20];
    ele[0][20] != ele[17][20];
    ele[0][20] != ele[18][20];
    ele[0][20] != ele[19][20];
    ele[0][20] != ele[2][18];
    ele[0][20] != ele[2][19];
    ele[0][20] != ele[2][20];
    ele[0][20] != ele[2][21];
    ele[0][20] != ele[2][22];
    ele[0][20] != ele[2][23];
    ele[0][20] != ele[20][20];
    ele[0][20] != ele[21][20];
    ele[0][20] != ele[22][20];
    ele[0][20] != ele[23][20];
    ele[0][20] != ele[24][20];
    ele[0][20] != ele[25][20];
    ele[0][20] != ele[26][20];
    ele[0][20] != ele[27][20];
    ele[0][20] != ele[28][20];
    ele[0][20] != ele[29][20];
    ele[0][20] != ele[3][18];
    ele[0][20] != ele[3][19];
    ele[0][20] != ele[3][20];
    ele[0][20] != ele[3][21];
    ele[0][20] != ele[3][22];
    ele[0][20] != ele[3][23];
    ele[0][20] != ele[30][20];
    ele[0][20] != ele[31][20];
    ele[0][20] != ele[32][20];
    ele[0][20] != ele[33][20];
    ele[0][20] != ele[34][20];
    ele[0][20] != ele[35][20];
    ele[0][20] != ele[4][18];
    ele[0][20] != ele[4][19];
    ele[0][20] != ele[4][20];
    ele[0][20] != ele[4][21];
    ele[0][20] != ele[4][22];
    ele[0][20] != ele[4][23];
    ele[0][20] != ele[5][18];
    ele[0][20] != ele[5][19];
    ele[0][20] != ele[5][20];
    ele[0][20] != ele[5][21];
    ele[0][20] != ele[5][22];
    ele[0][20] != ele[5][23];
    ele[0][20] != ele[6][20];
    ele[0][20] != ele[7][20];
    ele[0][20] != ele[8][20];
    ele[0][20] != ele[9][20];
    ele[0][21] != ele[0][22];
    ele[0][21] != ele[0][23];
    ele[0][21] != ele[0][24];
    ele[0][21] != ele[0][25];
    ele[0][21] != ele[0][26];
    ele[0][21] != ele[0][27];
    ele[0][21] != ele[0][28];
    ele[0][21] != ele[0][29];
    ele[0][21] != ele[0][30];
    ele[0][21] != ele[0][31];
    ele[0][21] != ele[0][32];
    ele[0][21] != ele[0][33];
    ele[0][21] != ele[0][34];
    ele[0][21] != ele[0][35];
    ele[0][21] != ele[1][18];
    ele[0][21] != ele[1][19];
    ele[0][21] != ele[1][20];
    ele[0][21] != ele[1][21];
    ele[0][21] != ele[1][22];
    ele[0][21] != ele[1][23];
    ele[0][21] != ele[10][21];
    ele[0][21] != ele[11][21];
    ele[0][21] != ele[12][21];
    ele[0][21] != ele[13][21];
    ele[0][21] != ele[14][21];
    ele[0][21] != ele[15][21];
    ele[0][21] != ele[16][21];
    ele[0][21] != ele[17][21];
    ele[0][21] != ele[18][21];
    ele[0][21] != ele[19][21];
    ele[0][21] != ele[2][18];
    ele[0][21] != ele[2][19];
    ele[0][21] != ele[2][20];
    ele[0][21] != ele[2][21];
    ele[0][21] != ele[2][22];
    ele[0][21] != ele[2][23];
    ele[0][21] != ele[20][21];
    ele[0][21] != ele[21][21];
    ele[0][21] != ele[22][21];
    ele[0][21] != ele[23][21];
    ele[0][21] != ele[24][21];
    ele[0][21] != ele[25][21];
    ele[0][21] != ele[26][21];
    ele[0][21] != ele[27][21];
    ele[0][21] != ele[28][21];
    ele[0][21] != ele[29][21];
    ele[0][21] != ele[3][18];
    ele[0][21] != ele[3][19];
    ele[0][21] != ele[3][20];
    ele[0][21] != ele[3][21];
    ele[0][21] != ele[3][22];
    ele[0][21] != ele[3][23];
    ele[0][21] != ele[30][21];
    ele[0][21] != ele[31][21];
    ele[0][21] != ele[32][21];
    ele[0][21] != ele[33][21];
    ele[0][21] != ele[34][21];
    ele[0][21] != ele[35][21];
    ele[0][21] != ele[4][18];
    ele[0][21] != ele[4][19];
    ele[0][21] != ele[4][20];
    ele[0][21] != ele[4][21];
    ele[0][21] != ele[4][22];
    ele[0][21] != ele[4][23];
    ele[0][21] != ele[5][18];
    ele[0][21] != ele[5][19];
    ele[0][21] != ele[5][20];
    ele[0][21] != ele[5][21];
    ele[0][21] != ele[5][22];
    ele[0][21] != ele[5][23];
    ele[0][21] != ele[6][21];
    ele[0][21] != ele[7][21];
    ele[0][21] != ele[8][21];
    ele[0][21] != ele[9][21];
    ele[0][22] != ele[0][23];
    ele[0][22] != ele[0][24];
    ele[0][22] != ele[0][25];
    ele[0][22] != ele[0][26];
    ele[0][22] != ele[0][27];
    ele[0][22] != ele[0][28];
    ele[0][22] != ele[0][29];
    ele[0][22] != ele[0][30];
    ele[0][22] != ele[0][31];
    ele[0][22] != ele[0][32];
    ele[0][22] != ele[0][33];
    ele[0][22] != ele[0][34];
    ele[0][22] != ele[0][35];
    ele[0][22] != ele[1][18];
    ele[0][22] != ele[1][19];
    ele[0][22] != ele[1][20];
    ele[0][22] != ele[1][21];
    ele[0][22] != ele[1][22];
    ele[0][22] != ele[1][23];
    ele[0][22] != ele[10][22];
    ele[0][22] != ele[11][22];
    ele[0][22] != ele[12][22];
    ele[0][22] != ele[13][22];
    ele[0][22] != ele[14][22];
    ele[0][22] != ele[15][22];
    ele[0][22] != ele[16][22];
    ele[0][22] != ele[17][22];
    ele[0][22] != ele[18][22];
    ele[0][22] != ele[19][22];
    ele[0][22] != ele[2][18];
    ele[0][22] != ele[2][19];
    ele[0][22] != ele[2][20];
    ele[0][22] != ele[2][21];
    ele[0][22] != ele[2][22];
    ele[0][22] != ele[2][23];
    ele[0][22] != ele[20][22];
    ele[0][22] != ele[21][22];
    ele[0][22] != ele[22][22];
    ele[0][22] != ele[23][22];
    ele[0][22] != ele[24][22];
    ele[0][22] != ele[25][22];
    ele[0][22] != ele[26][22];
    ele[0][22] != ele[27][22];
    ele[0][22] != ele[28][22];
    ele[0][22] != ele[29][22];
    ele[0][22] != ele[3][18];
    ele[0][22] != ele[3][19];
    ele[0][22] != ele[3][20];
    ele[0][22] != ele[3][21];
    ele[0][22] != ele[3][22];
    ele[0][22] != ele[3][23];
    ele[0][22] != ele[30][22];
    ele[0][22] != ele[31][22];
    ele[0][22] != ele[32][22];
    ele[0][22] != ele[33][22];
    ele[0][22] != ele[34][22];
    ele[0][22] != ele[35][22];
    ele[0][22] != ele[4][18];
    ele[0][22] != ele[4][19];
    ele[0][22] != ele[4][20];
    ele[0][22] != ele[4][21];
    ele[0][22] != ele[4][22];
    ele[0][22] != ele[4][23];
    ele[0][22] != ele[5][18];
    ele[0][22] != ele[5][19];
    ele[0][22] != ele[5][20];
    ele[0][22] != ele[5][21];
    ele[0][22] != ele[5][22];
    ele[0][22] != ele[5][23];
    ele[0][22] != ele[6][22];
    ele[0][22] != ele[7][22];
    ele[0][22] != ele[8][22];
    ele[0][22] != ele[9][22];
    ele[0][23] != ele[0][24];
    ele[0][23] != ele[0][25];
    ele[0][23] != ele[0][26];
    ele[0][23] != ele[0][27];
    ele[0][23] != ele[0][28];
    ele[0][23] != ele[0][29];
    ele[0][23] != ele[0][30];
    ele[0][23] != ele[0][31];
    ele[0][23] != ele[0][32];
    ele[0][23] != ele[0][33];
    ele[0][23] != ele[0][34];
    ele[0][23] != ele[0][35];
    ele[0][23] != ele[1][18];
    ele[0][23] != ele[1][19];
    ele[0][23] != ele[1][20];
    ele[0][23] != ele[1][21];
    ele[0][23] != ele[1][22];
    ele[0][23] != ele[1][23];
    ele[0][23] != ele[10][23];
    ele[0][23] != ele[11][23];
    ele[0][23] != ele[12][23];
    ele[0][23] != ele[13][23];
    ele[0][23] != ele[14][23];
    ele[0][23] != ele[15][23];
    ele[0][23] != ele[16][23];
    ele[0][23] != ele[17][23];
    ele[0][23] != ele[18][23];
    ele[0][23] != ele[19][23];
    ele[0][23] != ele[2][18];
    ele[0][23] != ele[2][19];
    ele[0][23] != ele[2][20];
    ele[0][23] != ele[2][21];
    ele[0][23] != ele[2][22];
    ele[0][23] != ele[2][23];
    ele[0][23] != ele[20][23];
    ele[0][23] != ele[21][23];
    ele[0][23] != ele[22][23];
    ele[0][23] != ele[23][23];
    ele[0][23] != ele[24][23];
    ele[0][23] != ele[25][23];
    ele[0][23] != ele[26][23];
    ele[0][23] != ele[27][23];
    ele[0][23] != ele[28][23];
    ele[0][23] != ele[29][23];
    ele[0][23] != ele[3][18];
    ele[0][23] != ele[3][19];
    ele[0][23] != ele[3][20];
    ele[0][23] != ele[3][21];
    ele[0][23] != ele[3][22];
    ele[0][23] != ele[3][23];
    ele[0][23] != ele[30][23];
    ele[0][23] != ele[31][23];
    ele[0][23] != ele[32][23];
    ele[0][23] != ele[33][23];
    ele[0][23] != ele[34][23];
    ele[0][23] != ele[35][23];
    ele[0][23] != ele[4][18];
    ele[0][23] != ele[4][19];
    ele[0][23] != ele[4][20];
    ele[0][23] != ele[4][21];
    ele[0][23] != ele[4][22];
    ele[0][23] != ele[4][23];
    ele[0][23] != ele[5][18];
    ele[0][23] != ele[5][19];
    ele[0][23] != ele[5][20];
    ele[0][23] != ele[5][21];
    ele[0][23] != ele[5][22];
    ele[0][23] != ele[5][23];
    ele[0][23] != ele[6][23];
    ele[0][23] != ele[7][23];
    ele[0][23] != ele[8][23];
    ele[0][23] != ele[9][23];
    ele[0][24] != ele[0][25];
    ele[0][24] != ele[0][26];
    ele[0][24] != ele[0][27];
    ele[0][24] != ele[0][28];
    ele[0][24] != ele[0][29];
    ele[0][24] != ele[0][30];
    ele[0][24] != ele[0][31];
    ele[0][24] != ele[0][32];
    ele[0][24] != ele[0][33];
    ele[0][24] != ele[0][34];
    ele[0][24] != ele[0][35];
    ele[0][24] != ele[1][24];
    ele[0][24] != ele[1][25];
    ele[0][24] != ele[1][26];
    ele[0][24] != ele[1][27];
    ele[0][24] != ele[1][28];
    ele[0][24] != ele[1][29];
    ele[0][24] != ele[10][24];
    ele[0][24] != ele[11][24];
    ele[0][24] != ele[12][24];
    ele[0][24] != ele[13][24];
    ele[0][24] != ele[14][24];
    ele[0][24] != ele[15][24];
    ele[0][24] != ele[16][24];
    ele[0][24] != ele[17][24];
    ele[0][24] != ele[18][24];
    ele[0][24] != ele[19][24];
    ele[0][24] != ele[2][24];
    ele[0][24] != ele[2][25];
    ele[0][24] != ele[2][26];
    ele[0][24] != ele[2][27];
    ele[0][24] != ele[2][28];
    ele[0][24] != ele[2][29];
    ele[0][24] != ele[20][24];
    ele[0][24] != ele[21][24];
    ele[0][24] != ele[22][24];
    ele[0][24] != ele[23][24];
    ele[0][24] != ele[24][24];
    ele[0][24] != ele[25][24];
    ele[0][24] != ele[26][24];
    ele[0][24] != ele[27][24];
    ele[0][24] != ele[28][24];
    ele[0][24] != ele[29][24];
    ele[0][24] != ele[3][24];
    ele[0][24] != ele[3][25];
    ele[0][24] != ele[3][26];
    ele[0][24] != ele[3][27];
    ele[0][24] != ele[3][28];
    ele[0][24] != ele[3][29];
    ele[0][24] != ele[30][24];
    ele[0][24] != ele[31][24];
    ele[0][24] != ele[32][24];
    ele[0][24] != ele[33][24];
    ele[0][24] != ele[34][24];
    ele[0][24] != ele[35][24];
    ele[0][24] != ele[4][24];
    ele[0][24] != ele[4][25];
    ele[0][24] != ele[4][26];
    ele[0][24] != ele[4][27];
    ele[0][24] != ele[4][28];
    ele[0][24] != ele[4][29];
    ele[0][24] != ele[5][24];
    ele[0][24] != ele[5][25];
    ele[0][24] != ele[5][26];
    ele[0][24] != ele[5][27];
    ele[0][24] != ele[5][28];
    ele[0][24] != ele[5][29];
    ele[0][24] != ele[6][24];
    ele[0][24] != ele[7][24];
    ele[0][24] != ele[8][24];
    ele[0][24] != ele[9][24];
    ele[0][25] != ele[0][26];
    ele[0][25] != ele[0][27];
    ele[0][25] != ele[0][28];
    ele[0][25] != ele[0][29];
    ele[0][25] != ele[0][30];
    ele[0][25] != ele[0][31];
    ele[0][25] != ele[0][32];
    ele[0][25] != ele[0][33];
    ele[0][25] != ele[0][34];
    ele[0][25] != ele[0][35];
    ele[0][25] != ele[1][24];
    ele[0][25] != ele[1][25];
    ele[0][25] != ele[1][26];
    ele[0][25] != ele[1][27];
    ele[0][25] != ele[1][28];
    ele[0][25] != ele[1][29];
    ele[0][25] != ele[10][25];
    ele[0][25] != ele[11][25];
    ele[0][25] != ele[12][25];
    ele[0][25] != ele[13][25];
    ele[0][25] != ele[14][25];
    ele[0][25] != ele[15][25];
    ele[0][25] != ele[16][25];
    ele[0][25] != ele[17][25];
    ele[0][25] != ele[18][25];
    ele[0][25] != ele[19][25];
    ele[0][25] != ele[2][24];
    ele[0][25] != ele[2][25];
    ele[0][25] != ele[2][26];
    ele[0][25] != ele[2][27];
    ele[0][25] != ele[2][28];
    ele[0][25] != ele[2][29];
    ele[0][25] != ele[20][25];
    ele[0][25] != ele[21][25];
    ele[0][25] != ele[22][25];
    ele[0][25] != ele[23][25];
    ele[0][25] != ele[24][25];
    ele[0][25] != ele[25][25];
    ele[0][25] != ele[26][25];
    ele[0][25] != ele[27][25];
    ele[0][25] != ele[28][25];
    ele[0][25] != ele[29][25];
    ele[0][25] != ele[3][24];
    ele[0][25] != ele[3][25];
    ele[0][25] != ele[3][26];
    ele[0][25] != ele[3][27];
    ele[0][25] != ele[3][28];
    ele[0][25] != ele[3][29];
    ele[0][25] != ele[30][25];
    ele[0][25] != ele[31][25];
    ele[0][25] != ele[32][25];
    ele[0][25] != ele[33][25];
    ele[0][25] != ele[34][25];
    ele[0][25] != ele[35][25];
    ele[0][25] != ele[4][24];
    ele[0][25] != ele[4][25];
    ele[0][25] != ele[4][26];
    ele[0][25] != ele[4][27];
    ele[0][25] != ele[4][28];
    ele[0][25] != ele[4][29];
    ele[0][25] != ele[5][24];
    ele[0][25] != ele[5][25];
    ele[0][25] != ele[5][26];
    ele[0][25] != ele[5][27];
    ele[0][25] != ele[5][28];
    ele[0][25] != ele[5][29];
    ele[0][25] != ele[6][25];
    ele[0][25] != ele[7][25];
    ele[0][25] != ele[8][25];
    ele[0][25] != ele[9][25];
    ele[0][26] != ele[0][27];
    ele[0][26] != ele[0][28];
    ele[0][26] != ele[0][29];
    ele[0][26] != ele[0][30];
    ele[0][26] != ele[0][31];
    ele[0][26] != ele[0][32];
    ele[0][26] != ele[0][33];
    ele[0][26] != ele[0][34];
    ele[0][26] != ele[0][35];
    ele[0][26] != ele[1][24];
    ele[0][26] != ele[1][25];
    ele[0][26] != ele[1][26];
    ele[0][26] != ele[1][27];
    ele[0][26] != ele[1][28];
    ele[0][26] != ele[1][29];
    ele[0][26] != ele[10][26];
    ele[0][26] != ele[11][26];
    ele[0][26] != ele[12][26];
    ele[0][26] != ele[13][26];
    ele[0][26] != ele[14][26];
    ele[0][26] != ele[15][26];
    ele[0][26] != ele[16][26];
    ele[0][26] != ele[17][26];
    ele[0][26] != ele[18][26];
    ele[0][26] != ele[19][26];
    ele[0][26] != ele[2][24];
    ele[0][26] != ele[2][25];
    ele[0][26] != ele[2][26];
    ele[0][26] != ele[2][27];
    ele[0][26] != ele[2][28];
    ele[0][26] != ele[2][29];
    ele[0][26] != ele[20][26];
    ele[0][26] != ele[21][26];
    ele[0][26] != ele[22][26];
    ele[0][26] != ele[23][26];
    ele[0][26] != ele[24][26];
    ele[0][26] != ele[25][26];
    ele[0][26] != ele[26][26];
    ele[0][26] != ele[27][26];
    ele[0][26] != ele[28][26];
    ele[0][26] != ele[29][26];
    ele[0][26] != ele[3][24];
    ele[0][26] != ele[3][25];
    ele[0][26] != ele[3][26];
    ele[0][26] != ele[3][27];
    ele[0][26] != ele[3][28];
    ele[0][26] != ele[3][29];
    ele[0][26] != ele[30][26];
    ele[0][26] != ele[31][26];
    ele[0][26] != ele[32][26];
    ele[0][26] != ele[33][26];
    ele[0][26] != ele[34][26];
    ele[0][26] != ele[35][26];
    ele[0][26] != ele[4][24];
    ele[0][26] != ele[4][25];
    ele[0][26] != ele[4][26];
    ele[0][26] != ele[4][27];
    ele[0][26] != ele[4][28];
    ele[0][26] != ele[4][29];
    ele[0][26] != ele[5][24];
    ele[0][26] != ele[5][25];
    ele[0][26] != ele[5][26];
    ele[0][26] != ele[5][27];
    ele[0][26] != ele[5][28];
    ele[0][26] != ele[5][29];
    ele[0][26] != ele[6][26];
    ele[0][26] != ele[7][26];
    ele[0][26] != ele[8][26];
    ele[0][26] != ele[9][26];
    ele[0][27] != ele[0][28];
    ele[0][27] != ele[0][29];
    ele[0][27] != ele[0][30];
    ele[0][27] != ele[0][31];
    ele[0][27] != ele[0][32];
    ele[0][27] != ele[0][33];
    ele[0][27] != ele[0][34];
    ele[0][27] != ele[0][35];
    ele[0][27] != ele[1][24];
    ele[0][27] != ele[1][25];
    ele[0][27] != ele[1][26];
    ele[0][27] != ele[1][27];
    ele[0][27] != ele[1][28];
    ele[0][27] != ele[1][29];
    ele[0][27] != ele[10][27];
    ele[0][27] != ele[11][27];
    ele[0][27] != ele[12][27];
    ele[0][27] != ele[13][27];
    ele[0][27] != ele[14][27];
    ele[0][27] != ele[15][27];
    ele[0][27] != ele[16][27];
    ele[0][27] != ele[17][27];
    ele[0][27] != ele[18][27];
    ele[0][27] != ele[19][27];
    ele[0][27] != ele[2][24];
    ele[0][27] != ele[2][25];
    ele[0][27] != ele[2][26];
    ele[0][27] != ele[2][27];
    ele[0][27] != ele[2][28];
    ele[0][27] != ele[2][29];
    ele[0][27] != ele[20][27];
    ele[0][27] != ele[21][27];
    ele[0][27] != ele[22][27];
    ele[0][27] != ele[23][27];
    ele[0][27] != ele[24][27];
    ele[0][27] != ele[25][27];
    ele[0][27] != ele[26][27];
    ele[0][27] != ele[27][27];
    ele[0][27] != ele[28][27];
    ele[0][27] != ele[29][27];
    ele[0][27] != ele[3][24];
    ele[0][27] != ele[3][25];
    ele[0][27] != ele[3][26];
    ele[0][27] != ele[3][27];
    ele[0][27] != ele[3][28];
    ele[0][27] != ele[3][29];
    ele[0][27] != ele[30][27];
    ele[0][27] != ele[31][27];
    ele[0][27] != ele[32][27];
    ele[0][27] != ele[33][27];
    ele[0][27] != ele[34][27];
    ele[0][27] != ele[35][27];
    ele[0][27] != ele[4][24];
    ele[0][27] != ele[4][25];
    ele[0][27] != ele[4][26];
    ele[0][27] != ele[4][27];
    ele[0][27] != ele[4][28];
    ele[0][27] != ele[4][29];
    ele[0][27] != ele[5][24];
    ele[0][27] != ele[5][25];
    ele[0][27] != ele[5][26];
    ele[0][27] != ele[5][27];
    ele[0][27] != ele[5][28];
    ele[0][27] != ele[5][29];
    ele[0][27] != ele[6][27];
    ele[0][27] != ele[7][27];
    ele[0][27] != ele[8][27];
    ele[0][27] != ele[9][27];
    ele[0][28] != ele[0][29];
    ele[0][28] != ele[0][30];
    ele[0][28] != ele[0][31];
    ele[0][28] != ele[0][32];
    ele[0][28] != ele[0][33];
    ele[0][28] != ele[0][34];
    ele[0][28] != ele[0][35];
    ele[0][28] != ele[1][24];
    ele[0][28] != ele[1][25];
    ele[0][28] != ele[1][26];
    ele[0][28] != ele[1][27];
    ele[0][28] != ele[1][28];
    ele[0][28] != ele[1][29];
    ele[0][28] != ele[10][28];
    ele[0][28] != ele[11][28];
    ele[0][28] != ele[12][28];
    ele[0][28] != ele[13][28];
    ele[0][28] != ele[14][28];
    ele[0][28] != ele[15][28];
    ele[0][28] != ele[16][28];
    ele[0][28] != ele[17][28];
    ele[0][28] != ele[18][28];
    ele[0][28] != ele[19][28];
    ele[0][28] != ele[2][24];
    ele[0][28] != ele[2][25];
    ele[0][28] != ele[2][26];
    ele[0][28] != ele[2][27];
    ele[0][28] != ele[2][28];
    ele[0][28] != ele[2][29];
    ele[0][28] != ele[20][28];
    ele[0][28] != ele[21][28];
    ele[0][28] != ele[22][28];
    ele[0][28] != ele[23][28];
    ele[0][28] != ele[24][28];
    ele[0][28] != ele[25][28];
    ele[0][28] != ele[26][28];
    ele[0][28] != ele[27][28];
    ele[0][28] != ele[28][28];
    ele[0][28] != ele[29][28];
    ele[0][28] != ele[3][24];
    ele[0][28] != ele[3][25];
    ele[0][28] != ele[3][26];
    ele[0][28] != ele[3][27];
    ele[0][28] != ele[3][28];
    ele[0][28] != ele[3][29];
    ele[0][28] != ele[30][28];
    ele[0][28] != ele[31][28];
    ele[0][28] != ele[32][28];
    ele[0][28] != ele[33][28];
    ele[0][28] != ele[34][28];
    ele[0][28] != ele[35][28];
    ele[0][28] != ele[4][24];
    ele[0][28] != ele[4][25];
    ele[0][28] != ele[4][26];
    ele[0][28] != ele[4][27];
    ele[0][28] != ele[4][28];
    ele[0][28] != ele[4][29];
    ele[0][28] != ele[5][24];
    ele[0][28] != ele[5][25];
    ele[0][28] != ele[5][26];
    ele[0][28] != ele[5][27];
    ele[0][28] != ele[5][28];
    ele[0][28] != ele[5][29];
    ele[0][28] != ele[6][28];
    ele[0][28] != ele[7][28];
    ele[0][28] != ele[8][28];
    ele[0][28] != ele[9][28];
    ele[0][29] != ele[0][30];
    ele[0][29] != ele[0][31];
    ele[0][29] != ele[0][32];
    ele[0][29] != ele[0][33];
    ele[0][29] != ele[0][34];
    ele[0][29] != ele[0][35];
    ele[0][29] != ele[1][24];
    ele[0][29] != ele[1][25];
    ele[0][29] != ele[1][26];
    ele[0][29] != ele[1][27];
    ele[0][29] != ele[1][28];
    ele[0][29] != ele[1][29];
    ele[0][29] != ele[10][29];
    ele[0][29] != ele[11][29];
    ele[0][29] != ele[12][29];
    ele[0][29] != ele[13][29];
    ele[0][29] != ele[14][29];
    ele[0][29] != ele[15][29];
    ele[0][29] != ele[16][29];
    ele[0][29] != ele[17][29];
    ele[0][29] != ele[18][29];
    ele[0][29] != ele[19][29];
    ele[0][29] != ele[2][24];
    ele[0][29] != ele[2][25];
    ele[0][29] != ele[2][26];
    ele[0][29] != ele[2][27];
    ele[0][29] != ele[2][28];
    ele[0][29] != ele[2][29];
    ele[0][29] != ele[20][29];
    ele[0][29] != ele[21][29];
    ele[0][29] != ele[22][29];
    ele[0][29] != ele[23][29];
    ele[0][29] != ele[24][29];
    ele[0][29] != ele[25][29];
    ele[0][29] != ele[26][29];
    ele[0][29] != ele[27][29];
    ele[0][29] != ele[28][29];
    ele[0][29] != ele[29][29];
    ele[0][29] != ele[3][24];
    ele[0][29] != ele[3][25];
    ele[0][29] != ele[3][26];
    ele[0][29] != ele[3][27];
    ele[0][29] != ele[3][28];
    ele[0][29] != ele[3][29];
    ele[0][29] != ele[30][29];
    ele[0][29] != ele[31][29];
    ele[0][29] != ele[32][29];
    ele[0][29] != ele[33][29];
    ele[0][29] != ele[34][29];
    ele[0][29] != ele[35][29];
    ele[0][29] != ele[4][24];
    ele[0][29] != ele[4][25];
    ele[0][29] != ele[4][26];
    ele[0][29] != ele[4][27];
    ele[0][29] != ele[4][28];
    ele[0][29] != ele[4][29];
    ele[0][29] != ele[5][24];
    ele[0][29] != ele[5][25];
    ele[0][29] != ele[5][26];
    ele[0][29] != ele[5][27];
    ele[0][29] != ele[5][28];
    ele[0][29] != ele[5][29];
    ele[0][29] != ele[6][29];
    ele[0][29] != ele[7][29];
    ele[0][29] != ele[8][29];
    ele[0][29] != ele[9][29];
    ele[0][3] != ele[0][10];
    ele[0][3] != ele[0][11];
    ele[0][3] != ele[0][12];
    ele[0][3] != ele[0][13];
    ele[0][3] != ele[0][14];
    ele[0][3] != ele[0][15];
    ele[0][3] != ele[0][16];
    ele[0][3] != ele[0][17];
    ele[0][3] != ele[0][18];
    ele[0][3] != ele[0][19];
    ele[0][3] != ele[0][20];
    ele[0][3] != ele[0][21];
    ele[0][3] != ele[0][22];
    ele[0][3] != ele[0][23];
    ele[0][3] != ele[0][24];
    ele[0][3] != ele[0][25];
    ele[0][3] != ele[0][26];
    ele[0][3] != ele[0][27];
    ele[0][3] != ele[0][28];
    ele[0][3] != ele[0][29];
    ele[0][3] != ele[0][30];
    ele[0][3] != ele[0][31];
    ele[0][3] != ele[0][32];
    ele[0][3] != ele[0][33];
    ele[0][3] != ele[0][34];
    ele[0][3] != ele[0][35];
    ele[0][3] != ele[0][4];
    ele[0][3] != ele[0][5];
    ele[0][3] != ele[0][6];
    ele[0][3] != ele[0][7];
    ele[0][3] != ele[0][8];
    ele[0][3] != ele[0][9];
    ele[0][3] != ele[1][0];
    ele[0][3] != ele[1][1];
    ele[0][3] != ele[1][2];
    ele[0][3] != ele[1][3];
    ele[0][3] != ele[1][4];
    ele[0][3] != ele[1][5];
    ele[0][3] != ele[10][3];
    ele[0][3] != ele[11][3];
    ele[0][3] != ele[12][3];
    ele[0][3] != ele[13][3];
    ele[0][3] != ele[14][3];
    ele[0][3] != ele[15][3];
    ele[0][3] != ele[16][3];
    ele[0][3] != ele[17][3];
    ele[0][3] != ele[18][3];
    ele[0][3] != ele[19][3];
    ele[0][3] != ele[2][0];
    ele[0][3] != ele[2][1];
    ele[0][3] != ele[2][2];
    ele[0][3] != ele[2][3];
    ele[0][3] != ele[2][4];
    ele[0][3] != ele[2][5];
    ele[0][3] != ele[20][3];
    ele[0][3] != ele[21][3];
    ele[0][3] != ele[22][3];
    ele[0][3] != ele[23][3];
    ele[0][3] != ele[24][3];
    ele[0][3] != ele[25][3];
    ele[0][3] != ele[26][3];
    ele[0][3] != ele[27][3];
    ele[0][3] != ele[28][3];
    ele[0][3] != ele[29][3];
    ele[0][3] != ele[3][0];
    ele[0][3] != ele[3][1];
    ele[0][3] != ele[3][2];
    ele[0][3] != ele[3][3];
    ele[0][3] != ele[3][4];
    ele[0][3] != ele[3][5];
    ele[0][3] != ele[30][3];
    ele[0][3] != ele[31][3];
    ele[0][3] != ele[32][3];
    ele[0][3] != ele[33][3];
    ele[0][3] != ele[34][3];
    ele[0][3] != ele[35][3];
    ele[0][3] != ele[4][0];
    ele[0][3] != ele[4][1];
    ele[0][3] != ele[4][2];
    ele[0][3] != ele[4][3];
    ele[0][3] != ele[4][4];
    ele[0][3] != ele[4][5];
    ele[0][3] != ele[5][0];
    ele[0][3] != ele[5][1];
    ele[0][3] != ele[5][2];
    ele[0][3] != ele[5][3];
    ele[0][3] != ele[5][4];
    ele[0][3] != ele[5][5];
    ele[0][3] != ele[6][3];
    ele[0][3] != ele[7][3];
    ele[0][3] != ele[8][3];
    ele[0][3] != ele[9][3];
    ele[0][30] != ele[0][31];
    ele[0][30] != ele[0][32];
    ele[0][30] != ele[0][33];
    ele[0][30] != ele[0][34];
    ele[0][30] != ele[0][35];
    ele[0][30] != ele[1][30];
    ele[0][30] != ele[1][31];
    ele[0][30] != ele[1][32];
    ele[0][30] != ele[1][33];
    ele[0][30] != ele[1][34];
    ele[0][30] != ele[1][35];
    ele[0][30] != ele[10][30];
    ele[0][30] != ele[11][30];
    ele[0][30] != ele[12][30];
    ele[0][30] != ele[13][30];
    ele[0][30] != ele[14][30];
    ele[0][30] != ele[15][30];
    ele[0][30] != ele[16][30];
    ele[0][30] != ele[17][30];
    ele[0][30] != ele[18][30];
    ele[0][30] != ele[19][30];
    ele[0][30] != ele[2][30];
    ele[0][30] != ele[2][31];
    ele[0][30] != ele[2][32];
    ele[0][30] != ele[2][33];
    ele[0][30] != ele[2][34];
    ele[0][30] != ele[2][35];
    ele[0][30] != ele[20][30];
    ele[0][30] != ele[21][30];
    ele[0][30] != ele[22][30];
    ele[0][30] != ele[23][30];
    ele[0][30] != ele[24][30];
    ele[0][30] != ele[25][30];
    ele[0][30] != ele[26][30];
    ele[0][30] != ele[27][30];
    ele[0][30] != ele[28][30];
    ele[0][30] != ele[29][30];
    ele[0][30] != ele[3][30];
    ele[0][30] != ele[3][31];
    ele[0][30] != ele[3][32];
    ele[0][30] != ele[3][33];
    ele[0][30] != ele[3][34];
    ele[0][30] != ele[3][35];
    ele[0][30] != ele[30][30];
    ele[0][30] != ele[31][30];
    ele[0][30] != ele[32][30];
    ele[0][30] != ele[33][30];
    ele[0][30] != ele[34][30];
    ele[0][30] != ele[35][30];
    ele[0][30] != ele[4][30];
    ele[0][30] != ele[4][31];
    ele[0][30] != ele[4][32];
    ele[0][30] != ele[4][33];
    ele[0][30] != ele[4][34];
    ele[0][30] != ele[4][35];
    ele[0][30] != ele[5][30];
    ele[0][30] != ele[5][31];
    ele[0][30] != ele[5][32];
    ele[0][30] != ele[5][33];
    ele[0][30] != ele[5][34];
    ele[0][30] != ele[5][35];
    ele[0][30] != ele[6][30];
    ele[0][30] != ele[7][30];
    ele[0][30] != ele[8][30];
    ele[0][30] != ele[9][30];
    ele[0][31] != ele[0][32];
    ele[0][31] != ele[0][33];
    ele[0][31] != ele[0][34];
    ele[0][31] != ele[0][35];
    ele[0][31] != ele[1][30];
    ele[0][31] != ele[1][31];
    ele[0][31] != ele[1][32];
    ele[0][31] != ele[1][33];
    ele[0][31] != ele[1][34];
    ele[0][31] != ele[1][35];
    ele[0][31] != ele[10][31];
    ele[0][31] != ele[11][31];
    ele[0][31] != ele[12][31];
    ele[0][31] != ele[13][31];
    ele[0][31] != ele[14][31];
    ele[0][31] != ele[15][31];
    ele[0][31] != ele[16][31];
    ele[0][31] != ele[17][31];
    ele[0][31] != ele[18][31];
    ele[0][31] != ele[19][31];
    ele[0][31] != ele[2][30];
    ele[0][31] != ele[2][31];
    ele[0][31] != ele[2][32];
    ele[0][31] != ele[2][33];
    ele[0][31] != ele[2][34];
    ele[0][31] != ele[2][35];
    ele[0][31] != ele[20][31];
    ele[0][31] != ele[21][31];
    ele[0][31] != ele[22][31];
    ele[0][31] != ele[23][31];
    ele[0][31] != ele[24][31];
    ele[0][31] != ele[25][31];
    ele[0][31] != ele[26][31];
    ele[0][31] != ele[27][31];
    ele[0][31] != ele[28][31];
    ele[0][31] != ele[29][31];
    ele[0][31] != ele[3][30];
    ele[0][31] != ele[3][31];
    ele[0][31] != ele[3][32];
    ele[0][31] != ele[3][33];
    ele[0][31] != ele[3][34];
    ele[0][31] != ele[3][35];
    ele[0][31] != ele[30][31];
    ele[0][31] != ele[31][31];
    ele[0][31] != ele[32][31];
    ele[0][31] != ele[33][31];
    ele[0][31] != ele[34][31];
    ele[0][31] != ele[35][31];
    ele[0][31] != ele[4][30];
    ele[0][31] != ele[4][31];
    ele[0][31] != ele[4][32];
    ele[0][31] != ele[4][33];
    ele[0][31] != ele[4][34];
    ele[0][31] != ele[4][35];
    ele[0][31] != ele[5][30];
    ele[0][31] != ele[5][31];
    ele[0][31] != ele[5][32];
    ele[0][31] != ele[5][33];
    ele[0][31] != ele[5][34];
    ele[0][31] != ele[5][35];
    ele[0][31] != ele[6][31];
    ele[0][31] != ele[7][31];
    ele[0][31] != ele[8][31];
    ele[0][31] != ele[9][31];
    ele[0][32] != ele[0][33];
    ele[0][32] != ele[0][34];
    ele[0][32] != ele[0][35];
    ele[0][32] != ele[1][30];
    ele[0][32] != ele[1][31];
    ele[0][32] != ele[1][32];
    ele[0][32] != ele[1][33];
    ele[0][32] != ele[1][34];
    ele[0][32] != ele[1][35];
    ele[0][32] != ele[10][32];
    ele[0][32] != ele[11][32];
    ele[0][32] != ele[12][32];
    ele[0][32] != ele[13][32];
    ele[0][32] != ele[14][32];
    ele[0][32] != ele[15][32];
    ele[0][32] != ele[16][32];
    ele[0][32] != ele[17][32];
    ele[0][32] != ele[18][32];
    ele[0][32] != ele[19][32];
    ele[0][32] != ele[2][30];
    ele[0][32] != ele[2][31];
    ele[0][32] != ele[2][32];
    ele[0][32] != ele[2][33];
    ele[0][32] != ele[2][34];
    ele[0][32] != ele[2][35];
    ele[0][32] != ele[20][32];
    ele[0][32] != ele[21][32];
    ele[0][32] != ele[22][32];
    ele[0][32] != ele[23][32];
    ele[0][32] != ele[24][32];
    ele[0][32] != ele[25][32];
    ele[0][32] != ele[26][32];
    ele[0][32] != ele[27][32];
    ele[0][32] != ele[28][32];
    ele[0][32] != ele[29][32];
    ele[0][32] != ele[3][30];
    ele[0][32] != ele[3][31];
    ele[0][32] != ele[3][32];
    ele[0][32] != ele[3][33];
    ele[0][32] != ele[3][34];
    ele[0][32] != ele[3][35];
    ele[0][32] != ele[30][32];
    ele[0][32] != ele[31][32];
    ele[0][32] != ele[32][32];
    ele[0][32] != ele[33][32];
    ele[0][32] != ele[34][32];
    ele[0][32] != ele[35][32];
    ele[0][32] != ele[4][30];
    ele[0][32] != ele[4][31];
    ele[0][32] != ele[4][32];
    ele[0][32] != ele[4][33];
    ele[0][32] != ele[4][34];
    ele[0][32] != ele[4][35];
    ele[0][32] != ele[5][30];
    ele[0][32] != ele[5][31];
    ele[0][32] != ele[5][32];
    ele[0][32] != ele[5][33];
    ele[0][32] != ele[5][34];
    ele[0][32] != ele[5][35];
    ele[0][32] != ele[6][32];
    ele[0][32] != ele[7][32];
    ele[0][32] != ele[8][32];
    ele[0][32] != ele[9][32];
    ele[0][33] != ele[0][34];
    ele[0][33] != ele[0][35];
    ele[0][33] != ele[1][30];
    ele[0][33] != ele[1][31];
    ele[0][33] != ele[1][32];
    ele[0][33] != ele[1][33];
    ele[0][33] != ele[1][34];
    ele[0][33] != ele[1][35];
    ele[0][33] != ele[10][33];
    ele[0][33] != ele[11][33];
    ele[0][33] != ele[12][33];
    ele[0][33] != ele[13][33];
    ele[0][33] != ele[14][33];
    ele[0][33] != ele[15][33];
    ele[0][33] != ele[16][33];
    ele[0][33] != ele[17][33];
    ele[0][33] != ele[18][33];
    ele[0][33] != ele[19][33];
    ele[0][33] != ele[2][30];
    ele[0][33] != ele[2][31];
    ele[0][33] != ele[2][32];
    ele[0][33] != ele[2][33];
    ele[0][33] != ele[2][34];
    ele[0][33] != ele[2][35];
    ele[0][33] != ele[20][33];
    ele[0][33] != ele[21][33];
    ele[0][33] != ele[22][33];
    ele[0][33] != ele[23][33];
    ele[0][33] != ele[24][33];
    ele[0][33] != ele[25][33];
    ele[0][33] != ele[26][33];
    ele[0][33] != ele[27][33];
    ele[0][33] != ele[28][33];
    ele[0][33] != ele[29][33];
    ele[0][33] != ele[3][30];
    ele[0][33] != ele[3][31];
    ele[0][33] != ele[3][32];
    ele[0][33] != ele[3][33];
    ele[0][33] != ele[3][34];
    ele[0][33] != ele[3][35];
    ele[0][33] != ele[30][33];
    ele[0][33] != ele[31][33];
    ele[0][33] != ele[32][33];
    ele[0][33] != ele[33][33];
    ele[0][33] != ele[34][33];
    ele[0][33] != ele[35][33];
    ele[0][33] != ele[4][30];
    ele[0][33] != ele[4][31];
    ele[0][33] != ele[4][32];
    ele[0][33] != ele[4][33];
    ele[0][33] != ele[4][34];
    ele[0][33] != ele[4][35];
    ele[0][33] != ele[5][30];
    ele[0][33] != ele[5][31];
    ele[0][33] != ele[5][32];
    ele[0][33] != ele[5][33];
    ele[0][33] != ele[5][34];
    ele[0][33] != ele[5][35];
    ele[0][33] != ele[6][33];
    ele[0][33] != ele[7][33];
    ele[0][33] != ele[8][33];
    ele[0][33] != ele[9][33];
    ele[0][34] != ele[0][35];
    ele[0][34] != ele[1][30];
    ele[0][34] != ele[1][31];
    ele[0][34] != ele[1][32];
    ele[0][34] != ele[1][33];
    ele[0][34] != ele[1][34];
    ele[0][34] != ele[1][35];
    ele[0][34] != ele[10][34];
    ele[0][34] != ele[11][34];
    ele[0][34] != ele[12][34];
    ele[0][34] != ele[13][34];
    ele[0][34] != ele[14][34];
    ele[0][34] != ele[15][34];
    ele[0][34] != ele[16][34];
    ele[0][34] != ele[17][34];
    ele[0][34] != ele[18][34];
    ele[0][34] != ele[19][34];
    ele[0][34] != ele[2][30];
    ele[0][34] != ele[2][31];
    ele[0][34] != ele[2][32];
    ele[0][34] != ele[2][33];
    ele[0][34] != ele[2][34];
    ele[0][34] != ele[2][35];
    ele[0][34] != ele[20][34];
    ele[0][34] != ele[21][34];
    ele[0][34] != ele[22][34];
    ele[0][34] != ele[23][34];
    ele[0][34] != ele[24][34];
    ele[0][34] != ele[25][34];
    ele[0][34] != ele[26][34];
    ele[0][34] != ele[27][34];
    ele[0][34] != ele[28][34];
    ele[0][34] != ele[29][34];
    ele[0][34] != ele[3][30];
    ele[0][34] != ele[3][31];
    ele[0][34] != ele[3][32];
    ele[0][34] != ele[3][33];
    ele[0][34] != ele[3][34];
    ele[0][34] != ele[3][35];
    ele[0][34] != ele[30][34];
    ele[0][34] != ele[31][34];
    ele[0][34] != ele[32][34];
    ele[0][34] != ele[33][34];
    ele[0][34] != ele[34][34];
    ele[0][34] != ele[35][34];
    ele[0][34] != ele[4][30];
    ele[0][34] != ele[4][31];
    ele[0][34] != ele[4][32];
    ele[0][34] != ele[4][33];
    ele[0][34] != ele[4][34];
    ele[0][34] != ele[4][35];
    ele[0][34] != ele[5][30];
    ele[0][34] != ele[5][31];
    ele[0][34] != ele[5][32];
    ele[0][34] != ele[5][33];
    ele[0][34] != ele[5][34];
    ele[0][34] != ele[5][35];
    ele[0][34] != ele[6][34];
    ele[0][34] != ele[7][34];
    ele[0][34] != ele[8][34];
    ele[0][34] != ele[9][34];
    ele[0][35] != ele[1][30];
    ele[0][35] != ele[1][31];
    ele[0][35] != ele[1][32];
    ele[0][35] != ele[1][33];
    ele[0][35] != ele[1][34];
    ele[0][35] != ele[1][35];
    ele[0][35] != ele[10][35];
    ele[0][35] != ele[11][35];
    ele[0][35] != ele[12][35];
    ele[0][35] != ele[13][35];
    ele[0][35] != ele[14][35];
    ele[0][35] != ele[15][35];
    ele[0][35] != ele[16][35];
    ele[0][35] != ele[17][35];
    ele[0][35] != ele[18][35];
    ele[0][35] != ele[19][35];
    ele[0][35] != ele[2][30];
    ele[0][35] != ele[2][31];
    ele[0][35] != ele[2][32];
    ele[0][35] != ele[2][33];
    ele[0][35] != ele[2][34];
    ele[0][35] != ele[2][35];
    ele[0][35] != ele[20][35];
    ele[0][35] != ele[21][35];
    ele[0][35] != ele[22][35];
    ele[0][35] != ele[23][35];
    ele[0][35] != ele[24][35];
    ele[0][35] != ele[25][35];
    ele[0][35] != ele[26][35];
    ele[0][35] != ele[27][35];
    ele[0][35] != ele[28][35];
    ele[0][35] != ele[29][35];
    ele[0][35] != ele[3][30];
    ele[0][35] != ele[3][31];
    ele[0][35] != ele[3][32];
    ele[0][35] != ele[3][33];
    ele[0][35] != ele[3][34];
    ele[0][35] != ele[3][35];
    ele[0][35] != ele[30][35];
    ele[0][35] != ele[31][35];
    ele[0][35] != ele[32][35];
    ele[0][35] != ele[33][35];
    ele[0][35] != ele[34][35];
    ele[0][35] != ele[35][35];
    ele[0][35] != ele[4][30];
    ele[0][35] != ele[4][31];
    ele[0][35] != ele[4][32];
    ele[0][35] != ele[4][33];
    ele[0][35] != ele[4][34];
    ele[0][35] != ele[4][35];
    ele[0][35] != ele[5][30];
    ele[0][35] != ele[5][31];
    ele[0][35] != ele[5][32];
    ele[0][35] != ele[5][33];
    ele[0][35] != ele[5][34];
    ele[0][35] != ele[5][35];
    ele[0][35] != ele[6][35];
    ele[0][35] != ele[7][35];
    ele[0][35] != ele[8][35];
    ele[0][35] != ele[9][35];
    ele[0][4] != ele[0][10];
    ele[0][4] != ele[0][11];
    ele[0][4] != ele[0][12];
    ele[0][4] != ele[0][13];
    ele[0][4] != ele[0][14];
    ele[0][4] != ele[0][15];
    ele[0][4] != ele[0][16];
    ele[0][4] != ele[0][17];
    ele[0][4] != ele[0][18];
    ele[0][4] != ele[0][19];
    ele[0][4] != ele[0][20];
    ele[0][4] != ele[0][21];
    ele[0][4] != ele[0][22];
    ele[0][4] != ele[0][23];
    ele[0][4] != ele[0][24];
    ele[0][4] != ele[0][25];
    ele[0][4] != ele[0][26];
    ele[0][4] != ele[0][27];
    ele[0][4] != ele[0][28];
    ele[0][4] != ele[0][29];
    ele[0][4] != ele[0][30];
    ele[0][4] != ele[0][31];
    ele[0][4] != ele[0][32];
    ele[0][4] != ele[0][33];
    ele[0][4] != ele[0][34];
    ele[0][4] != ele[0][35];
    ele[0][4] != ele[0][5];
    ele[0][4] != ele[0][6];
    ele[0][4] != ele[0][7];
    ele[0][4] != ele[0][8];
    ele[0][4] != ele[0][9];
    ele[0][4] != ele[1][0];
    ele[0][4] != ele[1][1];
    ele[0][4] != ele[1][2];
    ele[0][4] != ele[1][3];
    ele[0][4] != ele[1][4];
    ele[0][4] != ele[1][5];
    ele[0][4] != ele[10][4];
    ele[0][4] != ele[11][4];
    ele[0][4] != ele[12][4];
    ele[0][4] != ele[13][4];
    ele[0][4] != ele[14][4];
    ele[0][4] != ele[15][4];
    ele[0][4] != ele[16][4];
    ele[0][4] != ele[17][4];
    ele[0][4] != ele[18][4];
    ele[0][4] != ele[19][4];
    ele[0][4] != ele[2][0];
    ele[0][4] != ele[2][1];
    ele[0][4] != ele[2][2];
    ele[0][4] != ele[2][3];
    ele[0][4] != ele[2][4];
    ele[0][4] != ele[2][5];
    ele[0][4] != ele[20][4];
    ele[0][4] != ele[21][4];
    ele[0][4] != ele[22][4];
    ele[0][4] != ele[23][4];
    ele[0][4] != ele[24][4];
    ele[0][4] != ele[25][4];
    ele[0][4] != ele[26][4];
    ele[0][4] != ele[27][4];
    ele[0][4] != ele[28][4];
    ele[0][4] != ele[29][4];
    ele[0][4] != ele[3][0];
    ele[0][4] != ele[3][1];
    ele[0][4] != ele[3][2];
    ele[0][4] != ele[3][3];
    ele[0][4] != ele[3][4];
    ele[0][4] != ele[3][5];
    ele[0][4] != ele[30][4];
    ele[0][4] != ele[31][4];
    ele[0][4] != ele[32][4];
    ele[0][4] != ele[33][4];
    ele[0][4] != ele[34][4];
    ele[0][4] != ele[35][4];
    ele[0][4] != ele[4][0];
    ele[0][4] != ele[4][1];
    ele[0][4] != ele[4][2];
    ele[0][4] != ele[4][3];
    ele[0][4] != ele[4][4];
    ele[0][4] != ele[4][5];
    ele[0][4] != ele[5][0];
    ele[0][4] != ele[5][1];
    ele[0][4] != ele[5][2];
    ele[0][4] != ele[5][3];
    ele[0][4] != ele[5][4];
    ele[0][4] != ele[5][5];
    ele[0][4] != ele[6][4];
    ele[0][4] != ele[7][4];
    ele[0][4] != ele[8][4];
    ele[0][4] != ele[9][4];
    ele[0][5] != ele[0][10];
    ele[0][5] != ele[0][11];
    ele[0][5] != ele[0][12];
    ele[0][5] != ele[0][13];
    ele[0][5] != ele[0][14];
    ele[0][5] != ele[0][15];
    ele[0][5] != ele[0][16];
    ele[0][5] != ele[0][17];
    ele[0][5] != ele[0][18];
    ele[0][5] != ele[0][19];
    ele[0][5] != ele[0][20];
    ele[0][5] != ele[0][21];
    ele[0][5] != ele[0][22];
    ele[0][5] != ele[0][23];
    ele[0][5] != ele[0][24];
    ele[0][5] != ele[0][25];
    ele[0][5] != ele[0][26];
    ele[0][5] != ele[0][27];
    ele[0][5] != ele[0][28];
    ele[0][5] != ele[0][29];
    ele[0][5] != ele[0][30];
    ele[0][5] != ele[0][31];
    ele[0][5] != ele[0][32];
    ele[0][5] != ele[0][33];
    ele[0][5] != ele[0][34];
    ele[0][5] != ele[0][35];
    ele[0][5] != ele[0][6];
    ele[0][5] != ele[0][7];
    ele[0][5] != ele[0][8];
    ele[0][5] != ele[0][9];
    ele[0][5] != ele[1][0];
    ele[0][5] != ele[1][1];
    ele[0][5] != ele[1][2];
    ele[0][5] != ele[1][3];
    ele[0][5] != ele[1][4];
    ele[0][5] != ele[1][5];
    ele[0][5] != ele[10][5];
    ele[0][5] != ele[11][5];
    ele[0][5] != ele[12][5];
    ele[0][5] != ele[13][5];
    ele[0][5] != ele[14][5];
    ele[0][5] != ele[15][5];
    ele[0][5] != ele[16][5];
    ele[0][5] != ele[17][5];
    ele[0][5] != ele[18][5];
    ele[0][5] != ele[19][5];
    ele[0][5] != ele[2][0];
    ele[0][5] != ele[2][1];
    ele[0][5] != ele[2][2];
    ele[0][5] != ele[2][3];
    ele[0][5] != ele[2][4];
    ele[0][5] != ele[2][5];
    ele[0][5] != ele[20][5];
    ele[0][5] != ele[21][5];
    ele[0][5] != ele[22][5];
    ele[0][5] != ele[23][5];
    ele[0][5] != ele[24][5];
    ele[0][5] != ele[25][5];
    ele[0][5] != ele[26][5];
    ele[0][5] != ele[27][5];
    ele[0][5] != ele[28][5];
    ele[0][5] != ele[29][5];
    ele[0][5] != ele[3][0];
    ele[0][5] != ele[3][1];
    ele[0][5] != ele[3][2];
    ele[0][5] != ele[3][3];
    ele[0][5] != ele[3][4];
    ele[0][5] != ele[3][5];
    ele[0][5] != ele[30][5];
    ele[0][5] != ele[31][5];
    ele[0][5] != ele[32][5];
    ele[0][5] != ele[33][5];
    ele[0][5] != ele[34][5];
    ele[0][5] != ele[35][5];
    ele[0][5] != ele[4][0];
    ele[0][5] != ele[4][1];
    ele[0][5] != ele[4][2];
    ele[0][5] != ele[4][3];
    ele[0][5] != ele[4][4];
    ele[0][5] != ele[4][5];
    ele[0][5] != ele[5][0];
    ele[0][5] != ele[5][1];
    ele[0][5] != ele[5][2];
    ele[0][5] != ele[5][3];
    ele[0][5] != ele[5][4];
    ele[0][5] != ele[5][5];
    ele[0][5] != ele[6][5];
    ele[0][5] != ele[7][5];
    ele[0][5] != ele[8][5];
    ele[0][5] != ele[9][5];
    ele[0][6] != ele[0][10];
    ele[0][6] != ele[0][11];
    ele[0][6] != ele[0][12];
    ele[0][6] != ele[0][13];
    ele[0][6] != ele[0][14];
    ele[0][6] != ele[0][15];
    ele[0][6] != ele[0][16];
    ele[0][6] != ele[0][17];
    ele[0][6] != ele[0][18];
    ele[0][6] != ele[0][19];
    ele[0][6] != ele[0][20];
    ele[0][6] != ele[0][21];
    ele[0][6] != ele[0][22];
    ele[0][6] != ele[0][23];
    ele[0][6] != ele[0][24];
    ele[0][6] != ele[0][25];
    ele[0][6] != ele[0][26];
    ele[0][6] != ele[0][27];
    ele[0][6] != ele[0][28];
    ele[0][6] != ele[0][29];
    ele[0][6] != ele[0][30];
    ele[0][6] != ele[0][31];
    ele[0][6] != ele[0][32];
    ele[0][6] != ele[0][33];
    ele[0][6] != ele[0][34];
    ele[0][6] != ele[0][35];
    ele[0][6] != ele[0][7];
    ele[0][6] != ele[0][8];
    ele[0][6] != ele[0][9];
    ele[0][6] != ele[1][10];
    ele[0][6] != ele[1][11];
    ele[0][6] != ele[1][6];
    ele[0][6] != ele[1][7];
    ele[0][6] != ele[1][8];
    ele[0][6] != ele[1][9];
    ele[0][6] != ele[10][6];
    ele[0][6] != ele[11][6];
    ele[0][6] != ele[12][6];
    ele[0][6] != ele[13][6];
    ele[0][6] != ele[14][6];
    ele[0][6] != ele[15][6];
    ele[0][6] != ele[16][6];
    ele[0][6] != ele[17][6];
    ele[0][6] != ele[18][6];
    ele[0][6] != ele[19][6];
    ele[0][6] != ele[2][10];
    ele[0][6] != ele[2][11];
    ele[0][6] != ele[2][6];
    ele[0][6] != ele[2][7];
    ele[0][6] != ele[2][8];
    ele[0][6] != ele[2][9];
    ele[0][6] != ele[20][6];
    ele[0][6] != ele[21][6];
    ele[0][6] != ele[22][6];
    ele[0][6] != ele[23][6];
    ele[0][6] != ele[24][6];
    ele[0][6] != ele[25][6];
    ele[0][6] != ele[26][6];
    ele[0][6] != ele[27][6];
    ele[0][6] != ele[28][6];
    ele[0][6] != ele[29][6];
    ele[0][6] != ele[3][10];
    ele[0][6] != ele[3][11];
    ele[0][6] != ele[3][6];
    ele[0][6] != ele[3][7];
    ele[0][6] != ele[3][8];
    ele[0][6] != ele[3][9];
    ele[0][6] != ele[30][6];
    ele[0][6] != ele[31][6];
    ele[0][6] != ele[32][6];
    ele[0][6] != ele[33][6];
    ele[0][6] != ele[34][6];
    ele[0][6] != ele[35][6];
    ele[0][6] != ele[4][10];
    ele[0][6] != ele[4][11];
    ele[0][6] != ele[4][6];
    ele[0][6] != ele[4][7];
    ele[0][6] != ele[4][8];
    ele[0][6] != ele[4][9];
    ele[0][6] != ele[5][10];
    ele[0][6] != ele[5][11];
    ele[0][6] != ele[5][6];
    ele[0][6] != ele[5][7];
    ele[0][6] != ele[5][8];
    ele[0][6] != ele[5][9];
    ele[0][6] != ele[6][6];
    ele[0][6] != ele[7][6];
    ele[0][6] != ele[8][6];
    ele[0][6] != ele[9][6];
    ele[0][7] != ele[0][10];
    ele[0][7] != ele[0][11];
    ele[0][7] != ele[0][12];
    ele[0][7] != ele[0][13];
    ele[0][7] != ele[0][14];
    ele[0][7] != ele[0][15];
    ele[0][7] != ele[0][16];
    ele[0][7] != ele[0][17];
    ele[0][7] != ele[0][18];
    ele[0][7] != ele[0][19];
    ele[0][7] != ele[0][20];
    ele[0][7] != ele[0][21];
    ele[0][7] != ele[0][22];
    ele[0][7] != ele[0][23];
    ele[0][7] != ele[0][24];
    ele[0][7] != ele[0][25];
    ele[0][7] != ele[0][26];
    ele[0][7] != ele[0][27];
    ele[0][7] != ele[0][28];
    ele[0][7] != ele[0][29];
    ele[0][7] != ele[0][30];
    ele[0][7] != ele[0][31];
    ele[0][7] != ele[0][32];
    ele[0][7] != ele[0][33];
    ele[0][7] != ele[0][34];
    ele[0][7] != ele[0][35];
    ele[0][7] != ele[0][8];
    ele[0][7] != ele[0][9];
    ele[0][7] != ele[1][10];
    ele[0][7] != ele[1][11];
    ele[0][7] != ele[1][6];
    ele[0][7] != ele[1][7];
    ele[0][7] != ele[1][8];
    ele[0][7] != ele[1][9];
    ele[0][7] != ele[10][7];
    ele[0][7] != ele[11][7];
    ele[0][7] != ele[12][7];
    ele[0][7] != ele[13][7];
    ele[0][7] != ele[14][7];
    ele[0][7] != ele[15][7];
    ele[0][7] != ele[16][7];
    ele[0][7] != ele[17][7];
    ele[0][7] != ele[18][7];
    ele[0][7] != ele[19][7];
    ele[0][7] != ele[2][10];
    ele[0][7] != ele[2][11];
    ele[0][7] != ele[2][6];
    ele[0][7] != ele[2][7];
    ele[0][7] != ele[2][8];
    ele[0][7] != ele[2][9];
    ele[0][7] != ele[20][7];
    ele[0][7] != ele[21][7];
    ele[0][7] != ele[22][7];
    ele[0][7] != ele[23][7];
    ele[0][7] != ele[24][7];
    ele[0][7] != ele[25][7];
    ele[0][7] != ele[26][7];
    ele[0][7] != ele[27][7];
    ele[0][7] != ele[28][7];
    ele[0][7] != ele[29][7];
    ele[0][7] != ele[3][10];
    ele[0][7] != ele[3][11];
    ele[0][7] != ele[3][6];
    ele[0][7] != ele[3][7];
    ele[0][7] != ele[3][8];
    ele[0][7] != ele[3][9];
    ele[0][7] != ele[30][7];
    ele[0][7] != ele[31][7];
    ele[0][7] != ele[32][7];
    ele[0][7] != ele[33][7];
    ele[0][7] != ele[34][7];
    ele[0][7] != ele[35][7];
    ele[0][7] != ele[4][10];
    ele[0][7] != ele[4][11];
    ele[0][7] != ele[4][6];
    ele[0][7] != ele[4][7];
    ele[0][7] != ele[4][8];
    ele[0][7] != ele[4][9];
    ele[0][7] != ele[5][10];
    ele[0][7] != ele[5][11];
    ele[0][7] != ele[5][6];
    ele[0][7] != ele[5][7];
    ele[0][7] != ele[5][8];
    ele[0][7] != ele[5][9];
    ele[0][7] != ele[6][7];
    ele[0][7] != ele[7][7];
    ele[0][7] != ele[8][7];
    ele[0][7] != ele[9][7];
    ele[0][8] != ele[0][10];
    ele[0][8] != ele[0][11];
    ele[0][8] != ele[0][12];
    ele[0][8] != ele[0][13];
    ele[0][8] != ele[0][14];
    ele[0][8] != ele[0][15];
    ele[0][8] != ele[0][16];
    ele[0][8] != ele[0][17];
    ele[0][8] != ele[0][18];
    ele[0][8] != ele[0][19];
    ele[0][8] != ele[0][20];
    ele[0][8] != ele[0][21];
    ele[0][8] != ele[0][22];
    ele[0][8] != ele[0][23];
    ele[0][8] != ele[0][24];
    ele[0][8] != ele[0][25];
    ele[0][8] != ele[0][26];
    ele[0][8] != ele[0][27];
    ele[0][8] != ele[0][28];
    ele[0][8] != ele[0][29];
    ele[0][8] != ele[0][30];
    ele[0][8] != ele[0][31];
    ele[0][8] != ele[0][32];
    ele[0][8] != ele[0][33];
    ele[0][8] != ele[0][34];
    ele[0][8] != ele[0][35];
    ele[0][8] != ele[0][9];
    ele[0][8] != ele[1][10];
    ele[0][8] != ele[1][11];
    ele[0][8] != ele[1][6];
    ele[0][8] != ele[1][7];
    ele[0][8] != ele[1][8];
    ele[0][8] != ele[1][9];
    ele[0][8] != ele[10][8];
    ele[0][8] != ele[11][8];
    ele[0][8] != ele[12][8];
    ele[0][8] != ele[13][8];
    ele[0][8] != ele[14][8];
    ele[0][8] != ele[15][8];
    ele[0][8] != ele[16][8];
    ele[0][8] != ele[17][8];
    ele[0][8] != ele[18][8];
    ele[0][8] != ele[19][8];
    ele[0][8] != ele[2][10];
    ele[0][8] != ele[2][11];
    ele[0][8] != ele[2][6];
    ele[0][8] != ele[2][7];
    ele[0][8] != ele[2][8];
    ele[0][8] != ele[2][9];
    ele[0][8] != ele[20][8];
    ele[0][8] != ele[21][8];
    ele[0][8] != ele[22][8];
    ele[0][8] != ele[23][8];
    ele[0][8] != ele[24][8];
    ele[0][8] != ele[25][8];
    ele[0][8] != ele[26][8];
    ele[0][8] != ele[27][8];
    ele[0][8] != ele[28][8];
    ele[0][8] != ele[29][8];
    ele[0][8] != ele[3][10];
    ele[0][8] != ele[3][11];
    ele[0][8] != ele[3][6];
    ele[0][8] != ele[3][7];
    ele[0][8] != ele[3][8];
    ele[0][8] != ele[3][9];
    ele[0][8] != ele[30][8];
    ele[0][8] != ele[31][8];
    ele[0][8] != ele[32][8];
    ele[0][8] != ele[33][8];
    ele[0][8] != ele[34][8];
    ele[0][8] != ele[35][8];
    ele[0][8] != ele[4][10];
    ele[0][8] != ele[4][11];
    ele[0][8] != ele[4][6];
    ele[0][8] != ele[4][7];
    ele[0][8] != ele[4][8];
    ele[0][8] != ele[4][9];
    ele[0][8] != ele[5][10];
    ele[0][8] != ele[5][11];
    ele[0][8] != ele[5][6];
    ele[0][8] != ele[5][7];
    ele[0][8] != ele[5][8];
    ele[0][8] != ele[5][9];
    ele[0][8] != ele[6][8];
    ele[0][8] != ele[7][8];
    ele[0][8] != ele[8][8];
    ele[0][8] != ele[9][8];
    ele[0][9] != ele[0][10];
    ele[0][9] != ele[0][11];
    ele[0][9] != ele[0][12];
    ele[0][9] != ele[0][13];
    ele[0][9] != ele[0][14];
    ele[0][9] != ele[0][15];
    ele[0][9] != ele[0][16];
    ele[0][9] != ele[0][17];
    ele[0][9] != ele[0][18];
    ele[0][9] != ele[0][19];
    ele[0][9] != ele[0][20];
    ele[0][9] != ele[0][21];
    ele[0][9] != ele[0][22];
    ele[0][9] != ele[0][23];
    ele[0][9] != ele[0][24];
    ele[0][9] != ele[0][25];
    ele[0][9] != ele[0][26];
    ele[0][9] != ele[0][27];
    ele[0][9] != ele[0][28];
    ele[0][9] != ele[0][29];
    ele[0][9] != ele[0][30];
    ele[0][9] != ele[0][31];
    ele[0][9] != ele[0][32];
    ele[0][9] != ele[0][33];
    ele[0][9] != ele[0][34];
    ele[0][9] != ele[0][35];
    ele[0][9] != ele[1][10];
    ele[0][9] != ele[1][11];
    ele[0][9] != ele[1][6];
    ele[0][9] != ele[1][7];
    ele[0][9] != ele[1][8];
    ele[0][9] != ele[1][9];
    ele[0][9] != ele[10][9];
    ele[0][9] != ele[11][9];
    ele[0][9] != ele[12][9];
    ele[0][9] != ele[13][9];
    ele[0][9] != ele[14][9];
    ele[0][9] != ele[15][9];
    ele[0][9] != ele[16][9];
    ele[0][9] != ele[17][9];
    ele[0][9] != ele[18][9];
    ele[0][9] != ele[19][9];
    ele[0][9] != ele[2][10];
    ele[0][9] != ele[2][11];
    ele[0][9] != ele[2][6];
    ele[0][9] != ele[2][7];
    ele[0][9] != ele[2][8];
    ele[0][9] != ele[2][9];
    ele[0][9] != ele[20][9];
    ele[0][9] != ele[21][9];
    ele[0][9] != ele[22][9];
    ele[0][9] != ele[23][9];
    ele[0][9] != ele[24][9];
    ele[0][9] != ele[25][9];
    ele[0][9] != ele[26][9];
    ele[0][9] != ele[27][9];
    ele[0][9] != ele[28][9];
    ele[0][9] != ele[29][9];
    ele[0][9] != ele[3][10];
    ele[0][9] != ele[3][11];
    ele[0][9] != ele[3][6];
    ele[0][9] != ele[3][7];
    ele[0][9] != ele[3][8];
    ele[0][9] != ele[3][9];
    ele[0][9] != ele[30][9];
    ele[0][9] != ele[31][9];
    ele[0][9] != ele[32][9];
    ele[0][9] != ele[33][9];
    ele[0][9] != ele[34][9];
    ele[0][9] != ele[35][9];
    ele[0][9] != ele[4][10];
    ele[0][9] != ele[4][11];
    ele[0][9] != ele[4][6];
    ele[0][9] != ele[4][7];
    ele[0][9] != ele[4][8];
    ele[0][9] != ele[4][9];
    ele[0][9] != ele[5][10];
    ele[0][9] != ele[5][11];
    ele[0][9] != ele[5][6];
    ele[0][9] != ele[5][7];
    ele[0][9] != ele[5][8];
    ele[0][9] != ele[5][9];
    ele[0][9] != ele[6][9];
    ele[0][9] != ele[7][9];
    ele[0][9] != ele[8][9];
    ele[0][9] != ele[9][9];
    ele[1][0] != ele[1][1];
    ele[1][0] != ele[1][10];
    ele[1][0] != ele[1][11];
    ele[1][0] != ele[1][12];
    ele[1][0] != ele[1][13];
    ele[1][0] != ele[1][14];
    ele[1][0] != ele[1][15];
    ele[1][0] != ele[1][16];
    ele[1][0] != ele[1][17];
    ele[1][0] != ele[1][18];
    ele[1][0] != ele[1][19];
    ele[1][0] != ele[1][2];
    ele[1][0] != ele[1][20];
    ele[1][0] != ele[1][21];
    ele[1][0] != ele[1][22];
    ele[1][0] != ele[1][23];
    ele[1][0] != ele[1][24];
    ele[1][0] != ele[1][25];
    ele[1][0] != ele[1][26];
    ele[1][0] != ele[1][27];
    ele[1][0] != ele[1][28];
    ele[1][0] != ele[1][29];
    ele[1][0] != ele[1][3];
    ele[1][0] != ele[1][30];
    ele[1][0] != ele[1][31];
    ele[1][0] != ele[1][32];
    ele[1][0] != ele[1][33];
    ele[1][0] != ele[1][34];
    ele[1][0] != ele[1][35];
    ele[1][0] != ele[1][4];
    ele[1][0] != ele[1][5];
    ele[1][0] != ele[1][6];
    ele[1][0] != ele[1][7];
    ele[1][0] != ele[1][8];
    ele[1][0] != ele[1][9];
    ele[1][0] != ele[10][0];
    ele[1][0] != ele[11][0];
    ele[1][0] != ele[12][0];
    ele[1][0] != ele[13][0];
    ele[1][0] != ele[14][0];
    ele[1][0] != ele[15][0];
    ele[1][0] != ele[16][0];
    ele[1][0] != ele[17][0];
    ele[1][0] != ele[18][0];
    ele[1][0] != ele[19][0];
    ele[1][0] != ele[2][0];
    ele[1][0] != ele[2][1];
    ele[1][0] != ele[2][2];
    ele[1][0] != ele[2][3];
    ele[1][0] != ele[2][4];
    ele[1][0] != ele[2][5];
    ele[1][0] != ele[20][0];
    ele[1][0] != ele[21][0];
    ele[1][0] != ele[22][0];
    ele[1][0] != ele[23][0];
    ele[1][0] != ele[24][0];
    ele[1][0] != ele[25][0];
    ele[1][0] != ele[26][0];
    ele[1][0] != ele[27][0];
    ele[1][0] != ele[28][0];
    ele[1][0] != ele[29][0];
    ele[1][0] != ele[3][0];
    ele[1][0] != ele[3][1];
    ele[1][0] != ele[3][2];
    ele[1][0] != ele[3][3];
    ele[1][0] != ele[3][4];
    ele[1][0] != ele[3][5];
    ele[1][0] != ele[30][0];
    ele[1][0] != ele[31][0];
    ele[1][0] != ele[32][0];
    ele[1][0] != ele[33][0];
    ele[1][0] != ele[34][0];
    ele[1][0] != ele[35][0];
    ele[1][0] != ele[4][0];
    ele[1][0] != ele[4][1];
    ele[1][0] != ele[4][2];
    ele[1][0] != ele[4][3];
    ele[1][0] != ele[4][4];
    ele[1][0] != ele[4][5];
    ele[1][0] != ele[5][0];
    ele[1][0] != ele[5][1];
    ele[1][0] != ele[5][2];
    ele[1][0] != ele[5][3];
    ele[1][0] != ele[5][4];
    ele[1][0] != ele[5][5];
    ele[1][0] != ele[6][0];
    ele[1][0] != ele[7][0];
    ele[1][0] != ele[8][0];
    ele[1][0] != ele[9][0];
    ele[1][1] != ele[1][10];
    ele[1][1] != ele[1][11];
    ele[1][1] != ele[1][12];
    ele[1][1] != ele[1][13];
    ele[1][1] != ele[1][14];
    ele[1][1] != ele[1][15];
    ele[1][1] != ele[1][16];
    ele[1][1] != ele[1][17];
    ele[1][1] != ele[1][18];
    ele[1][1] != ele[1][19];
    ele[1][1] != ele[1][2];
    ele[1][1] != ele[1][20];
    ele[1][1] != ele[1][21];
    ele[1][1] != ele[1][22];
    ele[1][1] != ele[1][23];
    ele[1][1] != ele[1][24];
    ele[1][1] != ele[1][25];
    ele[1][1] != ele[1][26];
    ele[1][1] != ele[1][27];
    ele[1][1] != ele[1][28];
    ele[1][1] != ele[1][29];
    ele[1][1] != ele[1][3];
    ele[1][1] != ele[1][30];
    ele[1][1] != ele[1][31];
    ele[1][1] != ele[1][32];
    ele[1][1] != ele[1][33];
    ele[1][1] != ele[1][34];
    ele[1][1] != ele[1][35];
    ele[1][1] != ele[1][4];
    ele[1][1] != ele[1][5];
    ele[1][1] != ele[1][6];
    ele[1][1] != ele[1][7];
    ele[1][1] != ele[1][8];
    ele[1][1] != ele[1][9];
    ele[1][1] != ele[10][1];
    ele[1][1] != ele[11][1];
    ele[1][1] != ele[12][1];
    ele[1][1] != ele[13][1];
    ele[1][1] != ele[14][1];
    ele[1][1] != ele[15][1];
    ele[1][1] != ele[16][1];
    ele[1][1] != ele[17][1];
    ele[1][1] != ele[18][1];
    ele[1][1] != ele[19][1];
    ele[1][1] != ele[2][0];
    ele[1][1] != ele[2][1];
    ele[1][1] != ele[2][2];
    ele[1][1] != ele[2][3];
    ele[1][1] != ele[2][4];
    ele[1][1] != ele[2][5];
    ele[1][1] != ele[20][1];
    ele[1][1] != ele[21][1];
    ele[1][1] != ele[22][1];
    ele[1][1] != ele[23][1];
    ele[1][1] != ele[24][1];
    ele[1][1] != ele[25][1];
    ele[1][1] != ele[26][1];
    ele[1][1] != ele[27][1];
    ele[1][1] != ele[28][1];
    ele[1][1] != ele[29][1];
    ele[1][1] != ele[3][0];
    ele[1][1] != ele[3][1];
    ele[1][1] != ele[3][2];
    ele[1][1] != ele[3][3];
    ele[1][1] != ele[3][4];
    ele[1][1] != ele[3][5];
    ele[1][1] != ele[30][1];
    ele[1][1] != ele[31][1];
    ele[1][1] != ele[32][1];
    ele[1][1] != ele[33][1];
    ele[1][1] != ele[34][1];
    ele[1][1] != ele[35][1];
    ele[1][1] != ele[4][0];
    ele[1][1] != ele[4][1];
    ele[1][1] != ele[4][2];
    ele[1][1] != ele[4][3];
    ele[1][1] != ele[4][4];
    ele[1][1] != ele[4][5];
    ele[1][1] != ele[5][0];
    ele[1][1] != ele[5][1];
    ele[1][1] != ele[5][2];
    ele[1][1] != ele[5][3];
    ele[1][1] != ele[5][4];
    ele[1][1] != ele[5][5];
    ele[1][1] != ele[6][1];
    ele[1][1] != ele[7][1];
    ele[1][1] != ele[8][1];
    ele[1][1] != ele[9][1];
    ele[1][10] != ele[1][11];
    ele[1][10] != ele[1][12];
    ele[1][10] != ele[1][13];
    ele[1][10] != ele[1][14];
    ele[1][10] != ele[1][15];
    ele[1][10] != ele[1][16];
    ele[1][10] != ele[1][17];
    ele[1][10] != ele[1][18];
    ele[1][10] != ele[1][19];
    ele[1][10] != ele[1][20];
    ele[1][10] != ele[1][21];
    ele[1][10] != ele[1][22];
    ele[1][10] != ele[1][23];
    ele[1][10] != ele[1][24];
    ele[1][10] != ele[1][25];
    ele[1][10] != ele[1][26];
    ele[1][10] != ele[1][27];
    ele[1][10] != ele[1][28];
    ele[1][10] != ele[1][29];
    ele[1][10] != ele[1][30];
    ele[1][10] != ele[1][31];
    ele[1][10] != ele[1][32];
    ele[1][10] != ele[1][33];
    ele[1][10] != ele[1][34];
    ele[1][10] != ele[1][35];
    ele[1][10] != ele[10][10];
    ele[1][10] != ele[11][10];
    ele[1][10] != ele[12][10];
    ele[1][10] != ele[13][10];
    ele[1][10] != ele[14][10];
    ele[1][10] != ele[15][10];
    ele[1][10] != ele[16][10];
    ele[1][10] != ele[17][10];
    ele[1][10] != ele[18][10];
    ele[1][10] != ele[19][10];
    ele[1][10] != ele[2][10];
    ele[1][10] != ele[2][11];
    ele[1][10] != ele[2][6];
    ele[1][10] != ele[2][7];
    ele[1][10] != ele[2][8];
    ele[1][10] != ele[2][9];
    ele[1][10] != ele[20][10];
    ele[1][10] != ele[21][10];
    ele[1][10] != ele[22][10];
    ele[1][10] != ele[23][10];
    ele[1][10] != ele[24][10];
    ele[1][10] != ele[25][10];
    ele[1][10] != ele[26][10];
    ele[1][10] != ele[27][10];
    ele[1][10] != ele[28][10];
    ele[1][10] != ele[29][10];
    ele[1][10] != ele[3][10];
    ele[1][10] != ele[3][11];
    ele[1][10] != ele[3][6];
    ele[1][10] != ele[3][7];
    ele[1][10] != ele[3][8];
    ele[1][10] != ele[3][9];
    ele[1][10] != ele[30][10];
    ele[1][10] != ele[31][10];
    ele[1][10] != ele[32][10];
    ele[1][10] != ele[33][10];
    ele[1][10] != ele[34][10];
    ele[1][10] != ele[35][10];
    ele[1][10] != ele[4][10];
    ele[1][10] != ele[4][11];
    ele[1][10] != ele[4][6];
    ele[1][10] != ele[4][7];
    ele[1][10] != ele[4][8];
    ele[1][10] != ele[4][9];
    ele[1][10] != ele[5][10];
    ele[1][10] != ele[5][11];
    ele[1][10] != ele[5][6];
    ele[1][10] != ele[5][7];
    ele[1][10] != ele[5][8];
    ele[1][10] != ele[5][9];
    ele[1][10] != ele[6][10];
    ele[1][10] != ele[7][10];
    ele[1][10] != ele[8][10];
    ele[1][10] != ele[9][10];
    ele[1][11] != ele[1][12];
    ele[1][11] != ele[1][13];
    ele[1][11] != ele[1][14];
    ele[1][11] != ele[1][15];
    ele[1][11] != ele[1][16];
    ele[1][11] != ele[1][17];
    ele[1][11] != ele[1][18];
    ele[1][11] != ele[1][19];
    ele[1][11] != ele[1][20];
    ele[1][11] != ele[1][21];
    ele[1][11] != ele[1][22];
    ele[1][11] != ele[1][23];
    ele[1][11] != ele[1][24];
    ele[1][11] != ele[1][25];
    ele[1][11] != ele[1][26];
    ele[1][11] != ele[1][27];
    ele[1][11] != ele[1][28];
    ele[1][11] != ele[1][29];
    ele[1][11] != ele[1][30];
    ele[1][11] != ele[1][31];
    ele[1][11] != ele[1][32];
    ele[1][11] != ele[1][33];
    ele[1][11] != ele[1][34];
    ele[1][11] != ele[1][35];
    ele[1][11] != ele[10][11];
    ele[1][11] != ele[11][11];
    ele[1][11] != ele[12][11];
    ele[1][11] != ele[13][11];
    ele[1][11] != ele[14][11];
    ele[1][11] != ele[15][11];
    ele[1][11] != ele[16][11];
    ele[1][11] != ele[17][11];
    ele[1][11] != ele[18][11];
    ele[1][11] != ele[19][11];
    ele[1][11] != ele[2][10];
    ele[1][11] != ele[2][11];
    ele[1][11] != ele[2][6];
    ele[1][11] != ele[2][7];
    ele[1][11] != ele[2][8];
    ele[1][11] != ele[2][9];
    ele[1][11] != ele[20][11];
    ele[1][11] != ele[21][11];
    ele[1][11] != ele[22][11];
    ele[1][11] != ele[23][11];
    ele[1][11] != ele[24][11];
    ele[1][11] != ele[25][11];
    ele[1][11] != ele[26][11];
    ele[1][11] != ele[27][11];
    ele[1][11] != ele[28][11];
    ele[1][11] != ele[29][11];
    ele[1][11] != ele[3][10];
    ele[1][11] != ele[3][11];
    ele[1][11] != ele[3][6];
    ele[1][11] != ele[3][7];
    ele[1][11] != ele[3][8];
    ele[1][11] != ele[3][9];
    ele[1][11] != ele[30][11];
    ele[1][11] != ele[31][11];
    ele[1][11] != ele[32][11];
    ele[1][11] != ele[33][11];
    ele[1][11] != ele[34][11];
    ele[1][11] != ele[35][11];
    ele[1][11] != ele[4][10];
    ele[1][11] != ele[4][11];
    ele[1][11] != ele[4][6];
    ele[1][11] != ele[4][7];
    ele[1][11] != ele[4][8];
    ele[1][11] != ele[4][9];
    ele[1][11] != ele[5][10];
    ele[1][11] != ele[5][11];
    ele[1][11] != ele[5][6];
    ele[1][11] != ele[5][7];
    ele[1][11] != ele[5][8];
    ele[1][11] != ele[5][9];
    ele[1][11] != ele[6][11];
    ele[1][11] != ele[7][11];
    ele[1][11] != ele[8][11];
    ele[1][11] != ele[9][11];
    ele[1][12] != ele[1][13];
    ele[1][12] != ele[1][14];
    ele[1][12] != ele[1][15];
    ele[1][12] != ele[1][16];
    ele[1][12] != ele[1][17];
    ele[1][12] != ele[1][18];
    ele[1][12] != ele[1][19];
    ele[1][12] != ele[1][20];
    ele[1][12] != ele[1][21];
    ele[1][12] != ele[1][22];
    ele[1][12] != ele[1][23];
    ele[1][12] != ele[1][24];
    ele[1][12] != ele[1][25];
    ele[1][12] != ele[1][26];
    ele[1][12] != ele[1][27];
    ele[1][12] != ele[1][28];
    ele[1][12] != ele[1][29];
    ele[1][12] != ele[1][30];
    ele[1][12] != ele[1][31];
    ele[1][12] != ele[1][32];
    ele[1][12] != ele[1][33];
    ele[1][12] != ele[1][34];
    ele[1][12] != ele[1][35];
    ele[1][12] != ele[10][12];
    ele[1][12] != ele[11][12];
    ele[1][12] != ele[12][12];
    ele[1][12] != ele[13][12];
    ele[1][12] != ele[14][12];
    ele[1][12] != ele[15][12];
    ele[1][12] != ele[16][12];
    ele[1][12] != ele[17][12];
    ele[1][12] != ele[18][12];
    ele[1][12] != ele[19][12];
    ele[1][12] != ele[2][12];
    ele[1][12] != ele[2][13];
    ele[1][12] != ele[2][14];
    ele[1][12] != ele[2][15];
    ele[1][12] != ele[2][16];
    ele[1][12] != ele[2][17];
    ele[1][12] != ele[20][12];
    ele[1][12] != ele[21][12];
    ele[1][12] != ele[22][12];
    ele[1][12] != ele[23][12];
    ele[1][12] != ele[24][12];
    ele[1][12] != ele[25][12];
    ele[1][12] != ele[26][12];
    ele[1][12] != ele[27][12];
    ele[1][12] != ele[28][12];
    ele[1][12] != ele[29][12];
    ele[1][12] != ele[3][12];
    ele[1][12] != ele[3][13];
    ele[1][12] != ele[3][14];
    ele[1][12] != ele[3][15];
    ele[1][12] != ele[3][16];
    ele[1][12] != ele[3][17];
    ele[1][12] != ele[30][12];
    ele[1][12] != ele[31][12];
    ele[1][12] != ele[32][12];
    ele[1][12] != ele[33][12];
    ele[1][12] != ele[34][12];
    ele[1][12] != ele[35][12];
    ele[1][12] != ele[4][12];
    ele[1][12] != ele[4][13];
    ele[1][12] != ele[4][14];
    ele[1][12] != ele[4][15];
    ele[1][12] != ele[4][16];
    ele[1][12] != ele[4][17];
    ele[1][12] != ele[5][12];
    ele[1][12] != ele[5][13];
    ele[1][12] != ele[5][14];
    ele[1][12] != ele[5][15];
    ele[1][12] != ele[5][16];
    ele[1][12] != ele[5][17];
    ele[1][12] != ele[6][12];
    ele[1][12] != ele[7][12];
    ele[1][12] != ele[8][12];
    ele[1][12] != ele[9][12];
    ele[1][13] != ele[1][14];
    ele[1][13] != ele[1][15];
    ele[1][13] != ele[1][16];
    ele[1][13] != ele[1][17];
    ele[1][13] != ele[1][18];
    ele[1][13] != ele[1][19];
    ele[1][13] != ele[1][20];
    ele[1][13] != ele[1][21];
    ele[1][13] != ele[1][22];
    ele[1][13] != ele[1][23];
    ele[1][13] != ele[1][24];
    ele[1][13] != ele[1][25];
    ele[1][13] != ele[1][26];
    ele[1][13] != ele[1][27];
    ele[1][13] != ele[1][28];
    ele[1][13] != ele[1][29];
    ele[1][13] != ele[1][30];
    ele[1][13] != ele[1][31];
    ele[1][13] != ele[1][32];
    ele[1][13] != ele[1][33];
    ele[1][13] != ele[1][34];
    ele[1][13] != ele[1][35];
    ele[1][13] != ele[10][13];
    ele[1][13] != ele[11][13];
    ele[1][13] != ele[12][13];
    ele[1][13] != ele[13][13];
    ele[1][13] != ele[14][13];
    ele[1][13] != ele[15][13];
    ele[1][13] != ele[16][13];
    ele[1][13] != ele[17][13];
    ele[1][13] != ele[18][13];
    ele[1][13] != ele[19][13];
    ele[1][13] != ele[2][12];
    ele[1][13] != ele[2][13];
    ele[1][13] != ele[2][14];
    ele[1][13] != ele[2][15];
    ele[1][13] != ele[2][16];
    ele[1][13] != ele[2][17];
    ele[1][13] != ele[20][13];
    ele[1][13] != ele[21][13];
    ele[1][13] != ele[22][13];
    ele[1][13] != ele[23][13];
    ele[1][13] != ele[24][13];
    ele[1][13] != ele[25][13];
    ele[1][13] != ele[26][13];
    ele[1][13] != ele[27][13];
    ele[1][13] != ele[28][13];
    ele[1][13] != ele[29][13];
    ele[1][13] != ele[3][12];
    ele[1][13] != ele[3][13];
    ele[1][13] != ele[3][14];
    ele[1][13] != ele[3][15];
    ele[1][13] != ele[3][16];
    ele[1][13] != ele[3][17];
    ele[1][13] != ele[30][13];
    ele[1][13] != ele[31][13];
    ele[1][13] != ele[32][13];
    ele[1][13] != ele[33][13];
    ele[1][13] != ele[34][13];
    ele[1][13] != ele[35][13];
    ele[1][13] != ele[4][12];
    ele[1][13] != ele[4][13];
    ele[1][13] != ele[4][14];
    ele[1][13] != ele[4][15];
    ele[1][13] != ele[4][16];
    ele[1][13] != ele[4][17];
    ele[1][13] != ele[5][12];
    ele[1][13] != ele[5][13];
    ele[1][13] != ele[5][14];
    ele[1][13] != ele[5][15];
    ele[1][13] != ele[5][16];
    ele[1][13] != ele[5][17];
    ele[1][13] != ele[6][13];
    ele[1][13] != ele[7][13];
    ele[1][13] != ele[8][13];
    ele[1][13] != ele[9][13];
    ele[1][14] != ele[1][15];
    ele[1][14] != ele[1][16];
    ele[1][14] != ele[1][17];
    ele[1][14] != ele[1][18];
    ele[1][14] != ele[1][19];
    ele[1][14] != ele[1][20];
    ele[1][14] != ele[1][21];
    ele[1][14] != ele[1][22];
    ele[1][14] != ele[1][23];
    ele[1][14] != ele[1][24];
    ele[1][14] != ele[1][25];
    ele[1][14] != ele[1][26];
    ele[1][14] != ele[1][27];
    ele[1][14] != ele[1][28];
    ele[1][14] != ele[1][29];
    ele[1][14] != ele[1][30];
    ele[1][14] != ele[1][31];
    ele[1][14] != ele[1][32];
    ele[1][14] != ele[1][33];
    ele[1][14] != ele[1][34];
    ele[1][14] != ele[1][35];
    ele[1][14] != ele[10][14];
    ele[1][14] != ele[11][14];
    ele[1][14] != ele[12][14];
    ele[1][14] != ele[13][14];
    ele[1][14] != ele[14][14];
    ele[1][14] != ele[15][14];
    ele[1][14] != ele[16][14];
    ele[1][14] != ele[17][14];
    ele[1][14] != ele[18][14];
    ele[1][14] != ele[19][14];
    ele[1][14] != ele[2][12];
    ele[1][14] != ele[2][13];
    ele[1][14] != ele[2][14];
    ele[1][14] != ele[2][15];
    ele[1][14] != ele[2][16];
    ele[1][14] != ele[2][17];
    ele[1][14] != ele[20][14];
    ele[1][14] != ele[21][14];
    ele[1][14] != ele[22][14];
    ele[1][14] != ele[23][14];
    ele[1][14] != ele[24][14];
    ele[1][14] != ele[25][14];
    ele[1][14] != ele[26][14];
    ele[1][14] != ele[27][14];
    ele[1][14] != ele[28][14];
    ele[1][14] != ele[29][14];
    ele[1][14] != ele[3][12];
    ele[1][14] != ele[3][13];
    ele[1][14] != ele[3][14];
    ele[1][14] != ele[3][15];
    ele[1][14] != ele[3][16];
    ele[1][14] != ele[3][17];
    ele[1][14] != ele[30][14];
    ele[1][14] != ele[31][14];
    ele[1][14] != ele[32][14];
    ele[1][14] != ele[33][14];
    ele[1][14] != ele[34][14];
    ele[1][14] != ele[35][14];
    ele[1][14] != ele[4][12];
    ele[1][14] != ele[4][13];
    ele[1][14] != ele[4][14];
    ele[1][14] != ele[4][15];
    ele[1][14] != ele[4][16];
    ele[1][14] != ele[4][17];
    ele[1][14] != ele[5][12];
    ele[1][14] != ele[5][13];
    ele[1][14] != ele[5][14];
    ele[1][14] != ele[5][15];
    ele[1][14] != ele[5][16];
    ele[1][14] != ele[5][17];
    ele[1][14] != ele[6][14];
    ele[1][14] != ele[7][14];
    ele[1][14] != ele[8][14];
    ele[1][14] != ele[9][14];
    ele[1][15] != ele[1][16];
    ele[1][15] != ele[1][17];
    ele[1][15] != ele[1][18];
    ele[1][15] != ele[1][19];
    ele[1][15] != ele[1][20];
    ele[1][15] != ele[1][21];
    ele[1][15] != ele[1][22];
    ele[1][15] != ele[1][23];
    ele[1][15] != ele[1][24];
    ele[1][15] != ele[1][25];
    ele[1][15] != ele[1][26];
    ele[1][15] != ele[1][27];
    ele[1][15] != ele[1][28];
    ele[1][15] != ele[1][29];
    ele[1][15] != ele[1][30];
    ele[1][15] != ele[1][31];
    ele[1][15] != ele[1][32];
    ele[1][15] != ele[1][33];
    ele[1][15] != ele[1][34];
    ele[1][15] != ele[1][35];
    ele[1][15] != ele[10][15];
    ele[1][15] != ele[11][15];
    ele[1][15] != ele[12][15];
    ele[1][15] != ele[13][15];
    ele[1][15] != ele[14][15];
    ele[1][15] != ele[15][15];
    ele[1][15] != ele[16][15];
    ele[1][15] != ele[17][15];
    ele[1][15] != ele[18][15];
    ele[1][15] != ele[19][15];
    ele[1][15] != ele[2][12];
    ele[1][15] != ele[2][13];
    ele[1][15] != ele[2][14];
    ele[1][15] != ele[2][15];
    ele[1][15] != ele[2][16];
    ele[1][15] != ele[2][17];
    ele[1][15] != ele[20][15];
    ele[1][15] != ele[21][15];
    ele[1][15] != ele[22][15];
    ele[1][15] != ele[23][15];
    ele[1][15] != ele[24][15];
    ele[1][15] != ele[25][15];
    ele[1][15] != ele[26][15];
    ele[1][15] != ele[27][15];
    ele[1][15] != ele[28][15];
    ele[1][15] != ele[29][15];
    ele[1][15] != ele[3][12];
    ele[1][15] != ele[3][13];
    ele[1][15] != ele[3][14];
    ele[1][15] != ele[3][15];
    ele[1][15] != ele[3][16];
    ele[1][15] != ele[3][17];
    ele[1][15] != ele[30][15];
    ele[1][15] != ele[31][15];
    ele[1][15] != ele[32][15];
    ele[1][15] != ele[33][15];
    ele[1][15] != ele[34][15];
    ele[1][15] != ele[35][15];
    ele[1][15] != ele[4][12];
    ele[1][15] != ele[4][13];
    ele[1][15] != ele[4][14];
    ele[1][15] != ele[4][15];
    ele[1][15] != ele[4][16];
    ele[1][15] != ele[4][17];
    ele[1][15] != ele[5][12];
    ele[1][15] != ele[5][13];
    ele[1][15] != ele[5][14];
    ele[1][15] != ele[5][15];
    ele[1][15] != ele[5][16];
    ele[1][15] != ele[5][17];
    ele[1][15] != ele[6][15];
    ele[1][15] != ele[7][15];
    ele[1][15] != ele[8][15];
    ele[1][15] != ele[9][15];
    ele[1][16] != ele[1][17];
    ele[1][16] != ele[1][18];
    ele[1][16] != ele[1][19];
    ele[1][16] != ele[1][20];
    ele[1][16] != ele[1][21];
    ele[1][16] != ele[1][22];
    ele[1][16] != ele[1][23];
    ele[1][16] != ele[1][24];
    ele[1][16] != ele[1][25];
    ele[1][16] != ele[1][26];
    ele[1][16] != ele[1][27];
    ele[1][16] != ele[1][28];
    ele[1][16] != ele[1][29];
    ele[1][16] != ele[1][30];
    ele[1][16] != ele[1][31];
    ele[1][16] != ele[1][32];
    ele[1][16] != ele[1][33];
    ele[1][16] != ele[1][34];
    ele[1][16] != ele[1][35];
    ele[1][16] != ele[10][16];
    ele[1][16] != ele[11][16];
    ele[1][16] != ele[12][16];
    ele[1][16] != ele[13][16];
    ele[1][16] != ele[14][16];
    ele[1][16] != ele[15][16];
    ele[1][16] != ele[16][16];
    ele[1][16] != ele[17][16];
    ele[1][16] != ele[18][16];
    ele[1][16] != ele[19][16];
    ele[1][16] != ele[2][12];
    ele[1][16] != ele[2][13];
    ele[1][16] != ele[2][14];
    ele[1][16] != ele[2][15];
    ele[1][16] != ele[2][16];
    ele[1][16] != ele[2][17];
    ele[1][16] != ele[20][16];
    ele[1][16] != ele[21][16];
    ele[1][16] != ele[22][16];
    ele[1][16] != ele[23][16];
    ele[1][16] != ele[24][16];
    ele[1][16] != ele[25][16];
    ele[1][16] != ele[26][16];
    ele[1][16] != ele[27][16];
    ele[1][16] != ele[28][16];
    ele[1][16] != ele[29][16];
    ele[1][16] != ele[3][12];
    ele[1][16] != ele[3][13];
    ele[1][16] != ele[3][14];
    ele[1][16] != ele[3][15];
    ele[1][16] != ele[3][16];
    ele[1][16] != ele[3][17];
    ele[1][16] != ele[30][16];
    ele[1][16] != ele[31][16];
    ele[1][16] != ele[32][16];
    ele[1][16] != ele[33][16];
    ele[1][16] != ele[34][16];
    ele[1][16] != ele[35][16];
    ele[1][16] != ele[4][12];
    ele[1][16] != ele[4][13];
    ele[1][16] != ele[4][14];
    ele[1][16] != ele[4][15];
    ele[1][16] != ele[4][16];
    ele[1][16] != ele[4][17];
    ele[1][16] != ele[5][12];
    ele[1][16] != ele[5][13];
    ele[1][16] != ele[5][14];
    ele[1][16] != ele[5][15];
    ele[1][16] != ele[5][16];
    ele[1][16] != ele[5][17];
    ele[1][16] != ele[6][16];
    ele[1][16] != ele[7][16];
    ele[1][16] != ele[8][16];
    ele[1][16] != ele[9][16];
    ele[1][17] != ele[1][18];
    ele[1][17] != ele[1][19];
    ele[1][17] != ele[1][20];
    ele[1][17] != ele[1][21];
    ele[1][17] != ele[1][22];
    ele[1][17] != ele[1][23];
    ele[1][17] != ele[1][24];
    ele[1][17] != ele[1][25];
    ele[1][17] != ele[1][26];
    ele[1][17] != ele[1][27];
    ele[1][17] != ele[1][28];
    ele[1][17] != ele[1][29];
    ele[1][17] != ele[1][30];
    ele[1][17] != ele[1][31];
    ele[1][17] != ele[1][32];
    ele[1][17] != ele[1][33];
    ele[1][17] != ele[1][34];
    ele[1][17] != ele[1][35];
    ele[1][17] != ele[10][17];
    ele[1][17] != ele[11][17];
    ele[1][17] != ele[12][17];
    ele[1][17] != ele[13][17];
    ele[1][17] != ele[14][17];
    ele[1][17] != ele[15][17];
    ele[1][17] != ele[16][17];
    ele[1][17] != ele[17][17];
    ele[1][17] != ele[18][17];
    ele[1][17] != ele[19][17];
    ele[1][17] != ele[2][12];
    ele[1][17] != ele[2][13];
    ele[1][17] != ele[2][14];
    ele[1][17] != ele[2][15];
    ele[1][17] != ele[2][16];
    ele[1][17] != ele[2][17];
    ele[1][17] != ele[20][17];
    ele[1][17] != ele[21][17];
    ele[1][17] != ele[22][17];
    ele[1][17] != ele[23][17];
    ele[1][17] != ele[24][17];
    ele[1][17] != ele[25][17];
    ele[1][17] != ele[26][17];
    ele[1][17] != ele[27][17];
    ele[1][17] != ele[28][17];
    ele[1][17] != ele[29][17];
    ele[1][17] != ele[3][12];
    ele[1][17] != ele[3][13];
    ele[1][17] != ele[3][14];
    ele[1][17] != ele[3][15];
    ele[1][17] != ele[3][16];
    ele[1][17] != ele[3][17];
    ele[1][17] != ele[30][17];
    ele[1][17] != ele[31][17];
    ele[1][17] != ele[32][17];
    ele[1][17] != ele[33][17];
    ele[1][17] != ele[34][17];
    ele[1][17] != ele[35][17];
    ele[1][17] != ele[4][12];
    ele[1][17] != ele[4][13];
    ele[1][17] != ele[4][14];
    ele[1][17] != ele[4][15];
    ele[1][17] != ele[4][16];
    ele[1][17] != ele[4][17];
    ele[1][17] != ele[5][12];
    ele[1][17] != ele[5][13];
    ele[1][17] != ele[5][14];
    ele[1][17] != ele[5][15];
    ele[1][17] != ele[5][16];
    ele[1][17] != ele[5][17];
    ele[1][17] != ele[6][17];
    ele[1][17] != ele[7][17];
    ele[1][17] != ele[8][17];
    ele[1][17] != ele[9][17];
    ele[1][18] != ele[1][19];
    ele[1][18] != ele[1][20];
    ele[1][18] != ele[1][21];
    ele[1][18] != ele[1][22];
    ele[1][18] != ele[1][23];
    ele[1][18] != ele[1][24];
    ele[1][18] != ele[1][25];
    ele[1][18] != ele[1][26];
    ele[1][18] != ele[1][27];
    ele[1][18] != ele[1][28];
    ele[1][18] != ele[1][29];
    ele[1][18] != ele[1][30];
    ele[1][18] != ele[1][31];
    ele[1][18] != ele[1][32];
    ele[1][18] != ele[1][33];
    ele[1][18] != ele[1][34];
    ele[1][18] != ele[1][35];
    ele[1][18] != ele[10][18];
    ele[1][18] != ele[11][18];
    ele[1][18] != ele[12][18];
    ele[1][18] != ele[13][18];
    ele[1][18] != ele[14][18];
    ele[1][18] != ele[15][18];
    ele[1][18] != ele[16][18];
    ele[1][18] != ele[17][18];
    ele[1][18] != ele[18][18];
    ele[1][18] != ele[19][18];
    ele[1][18] != ele[2][18];
    ele[1][18] != ele[2][19];
    ele[1][18] != ele[2][20];
    ele[1][18] != ele[2][21];
    ele[1][18] != ele[2][22];
    ele[1][18] != ele[2][23];
    ele[1][18] != ele[20][18];
    ele[1][18] != ele[21][18];
    ele[1][18] != ele[22][18];
    ele[1][18] != ele[23][18];
    ele[1][18] != ele[24][18];
    ele[1][18] != ele[25][18];
    ele[1][18] != ele[26][18];
    ele[1][18] != ele[27][18];
    ele[1][18] != ele[28][18];
    ele[1][18] != ele[29][18];
    ele[1][18] != ele[3][18];
    ele[1][18] != ele[3][19];
    ele[1][18] != ele[3][20];
    ele[1][18] != ele[3][21];
    ele[1][18] != ele[3][22];
    ele[1][18] != ele[3][23];
    ele[1][18] != ele[30][18];
    ele[1][18] != ele[31][18];
    ele[1][18] != ele[32][18];
    ele[1][18] != ele[33][18];
    ele[1][18] != ele[34][18];
    ele[1][18] != ele[35][18];
    ele[1][18] != ele[4][18];
    ele[1][18] != ele[4][19];
    ele[1][18] != ele[4][20];
    ele[1][18] != ele[4][21];
    ele[1][18] != ele[4][22];
    ele[1][18] != ele[4][23];
    ele[1][18] != ele[5][18];
    ele[1][18] != ele[5][19];
    ele[1][18] != ele[5][20];
    ele[1][18] != ele[5][21];
    ele[1][18] != ele[5][22];
    ele[1][18] != ele[5][23];
    ele[1][18] != ele[6][18];
    ele[1][18] != ele[7][18];
    ele[1][18] != ele[8][18];
    ele[1][18] != ele[9][18];
    ele[1][19] != ele[1][20];
    ele[1][19] != ele[1][21];
    ele[1][19] != ele[1][22];
    ele[1][19] != ele[1][23];
    ele[1][19] != ele[1][24];
    ele[1][19] != ele[1][25];
    ele[1][19] != ele[1][26];
    ele[1][19] != ele[1][27];
    ele[1][19] != ele[1][28];
    ele[1][19] != ele[1][29];
    ele[1][19] != ele[1][30];
    ele[1][19] != ele[1][31];
    ele[1][19] != ele[1][32];
    ele[1][19] != ele[1][33];
    ele[1][19] != ele[1][34];
    ele[1][19] != ele[1][35];
    ele[1][19] != ele[10][19];
    ele[1][19] != ele[11][19];
    ele[1][19] != ele[12][19];
    ele[1][19] != ele[13][19];
    ele[1][19] != ele[14][19];
    ele[1][19] != ele[15][19];
    ele[1][19] != ele[16][19];
    ele[1][19] != ele[17][19];
    ele[1][19] != ele[18][19];
    ele[1][19] != ele[19][19];
    ele[1][19] != ele[2][18];
    ele[1][19] != ele[2][19];
    ele[1][19] != ele[2][20];
    ele[1][19] != ele[2][21];
    ele[1][19] != ele[2][22];
    ele[1][19] != ele[2][23];
    ele[1][19] != ele[20][19];
    ele[1][19] != ele[21][19];
    ele[1][19] != ele[22][19];
    ele[1][19] != ele[23][19];
    ele[1][19] != ele[24][19];
    ele[1][19] != ele[25][19];
    ele[1][19] != ele[26][19];
    ele[1][19] != ele[27][19];
    ele[1][19] != ele[28][19];
    ele[1][19] != ele[29][19];
    ele[1][19] != ele[3][18];
    ele[1][19] != ele[3][19];
    ele[1][19] != ele[3][20];
    ele[1][19] != ele[3][21];
    ele[1][19] != ele[3][22];
    ele[1][19] != ele[3][23];
    ele[1][19] != ele[30][19];
    ele[1][19] != ele[31][19];
    ele[1][19] != ele[32][19];
    ele[1][19] != ele[33][19];
    ele[1][19] != ele[34][19];
    ele[1][19] != ele[35][19];
    ele[1][19] != ele[4][18];
    ele[1][19] != ele[4][19];
    ele[1][19] != ele[4][20];
    ele[1][19] != ele[4][21];
    ele[1][19] != ele[4][22];
    ele[1][19] != ele[4][23];
    ele[1][19] != ele[5][18];
    ele[1][19] != ele[5][19];
    ele[1][19] != ele[5][20];
    ele[1][19] != ele[5][21];
    ele[1][19] != ele[5][22];
    ele[1][19] != ele[5][23];
    ele[1][19] != ele[6][19];
    ele[1][19] != ele[7][19];
    ele[1][19] != ele[8][19];
    ele[1][19] != ele[9][19];
    ele[1][2] != ele[1][10];
    ele[1][2] != ele[1][11];
    ele[1][2] != ele[1][12];
    ele[1][2] != ele[1][13];
    ele[1][2] != ele[1][14];
    ele[1][2] != ele[1][15];
    ele[1][2] != ele[1][16];
    ele[1][2] != ele[1][17];
    ele[1][2] != ele[1][18];
    ele[1][2] != ele[1][19];
    ele[1][2] != ele[1][20];
    ele[1][2] != ele[1][21];
    ele[1][2] != ele[1][22];
    ele[1][2] != ele[1][23];
    ele[1][2] != ele[1][24];
    ele[1][2] != ele[1][25];
    ele[1][2] != ele[1][26];
    ele[1][2] != ele[1][27];
    ele[1][2] != ele[1][28];
    ele[1][2] != ele[1][29];
    ele[1][2] != ele[1][3];
    ele[1][2] != ele[1][30];
    ele[1][2] != ele[1][31];
    ele[1][2] != ele[1][32];
    ele[1][2] != ele[1][33];
    ele[1][2] != ele[1][34];
    ele[1][2] != ele[1][35];
    ele[1][2] != ele[1][4];
    ele[1][2] != ele[1][5];
    ele[1][2] != ele[1][6];
    ele[1][2] != ele[1][7];
    ele[1][2] != ele[1][8];
    ele[1][2] != ele[1][9];
    ele[1][2] != ele[10][2];
    ele[1][2] != ele[11][2];
    ele[1][2] != ele[12][2];
    ele[1][2] != ele[13][2];
    ele[1][2] != ele[14][2];
    ele[1][2] != ele[15][2];
    ele[1][2] != ele[16][2];
    ele[1][2] != ele[17][2];
    ele[1][2] != ele[18][2];
    ele[1][2] != ele[19][2];
    ele[1][2] != ele[2][0];
    ele[1][2] != ele[2][1];
    ele[1][2] != ele[2][2];
    ele[1][2] != ele[2][3];
    ele[1][2] != ele[2][4];
    ele[1][2] != ele[2][5];
    ele[1][2] != ele[20][2];
    ele[1][2] != ele[21][2];
    ele[1][2] != ele[22][2];
    ele[1][2] != ele[23][2];
    ele[1][2] != ele[24][2];
    ele[1][2] != ele[25][2];
    ele[1][2] != ele[26][2];
    ele[1][2] != ele[27][2];
    ele[1][2] != ele[28][2];
    ele[1][2] != ele[29][2];
    ele[1][2] != ele[3][0];
    ele[1][2] != ele[3][1];
    ele[1][2] != ele[3][2];
    ele[1][2] != ele[3][3];
    ele[1][2] != ele[3][4];
    ele[1][2] != ele[3][5];
    ele[1][2] != ele[30][2];
    ele[1][2] != ele[31][2];
    ele[1][2] != ele[32][2];
    ele[1][2] != ele[33][2];
    ele[1][2] != ele[34][2];
    ele[1][2] != ele[35][2];
    ele[1][2] != ele[4][0];
    ele[1][2] != ele[4][1];
    ele[1][2] != ele[4][2];
    ele[1][2] != ele[4][3];
    ele[1][2] != ele[4][4];
    ele[1][2] != ele[4][5];
    ele[1][2] != ele[5][0];
    ele[1][2] != ele[5][1];
    ele[1][2] != ele[5][2];
    ele[1][2] != ele[5][3];
    ele[1][2] != ele[5][4];
    ele[1][2] != ele[5][5];
    ele[1][2] != ele[6][2];
    ele[1][2] != ele[7][2];
    ele[1][2] != ele[8][2];
    ele[1][2] != ele[9][2];
    ele[1][20] != ele[1][21];
    ele[1][20] != ele[1][22];
    ele[1][20] != ele[1][23];
    ele[1][20] != ele[1][24];
    ele[1][20] != ele[1][25];
    ele[1][20] != ele[1][26];
    ele[1][20] != ele[1][27];
    ele[1][20] != ele[1][28];
    ele[1][20] != ele[1][29];
    ele[1][20] != ele[1][30];
    ele[1][20] != ele[1][31];
    ele[1][20] != ele[1][32];
    ele[1][20] != ele[1][33];
    ele[1][20] != ele[1][34];
    ele[1][20] != ele[1][35];
    ele[1][20] != ele[10][20];
    ele[1][20] != ele[11][20];
    ele[1][20] != ele[12][20];
    ele[1][20] != ele[13][20];
    ele[1][20] != ele[14][20];
    ele[1][20] != ele[15][20];
    ele[1][20] != ele[16][20];
    ele[1][20] != ele[17][20];
    ele[1][20] != ele[18][20];
    ele[1][20] != ele[19][20];
    ele[1][20] != ele[2][18];
    ele[1][20] != ele[2][19];
    ele[1][20] != ele[2][20];
    ele[1][20] != ele[2][21];
    ele[1][20] != ele[2][22];
    ele[1][20] != ele[2][23];
    ele[1][20] != ele[20][20];
    ele[1][20] != ele[21][20];
    ele[1][20] != ele[22][20];
    ele[1][20] != ele[23][20];
    ele[1][20] != ele[24][20];
    ele[1][20] != ele[25][20];
    ele[1][20] != ele[26][20];
    ele[1][20] != ele[27][20];
    ele[1][20] != ele[28][20];
    ele[1][20] != ele[29][20];
    ele[1][20] != ele[3][18];
    ele[1][20] != ele[3][19];
    ele[1][20] != ele[3][20];
    ele[1][20] != ele[3][21];
    ele[1][20] != ele[3][22];
    ele[1][20] != ele[3][23];
    ele[1][20] != ele[30][20];
    ele[1][20] != ele[31][20];
    ele[1][20] != ele[32][20];
    ele[1][20] != ele[33][20];
    ele[1][20] != ele[34][20];
    ele[1][20] != ele[35][20];
    ele[1][20] != ele[4][18];
    ele[1][20] != ele[4][19];
    ele[1][20] != ele[4][20];
    ele[1][20] != ele[4][21];
    ele[1][20] != ele[4][22];
    ele[1][20] != ele[4][23];
    ele[1][20] != ele[5][18];
    ele[1][20] != ele[5][19];
    ele[1][20] != ele[5][20];
    ele[1][20] != ele[5][21];
    ele[1][20] != ele[5][22];
    ele[1][20] != ele[5][23];
    ele[1][20] != ele[6][20];
    ele[1][20] != ele[7][20];
    ele[1][20] != ele[8][20];
    ele[1][20] != ele[9][20];
    ele[1][21] != ele[1][22];
    ele[1][21] != ele[1][23];
    ele[1][21] != ele[1][24];
    ele[1][21] != ele[1][25];
    ele[1][21] != ele[1][26];
    ele[1][21] != ele[1][27];
    ele[1][21] != ele[1][28];
    ele[1][21] != ele[1][29];
    ele[1][21] != ele[1][30];
    ele[1][21] != ele[1][31];
    ele[1][21] != ele[1][32];
    ele[1][21] != ele[1][33];
    ele[1][21] != ele[1][34];
    ele[1][21] != ele[1][35];
    ele[1][21] != ele[10][21];
    ele[1][21] != ele[11][21];
    ele[1][21] != ele[12][21];
    ele[1][21] != ele[13][21];
    ele[1][21] != ele[14][21];
    ele[1][21] != ele[15][21];
    ele[1][21] != ele[16][21];
    ele[1][21] != ele[17][21];
    ele[1][21] != ele[18][21];
    ele[1][21] != ele[19][21];
    ele[1][21] != ele[2][18];
    ele[1][21] != ele[2][19];
    ele[1][21] != ele[2][20];
    ele[1][21] != ele[2][21];
    ele[1][21] != ele[2][22];
    ele[1][21] != ele[2][23];
    ele[1][21] != ele[20][21];
    ele[1][21] != ele[21][21];
    ele[1][21] != ele[22][21];
    ele[1][21] != ele[23][21];
    ele[1][21] != ele[24][21];
    ele[1][21] != ele[25][21];
    ele[1][21] != ele[26][21];
    ele[1][21] != ele[27][21];
    ele[1][21] != ele[28][21];
    ele[1][21] != ele[29][21];
    ele[1][21] != ele[3][18];
    ele[1][21] != ele[3][19];
    ele[1][21] != ele[3][20];
    ele[1][21] != ele[3][21];
    ele[1][21] != ele[3][22];
    ele[1][21] != ele[3][23];
    ele[1][21] != ele[30][21];
    ele[1][21] != ele[31][21];
    ele[1][21] != ele[32][21];
    ele[1][21] != ele[33][21];
    ele[1][21] != ele[34][21];
    ele[1][21] != ele[35][21];
    ele[1][21] != ele[4][18];
    ele[1][21] != ele[4][19];
    ele[1][21] != ele[4][20];
    ele[1][21] != ele[4][21];
    ele[1][21] != ele[4][22];
    ele[1][21] != ele[4][23];
    ele[1][21] != ele[5][18];
    ele[1][21] != ele[5][19];
    ele[1][21] != ele[5][20];
    ele[1][21] != ele[5][21];
    ele[1][21] != ele[5][22];
    ele[1][21] != ele[5][23];
    ele[1][21] != ele[6][21];
    ele[1][21] != ele[7][21];
    ele[1][21] != ele[8][21];
    ele[1][21] != ele[9][21];
    ele[1][22] != ele[1][23];
    ele[1][22] != ele[1][24];
    ele[1][22] != ele[1][25];
    ele[1][22] != ele[1][26];
    ele[1][22] != ele[1][27];
    ele[1][22] != ele[1][28];
    ele[1][22] != ele[1][29];
    ele[1][22] != ele[1][30];
    ele[1][22] != ele[1][31];
    ele[1][22] != ele[1][32];
    ele[1][22] != ele[1][33];
    ele[1][22] != ele[1][34];
    ele[1][22] != ele[1][35];
    ele[1][22] != ele[10][22];
    ele[1][22] != ele[11][22];
    ele[1][22] != ele[12][22];
    ele[1][22] != ele[13][22];
    ele[1][22] != ele[14][22];
    ele[1][22] != ele[15][22];
    ele[1][22] != ele[16][22];
    ele[1][22] != ele[17][22];
    ele[1][22] != ele[18][22];
    ele[1][22] != ele[19][22];
    ele[1][22] != ele[2][18];
    ele[1][22] != ele[2][19];
    ele[1][22] != ele[2][20];
    ele[1][22] != ele[2][21];
    ele[1][22] != ele[2][22];
    ele[1][22] != ele[2][23];
    ele[1][22] != ele[20][22];
    ele[1][22] != ele[21][22];
    ele[1][22] != ele[22][22];
    ele[1][22] != ele[23][22];
    ele[1][22] != ele[24][22];
    ele[1][22] != ele[25][22];
    ele[1][22] != ele[26][22];
    ele[1][22] != ele[27][22];
    ele[1][22] != ele[28][22];
    ele[1][22] != ele[29][22];
    ele[1][22] != ele[3][18];
    ele[1][22] != ele[3][19];
    ele[1][22] != ele[3][20];
    ele[1][22] != ele[3][21];
    ele[1][22] != ele[3][22];
    ele[1][22] != ele[3][23];
    ele[1][22] != ele[30][22];
    ele[1][22] != ele[31][22];
    ele[1][22] != ele[32][22];
    ele[1][22] != ele[33][22];
    ele[1][22] != ele[34][22];
    ele[1][22] != ele[35][22];
    ele[1][22] != ele[4][18];
    ele[1][22] != ele[4][19];
    ele[1][22] != ele[4][20];
    ele[1][22] != ele[4][21];
    ele[1][22] != ele[4][22];
    ele[1][22] != ele[4][23];
    ele[1][22] != ele[5][18];
    ele[1][22] != ele[5][19];
    ele[1][22] != ele[5][20];
    ele[1][22] != ele[5][21];
    ele[1][22] != ele[5][22];
    ele[1][22] != ele[5][23];
    ele[1][22] != ele[6][22];
    ele[1][22] != ele[7][22];
    ele[1][22] != ele[8][22];
    ele[1][22] != ele[9][22];
    ele[1][23] != ele[1][24];
    ele[1][23] != ele[1][25];
    ele[1][23] != ele[1][26];
    ele[1][23] != ele[1][27];
    ele[1][23] != ele[1][28];
    ele[1][23] != ele[1][29];
    ele[1][23] != ele[1][30];
    ele[1][23] != ele[1][31];
    ele[1][23] != ele[1][32];
    ele[1][23] != ele[1][33];
    ele[1][23] != ele[1][34];
    ele[1][23] != ele[1][35];
    ele[1][23] != ele[10][23];
    ele[1][23] != ele[11][23];
    ele[1][23] != ele[12][23];
    ele[1][23] != ele[13][23];
    ele[1][23] != ele[14][23];
    ele[1][23] != ele[15][23];
    ele[1][23] != ele[16][23];
    ele[1][23] != ele[17][23];
    ele[1][23] != ele[18][23];
    ele[1][23] != ele[19][23];
    ele[1][23] != ele[2][18];
    ele[1][23] != ele[2][19];
    ele[1][23] != ele[2][20];
    ele[1][23] != ele[2][21];
    ele[1][23] != ele[2][22];
    ele[1][23] != ele[2][23];
    ele[1][23] != ele[20][23];
    ele[1][23] != ele[21][23];
    ele[1][23] != ele[22][23];
    ele[1][23] != ele[23][23];
    ele[1][23] != ele[24][23];
    ele[1][23] != ele[25][23];
    ele[1][23] != ele[26][23];
    ele[1][23] != ele[27][23];
    ele[1][23] != ele[28][23];
    ele[1][23] != ele[29][23];
    ele[1][23] != ele[3][18];
    ele[1][23] != ele[3][19];
    ele[1][23] != ele[3][20];
    ele[1][23] != ele[3][21];
    ele[1][23] != ele[3][22];
    ele[1][23] != ele[3][23];
    ele[1][23] != ele[30][23];
    ele[1][23] != ele[31][23];
    ele[1][23] != ele[32][23];
    ele[1][23] != ele[33][23];
    ele[1][23] != ele[34][23];
    ele[1][23] != ele[35][23];
    ele[1][23] != ele[4][18];
    ele[1][23] != ele[4][19];
    ele[1][23] != ele[4][20];
    ele[1][23] != ele[4][21];
    ele[1][23] != ele[4][22];
    ele[1][23] != ele[4][23];
    ele[1][23] != ele[5][18];
    ele[1][23] != ele[5][19];
    ele[1][23] != ele[5][20];
    ele[1][23] != ele[5][21];
    ele[1][23] != ele[5][22];
    ele[1][23] != ele[5][23];
    ele[1][23] != ele[6][23];
    ele[1][23] != ele[7][23];
    ele[1][23] != ele[8][23];
    ele[1][23] != ele[9][23];
    ele[1][24] != ele[1][25];
    ele[1][24] != ele[1][26];
    ele[1][24] != ele[1][27];
    ele[1][24] != ele[1][28];
    ele[1][24] != ele[1][29];
    ele[1][24] != ele[1][30];
    ele[1][24] != ele[1][31];
    ele[1][24] != ele[1][32];
    ele[1][24] != ele[1][33];
    ele[1][24] != ele[1][34];
    ele[1][24] != ele[1][35];
    ele[1][24] != ele[10][24];
    ele[1][24] != ele[11][24];
    ele[1][24] != ele[12][24];
    ele[1][24] != ele[13][24];
    ele[1][24] != ele[14][24];
    ele[1][24] != ele[15][24];
    ele[1][24] != ele[16][24];
    ele[1][24] != ele[17][24];
    ele[1][24] != ele[18][24];
    ele[1][24] != ele[19][24];
    ele[1][24] != ele[2][24];
    ele[1][24] != ele[2][25];
    ele[1][24] != ele[2][26];
    ele[1][24] != ele[2][27];
    ele[1][24] != ele[2][28];
    ele[1][24] != ele[2][29];
    ele[1][24] != ele[20][24];
    ele[1][24] != ele[21][24];
    ele[1][24] != ele[22][24];
    ele[1][24] != ele[23][24];
    ele[1][24] != ele[24][24];
    ele[1][24] != ele[25][24];
    ele[1][24] != ele[26][24];
    ele[1][24] != ele[27][24];
    ele[1][24] != ele[28][24];
    ele[1][24] != ele[29][24];
    ele[1][24] != ele[3][24];
    ele[1][24] != ele[3][25];
    ele[1][24] != ele[3][26];
    ele[1][24] != ele[3][27];
    ele[1][24] != ele[3][28];
    ele[1][24] != ele[3][29];
    ele[1][24] != ele[30][24];
    ele[1][24] != ele[31][24];
    ele[1][24] != ele[32][24];
    ele[1][24] != ele[33][24];
    ele[1][24] != ele[34][24];
    ele[1][24] != ele[35][24];
    ele[1][24] != ele[4][24];
    ele[1][24] != ele[4][25];
    ele[1][24] != ele[4][26];
    ele[1][24] != ele[4][27];
    ele[1][24] != ele[4][28];
    ele[1][24] != ele[4][29];
    ele[1][24] != ele[5][24];
    ele[1][24] != ele[5][25];
    ele[1][24] != ele[5][26];
    ele[1][24] != ele[5][27];
    ele[1][24] != ele[5][28];
    ele[1][24] != ele[5][29];
    ele[1][24] != ele[6][24];
    ele[1][24] != ele[7][24];
    ele[1][24] != ele[8][24];
    ele[1][24] != ele[9][24];
    ele[1][25] != ele[1][26];
    ele[1][25] != ele[1][27];
    ele[1][25] != ele[1][28];
    ele[1][25] != ele[1][29];
    ele[1][25] != ele[1][30];
    ele[1][25] != ele[1][31];
    ele[1][25] != ele[1][32];
    ele[1][25] != ele[1][33];
    ele[1][25] != ele[1][34];
    ele[1][25] != ele[1][35];
    ele[1][25] != ele[10][25];
    ele[1][25] != ele[11][25];
    ele[1][25] != ele[12][25];
    ele[1][25] != ele[13][25];
    ele[1][25] != ele[14][25];
    ele[1][25] != ele[15][25];
    ele[1][25] != ele[16][25];
    ele[1][25] != ele[17][25];
    ele[1][25] != ele[18][25];
    ele[1][25] != ele[19][25];
    ele[1][25] != ele[2][24];
    ele[1][25] != ele[2][25];
    ele[1][25] != ele[2][26];
    ele[1][25] != ele[2][27];
    ele[1][25] != ele[2][28];
    ele[1][25] != ele[2][29];
    ele[1][25] != ele[20][25];
    ele[1][25] != ele[21][25];
    ele[1][25] != ele[22][25];
    ele[1][25] != ele[23][25];
    ele[1][25] != ele[24][25];
    ele[1][25] != ele[25][25];
    ele[1][25] != ele[26][25];
    ele[1][25] != ele[27][25];
    ele[1][25] != ele[28][25];
    ele[1][25] != ele[29][25];
    ele[1][25] != ele[3][24];
    ele[1][25] != ele[3][25];
    ele[1][25] != ele[3][26];
    ele[1][25] != ele[3][27];
    ele[1][25] != ele[3][28];
    ele[1][25] != ele[3][29];
    ele[1][25] != ele[30][25];
    ele[1][25] != ele[31][25];
    ele[1][25] != ele[32][25];
    ele[1][25] != ele[33][25];
    ele[1][25] != ele[34][25];
    ele[1][25] != ele[35][25];
    ele[1][25] != ele[4][24];
    ele[1][25] != ele[4][25];
    ele[1][25] != ele[4][26];
    ele[1][25] != ele[4][27];
    ele[1][25] != ele[4][28];
    ele[1][25] != ele[4][29];
    ele[1][25] != ele[5][24];
    ele[1][25] != ele[5][25];
    ele[1][25] != ele[5][26];
    ele[1][25] != ele[5][27];
    ele[1][25] != ele[5][28];
    ele[1][25] != ele[5][29];
    ele[1][25] != ele[6][25];
    ele[1][25] != ele[7][25];
    ele[1][25] != ele[8][25];
    ele[1][25] != ele[9][25];
    ele[1][26] != ele[1][27];
    ele[1][26] != ele[1][28];
    ele[1][26] != ele[1][29];
    ele[1][26] != ele[1][30];
    ele[1][26] != ele[1][31];
    ele[1][26] != ele[1][32];
    ele[1][26] != ele[1][33];
    ele[1][26] != ele[1][34];
    ele[1][26] != ele[1][35];
    ele[1][26] != ele[10][26];
    ele[1][26] != ele[11][26];
    ele[1][26] != ele[12][26];
    ele[1][26] != ele[13][26];
    ele[1][26] != ele[14][26];
    ele[1][26] != ele[15][26];
    ele[1][26] != ele[16][26];
    ele[1][26] != ele[17][26];
    ele[1][26] != ele[18][26];
    ele[1][26] != ele[19][26];
    ele[1][26] != ele[2][24];
    ele[1][26] != ele[2][25];
    ele[1][26] != ele[2][26];
    ele[1][26] != ele[2][27];
    ele[1][26] != ele[2][28];
    ele[1][26] != ele[2][29];
    ele[1][26] != ele[20][26];
    ele[1][26] != ele[21][26];
    ele[1][26] != ele[22][26];
    ele[1][26] != ele[23][26];
    ele[1][26] != ele[24][26];
    ele[1][26] != ele[25][26];
    ele[1][26] != ele[26][26];
    ele[1][26] != ele[27][26];
    ele[1][26] != ele[28][26];
    ele[1][26] != ele[29][26];
    ele[1][26] != ele[3][24];
    ele[1][26] != ele[3][25];
    ele[1][26] != ele[3][26];
    ele[1][26] != ele[3][27];
    ele[1][26] != ele[3][28];
    ele[1][26] != ele[3][29];
    ele[1][26] != ele[30][26];
    ele[1][26] != ele[31][26];
    ele[1][26] != ele[32][26];
    ele[1][26] != ele[33][26];
    ele[1][26] != ele[34][26];
    ele[1][26] != ele[35][26];
    ele[1][26] != ele[4][24];
    ele[1][26] != ele[4][25];
    ele[1][26] != ele[4][26];
    ele[1][26] != ele[4][27];
    ele[1][26] != ele[4][28];
    ele[1][26] != ele[4][29];
    ele[1][26] != ele[5][24];
    ele[1][26] != ele[5][25];
    ele[1][26] != ele[5][26];
    ele[1][26] != ele[5][27];
    ele[1][26] != ele[5][28];
    ele[1][26] != ele[5][29];
    ele[1][26] != ele[6][26];
    ele[1][26] != ele[7][26];
    ele[1][26] != ele[8][26];
    ele[1][26] != ele[9][26];
    ele[1][27] != ele[1][28];
    ele[1][27] != ele[1][29];
    ele[1][27] != ele[1][30];
    ele[1][27] != ele[1][31];
    ele[1][27] != ele[1][32];
    ele[1][27] != ele[1][33];
    ele[1][27] != ele[1][34];
    ele[1][27] != ele[1][35];
    ele[1][27] != ele[10][27];
    ele[1][27] != ele[11][27];
    ele[1][27] != ele[12][27];
    ele[1][27] != ele[13][27];
    ele[1][27] != ele[14][27];
    ele[1][27] != ele[15][27];
    ele[1][27] != ele[16][27];
    ele[1][27] != ele[17][27];
    ele[1][27] != ele[18][27];
    ele[1][27] != ele[19][27];
    ele[1][27] != ele[2][24];
    ele[1][27] != ele[2][25];
    ele[1][27] != ele[2][26];
    ele[1][27] != ele[2][27];
    ele[1][27] != ele[2][28];
    ele[1][27] != ele[2][29];
    ele[1][27] != ele[20][27];
    ele[1][27] != ele[21][27];
    ele[1][27] != ele[22][27];
    ele[1][27] != ele[23][27];
    ele[1][27] != ele[24][27];
    ele[1][27] != ele[25][27];
    ele[1][27] != ele[26][27];
    ele[1][27] != ele[27][27];
    ele[1][27] != ele[28][27];
    ele[1][27] != ele[29][27];
    ele[1][27] != ele[3][24];
    ele[1][27] != ele[3][25];
    ele[1][27] != ele[3][26];
    ele[1][27] != ele[3][27];
    ele[1][27] != ele[3][28];
    ele[1][27] != ele[3][29];
    ele[1][27] != ele[30][27];
    ele[1][27] != ele[31][27];
    ele[1][27] != ele[32][27];
    ele[1][27] != ele[33][27];
    ele[1][27] != ele[34][27];
    ele[1][27] != ele[35][27];
    ele[1][27] != ele[4][24];
    ele[1][27] != ele[4][25];
    ele[1][27] != ele[4][26];
    ele[1][27] != ele[4][27];
    ele[1][27] != ele[4][28];
    ele[1][27] != ele[4][29];
    ele[1][27] != ele[5][24];
    ele[1][27] != ele[5][25];
    ele[1][27] != ele[5][26];
    ele[1][27] != ele[5][27];
    ele[1][27] != ele[5][28];
    ele[1][27] != ele[5][29];
    ele[1][27] != ele[6][27];
    ele[1][27] != ele[7][27];
    ele[1][27] != ele[8][27];
    ele[1][27] != ele[9][27];
    ele[1][28] != ele[1][29];
    ele[1][28] != ele[1][30];
    ele[1][28] != ele[1][31];
    ele[1][28] != ele[1][32];
    ele[1][28] != ele[1][33];
    ele[1][28] != ele[1][34];
    ele[1][28] != ele[1][35];
    ele[1][28] != ele[10][28];
    ele[1][28] != ele[11][28];
    ele[1][28] != ele[12][28];
    ele[1][28] != ele[13][28];
    ele[1][28] != ele[14][28];
    ele[1][28] != ele[15][28];
    ele[1][28] != ele[16][28];
    ele[1][28] != ele[17][28];
    ele[1][28] != ele[18][28];
    ele[1][28] != ele[19][28];
    ele[1][28] != ele[2][24];
    ele[1][28] != ele[2][25];
    ele[1][28] != ele[2][26];
    ele[1][28] != ele[2][27];
    ele[1][28] != ele[2][28];
    ele[1][28] != ele[2][29];
    ele[1][28] != ele[20][28];
    ele[1][28] != ele[21][28];
    ele[1][28] != ele[22][28];
    ele[1][28] != ele[23][28];
    ele[1][28] != ele[24][28];
    ele[1][28] != ele[25][28];
    ele[1][28] != ele[26][28];
    ele[1][28] != ele[27][28];
    ele[1][28] != ele[28][28];
    ele[1][28] != ele[29][28];
    ele[1][28] != ele[3][24];
    ele[1][28] != ele[3][25];
    ele[1][28] != ele[3][26];
    ele[1][28] != ele[3][27];
    ele[1][28] != ele[3][28];
    ele[1][28] != ele[3][29];
    ele[1][28] != ele[30][28];
    ele[1][28] != ele[31][28];
    ele[1][28] != ele[32][28];
    ele[1][28] != ele[33][28];
    ele[1][28] != ele[34][28];
    ele[1][28] != ele[35][28];
    ele[1][28] != ele[4][24];
    ele[1][28] != ele[4][25];
    ele[1][28] != ele[4][26];
    ele[1][28] != ele[4][27];
    ele[1][28] != ele[4][28];
    ele[1][28] != ele[4][29];
    ele[1][28] != ele[5][24];
    ele[1][28] != ele[5][25];
    ele[1][28] != ele[5][26];
    ele[1][28] != ele[5][27];
    ele[1][28] != ele[5][28];
    ele[1][28] != ele[5][29];
    ele[1][28] != ele[6][28];
    ele[1][28] != ele[7][28];
    ele[1][28] != ele[8][28];
    ele[1][28] != ele[9][28];
    ele[1][29] != ele[1][30];
    ele[1][29] != ele[1][31];
    ele[1][29] != ele[1][32];
    ele[1][29] != ele[1][33];
    ele[1][29] != ele[1][34];
    ele[1][29] != ele[1][35];
    ele[1][29] != ele[10][29];
    ele[1][29] != ele[11][29];
    ele[1][29] != ele[12][29];
    ele[1][29] != ele[13][29];
    ele[1][29] != ele[14][29];
    ele[1][29] != ele[15][29];
    ele[1][29] != ele[16][29];
    ele[1][29] != ele[17][29];
    ele[1][29] != ele[18][29];
    ele[1][29] != ele[19][29];
    ele[1][29] != ele[2][24];
    ele[1][29] != ele[2][25];
    ele[1][29] != ele[2][26];
    ele[1][29] != ele[2][27];
    ele[1][29] != ele[2][28];
    ele[1][29] != ele[2][29];
    ele[1][29] != ele[20][29];
    ele[1][29] != ele[21][29];
    ele[1][29] != ele[22][29];
    ele[1][29] != ele[23][29];
    ele[1][29] != ele[24][29];
    ele[1][29] != ele[25][29];
    ele[1][29] != ele[26][29];
    ele[1][29] != ele[27][29];
    ele[1][29] != ele[28][29];
    ele[1][29] != ele[29][29];
    ele[1][29] != ele[3][24];
    ele[1][29] != ele[3][25];
    ele[1][29] != ele[3][26];
    ele[1][29] != ele[3][27];
    ele[1][29] != ele[3][28];
    ele[1][29] != ele[3][29];
    ele[1][29] != ele[30][29];
    ele[1][29] != ele[31][29];
    ele[1][29] != ele[32][29];
    ele[1][29] != ele[33][29];
    ele[1][29] != ele[34][29];
    ele[1][29] != ele[35][29];
    ele[1][29] != ele[4][24];
    ele[1][29] != ele[4][25];
    ele[1][29] != ele[4][26];
    ele[1][29] != ele[4][27];
    ele[1][29] != ele[4][28];
    ele[1][29] != ele[4][29];
    ele[1][29] != ele[5][24];
    ele[1][29] != ele[5][25];
    ele[1][29] != ele[5][26];
    ele[1][29] != ele[5][27];
    ele[1][29] != ele[5][28];
    ele[1][29] != ele[5][29];
    ele[1][29] != ele[6][29];
    ele[1][29] != ele[7][29];
    ele[1][29] != ele[8][29];
    ele[1][29] != ele[9][29];
    ele[1][3] != ele[1][10];
    ele[1][3] != ele[1][11];
    ele[1][3] != ele[1][12];
    ele[1][3] != ele[1][13];
    ele[1][3] != ele[1][14];
    ele[1][3] != ele[1][15];
    ele[1][3] != ele[1][16];
    ele[1][3] != ele[1][17];
    ele[1][3] != ele[1][18];
    ele[1][3] != ele[1][19];
    ele[1][3] != ele[1][20];
    ele[1][3] != ele[1][21];
    ele[1][3] != ele[1][22];
    ele[1][3] != ele[1][23];
    ele[1][3] != ele[1][24];
    ele[1][3] != ele[1][25];
    ele[1][3] != ele[1][26];
    ele[1][3] != ele[1][27];
    ele[1][3] != ele[1][28];
    ele[1][3] != ele[1][29];
    ele[1][3] != ele[1][30];
    ele[1][3] != ele[1][31];
    ele[1][3] != ele[1][32];
    ele[1][3] != ele[1][33];
    ele[1][3] != ele[1][34];
    ele[1][3] != ele[1][35];
    ele[1][3] != ele[1][4];
    ele[1][3] != ele[1][5];
    ele[1][3] != ele[1][6];
    ele[1][3] != ele[1][7];
    ele[1][3] != ele[1][8];
    ele[1][3] != ele[1][9];
    ele[1][3] != ele[10][3];
    ele[1][3] != ele[11][3];
    ele[1][3] != ele[12][3];
    ele[1][3] != ele[13][3];
    ele[1][3] != ele[14][3];
    ele[1][3] != ele[15][3];
    ele[1][3] != ele[16][3];
    ele[1][3] != ele[17][3];
    ele[1][3] != ele[18][3];
    ele[1][3] != ele[19][3];
    ele[1][3] != ele[2][0];
    ele[1][3] != ele[2][1];
    ele[1][3] != ele[2][2];
    ele[1][3] != ele[2][3];
    ele[1][3] != ele[2][4];
    ele[1][3] != ele[2][5];
    ele[1][3] != ele[20][3];
    ele[1][3] != ele[21][3];
    ele[1][3] != ele[22][3];
    ele[1][3] != ele[23][3];
    ele[1][3] != ele[24][3];
    ele[1][3] != ele[25][3];
    ele[1][3] != ele[26][3];
    ele[1][3] != ele[27][3];
    ele[1][3] != ele[28][3];
    ele[1][3] != ele[29][3];
    ele[1][3] != ele[3][0];
    ele[1][3] != ele[3][1];
    ele[1][3] != ele[3][2];
    ele[1][3] != ele[3][3];
    ele[1][3] != ele[3][4];
    ele[1][3] != ele[3][5];
    ele[1][3] != ele[30][3];
    ele[1][3] != ele[31][3];
    ele[1][3] != ele[32][3];
    ele[1][3] != ele[33][3];
    ele[1][3] != ele[34][3];
    ele[1][3] != ele[35][3];
    ele[1][3] != ele[4][0];
    ele[1][3] != ele[4][1];
    ele[1][3] != ele[4][2];
    ele[1][3] != ele[4][3];
    ele[1][3] != ele[4][4];
    ele[1][3] != ele[4][5];
    ele[1][3] != ele[5][0];
    ele[1][3] != ele[5][1];
    ele[1][3] != ele[5][2];
    ele[1][3] != ele[5][3];
    ele[1][3] != ele[5][4];
    ele[1][3] != ele[5][5];
    ele[1][3] != ele[6][3];
    ele[1][3] != ele[7][3];
    ele[1][3] != ele[8][3];
    ele[1][3] != ele[9][3];
    ele[1][30] != ele[1][31];
    ele[1][30] != ele[1][32];
    ele[1][30] != ele[1][33];
    ele[1][30] != ele[1][34];
    ele[1][30] != ele[1][35];
    ele[1][30] != ele[10][30];
    ele[1][30] != ele[11][30];
    ele[1][30] != ele[12][30];
    ele[1][30] != ele[13][30];
    ele[1][30] != ele[14][30];
    ele[1][30] != ele[15][30];
    ele[1][30] != ele[16][30];
    ele[1][30] != ele[17][30];
    ele[1][30] != ele[18][30];
    ele[1][30] != ele[19][30];
    ele[1][30] != ele[2][30];
    ele[1][30] != ele[2][31];
    ele[1][30] != ele[2][32];
    ele[1][30] != ele[2][33];
    ele[1][30] != ele[2][34];
    ele[1][30] != ele[2][35];
    ele[1][30] != ele[20][30];
    ele[1][30] != ele[21][30];
    ele[1][30] != ele[22][30];
    ele[1][30] != ele[23][30];
    ele[1][30] != ele[24][30];
    ele[1][30] != ele[25][30];
    ele[1][30] != ele[26][30];
    ele[1][30] != ele[27][30];
    ele[1][30] != ele[28][30];
    ele[1][30] != ele[29][30];
    ele[1][30] != ele[3][30];
    ele[1][30] != ele[3][31];
    ele[1][30] != ele[3][32];
    ele[1][30] != ele[3][33];
    ele[1][30] != ele[3][34];
    ele[1][30] != ele[3][35];
    ele[1][30] != ele[30][30];
    ele[1][30] != ele[31][30];
    ele[1][30] != ele[32][30];
    ele[1][30] != ele[33][30];
    ele[1][30] != ele[34][30];
    ele[1][30] != ele[35][30];
    ele[1][30] != ele[4][30];
    ele[1][30] != ele[4][31];
    ele[1][30] != ele[4][32];
    ele[1][30] != ele[4][33];
    ele[1][30] != ele[4][34];
    ele[1][30] != ele[4][35];
    ele[1][30] != ele[5][30];
    ele[1][30] != ele[5][31];
    ele[1][30] != ele[5][32];
    ele[1][30] != ele[5][33];
    ele[1][30] != ele[5][34];
    ele[1][30] != ele[5][35];
    ele[1][30] != ele[6][30];
    ele[1][30] != ele[7][30];
    ele[1][30] != ele[8][30];
    ele[1][30] != ele[9][30];
    ele[1][31] != ele[1][32];
    ele[1][31] != ele[1][33];
    ele[1][31] != ele[1][34];
    ele[1][31] != ele[1][35];
    ele[1][31] != ele[10][31];
    ele[1][31] != ele[11][31];
    ele[1][31] != ele[12][31];
    ele[1][31] != ele[13][31];
    ele[1][31] != ele[14][31];
    ele[1][31] != ele[15][31];
    ele[1][31] != ele[16][31];
    ele[1][31] != ele[17][31];
    ele[1][31] != ele[18][31];
    ele[1][31] != ele[19][31];
    ele[1][31] != ele[2][30];
    ele[1][31] != ele[2][31];
    ele[1][31] != ele[2][32];
    ele[1][31] != ele[2][33];
    ele[1][31] != ele[2][34];
    ele[1][31] != ele[2][35];
    ele[1][31] != ele[20][31];
    ele[1][31] != ele[21][31];
    ele[1][31] != ele[22][31];
    ele[1][31] != ele[23][31];
    ele[1][31] != ele[24][31];
    ele[1][31] != ele[25][31];
    ele[1][31] != ele[26][31];
    ele[1][31] != ele[27][31];
    ele[1][31] != ele[28][31];
    ele[1][31] != ele[29][31];
    ele[1][31] != ele[3][30];
    ele[1][31] != ele[3][31];
    ele[1][31] != ele[3][32];
    ele[1][31] != ele[3][33];
    ele[1][31] != ele[3][34];
    ele[1][31] != ele[3][35];
    ele[1][31] != ele[30][31];
    ele[1][31] != ele[31][31];
    ele[1][31] != ele[32][31];
    ele[1][31] != ele[33][31];
    ele[1][31] != ele[34][31];
    ele[1][31] != ele[35][31];
    ele[1][31] != ele[4][30];
    ele[1][31] != ele[4][31];
    ele[1][31] != ele[4][32];
    ele[1][31] != ele[4][33];
    ele[1][31] != ele[4][34];
    ele[1][31] != ele[4][35];
    ele[1][31] != ele[5][30];
    ele[1][31] != ele[5][31];
    ele[1][31] != ele[5][32];
    ele[1][31] != ele[5][33];
    ele[1][31] != ele[5][34];
    ele[1][31] != ele[5][35];
    ele[1][31] != ele[6][31];
    ele[1][31] != ele[7][31];
    ele[1][31] != ele[8][31];
    ele[1][31] != ele[9][31];
    ele[1][32] != ele[1][33];
    ele[1][32] != ele[1][34];
    ele[1][32] != ele[1][35];
    ele[1][32] != ele[10][32];
    ele[1][32] != ele[11][32];
    ele[1][32] != ele[12][32];
    ele[1][32] != ele[13][32];
    ele[1][32] != ele[14][32];
    ele[1][32] != ele[15][32];
    ele[1][32] != ele[16][32];
    ele[1][32] != ele[17][32];
    ele[1][32] != ele[18][32];
    ele[1][32] != ele[19][32];
    ele[1][32] != ele[2][30];
    ele[1][32] != ele[2][31];
    ele[1][32] != ele[2][32];
    ele[1][32] != ele[2][33];
    ele[1][32] != ele[2][34];
    ele[1][32] != ele[2][35];
    ele[1][32] != ele[20][32];
    ele[1][32] != ele[21][32];
    ele[1][32] != ele[22][32];
    ele[1][32] != ele[23][32];
    ele[1][32] != ele[24][32];
    ele[1][32] != ele[25][32];
    ele[1][32] != ele[26][32];
    ele[1][32] != ele[27][32];
    ele[1][32] != ele[28][32];
    ele[1][32] != ele[29][32];
    ele[1][32] != ele[3][30];
    ele[1][32] != ele[3][31];
    ele[1][32] != ele[3][32];
    ele[1][32] != ele[3][33];
    ele[1][32] != ele[3][34];
    ele[1][32] != ele[3][35];
    ele[1][32] != ele[30][32];
    ele[1][32] != ele[31][32];
    ele[1][32] != ele[32][32];
    ele[1][32] != ele[33][32];
    ele[1][32] != ele[34][32];
    ele[1][32] != ele[35][32];
    ele[1][32] != ele[4][30];
    ele[1][32] != ele[4][31];
    ele[1][32] != ele[4][32];
    ele[1][32] != ele[4][33];
    ele[1][32] != ele[4][34];
    ele[1][32] != ele[4][35];
    ele[1][32] != ele[5][30];
    ele[1][32] != ele[5][31];
    ele[1][32] != ele[5][32];
    ele[1][32] != ele[5][33];
    ele[1][32] != ele[5][34];
    ele[1][32] != ele[5][35];
    ele[1][32] != ele[6][32];
    ele[1][32] != ele[7][32];
    ele[1][32] != ele[8][32];
    ele[1][32] != ele[9][32];
    ele[1][33] != ele[1][34];
    ele[1][33] != ele[1][35];
    ele[1][33] != ele[10][33];
    ele[1][33] != ele[11][33];
    ele[1][33] != ele[12][33];
    ele[1][33] != ele[13][33];
    ele[1][33] != ele[14][33];
    ele[1][33] != ele[15][33];
    ele[1][33] != ele[16][33];
    ele[1][33] != ele[17][33];
    ele[1][33] != ele[18][33];
    ele[1][33] != ele[19][33];
    ele[1][33] != ele[2][30];
    ele[1][33] != ele[2][31];
    ele[1][33] != ele[2][32];
    ele[1][33] != ele[2][33];
    ele[1][33] != ele[2][34];
    ele[1][33] != ele[2][35];
    ele[1][33] != ele[20][33];
    ele[1][33] != ele[21][33];
    ele[1][33] != ele[22][33];
    ele[1][33] != ele[23][33];
    ele[1][33] != ele[24][33];
    ele[1][33] != ele[25][33];
    ele[1][33] != ele[26][33];
    ele[1][33] != ele[27][33];
    ele[1][33] != ele[28][33];
    ele[1][33] != ele[29][33];
    ele[1][33] != ele[3][30];
    ele[1][33] != ele[3][31];
    ele[1][33] != ele[3][32];
    ele[1][33] != ele[3][33];
    ele[1][33] != ele[3][34];
    ele[1][33] != ele[3][35];
    ele[1][33] != ele[30][33];
    ele[1][33] != ele[31][33];
    ele[1][33] != ele[32][33];
    ele[1][33] != ele[33][33];
    ele[1][33] != ele[34][33];
    ele[1][33] != ele[35][33];
    ele[1][33] != ele[4][30];
    ele[1][33] != ele[4][31];
    ele[1][33] != ele[4][32];
    ele[1][33] != ele[4][33];
    ele[1][33] != ele[4][34];
    ele[1][33] != ele[4][35];
    ele[1][33] != ele[5][30];
    ele[1][33] != ele[5][31];
    ele[1][33] != ele[5][32];
    ele[1][33] != ele[5][33];
    ele[1][33] != ele[5][34];
    ele[1][33] != ele[5][35];
    ele[1][33] != ele[6][33];
    ele[1][33] != ele[7][33];
    ele[1][33] != ele[8][33];
    ele[1][33] != ele[9][33];
    ele[1][34] != ele[1][35];
    ele[1][34] != ele[10][34];
    ele[1][34] != ele[11][34];
    ele[1][34] != ele[12][34];
    ele[1][34] != ele[13][34];
    ele[1][34] != ele[14][34];
    ele[1][34] != ele[15][34];
    ele[1][34] != ele[16][34];
    ele[1][34] != ele[17][34];
    ele[1][34] != ele[18][34];
    ele[1][34] != ele[19][34];
    ele[1][34] != ele[2][30];
    ele[1][34] != ele[2][31];
    ele[1][34] != ele[2][32];
    ele[1][34] != ele[2][33];
    ele[1][34] != ele[2][34];
    ele[1][34] != ele[2][35];
    ele[1][34] != ele[20][34];
    ele[1][34] != ele[21][34];
    ele[1][34] != ele[22][34];
    ele[1][34] != ele[23][34];
    ele[1][34] != ele[24][34];
    ele[1][34] != ele[25][34];
    ele[1][34] != ele[26][34];
    ele[1][34] != ele[27][34];
    ele[1][34] != ele[28][34];
    ele[1][34] != ele[29][34];
    ele[1][34] != ele[3][30];
    ele[1][34] != ele[3][31];
    ele[1][34] != ele[3][32];
    ele[1][34] != ele[3][33];
    ele[1][34] != ele[3][34];
    ele[1][34] != ele[3][35];
    ele[1][34] != ele[30][34];
    ele[1][34] != ele[31][34];
    ele[1][34] != ele[32][34];
    ele[1][34] != ele[33][34];
    ele[1][34] != ele[34][34];
    ele[1][34] != ele[35][34];
    ele[1][34] != ele[4][30];
    ele[1][34] != ele[4][31];
    ele[1][34] != ele[4][32];
    ele[1][34] != ele[4][33];
    ele[1][34] != ele[4][34];
    ele[1][34] != ele[4][35];
    ele[1][34] != ele[5][30];
    ele[1][34] != ele[5][31];
    ele[1][34] != ele[5][32];
    ele[1][34] != ele[5][33];
    ele[1][34] != ele[5][34];
    ele[1][34] != ele[5][35];
    ele[1][34] != ele[6][34];
    ele[1][34] != ele[7][34];
    ele[1][34] != ele[8][34];
    ele[1][34] != ele[9][34];
    ele[1][35] != ele[10][35];
    ele[1][35] != ele[11][35];
    ele[1][35] != ele[12][35];
    ele[1][35] != ele[13][35];
    ele[1][35] != ele[14][35];
    ele[1][35] != ele[15][35];
    ele[1][35] != ele[16][35];
    ele[1][35] != ele[17][35];
    ele[1][35] != ele[18][35];
    ele[1][35] != ele[19][35];
    ele[1][35] != ele[2][30];
    ele[1][35] != ele[2][31];
    ele[1][35] != ele[2][32];
    ele[1][35] != ele[2][33];
    ele[1][35] != ele[2][34];
    ele[1][35] != ele[2][35];
    ele[1][35] != ele[20][35];
    ele[1][35] != ele[21][35];
    ele[1][35] != ele[22][35];
    ele[1][35] != ele[23][35];
    ele[1][35] != ele[24][35];
    ele[1][35] != ele[25][35];
    ele[1][35] != ele[26][35];
    ele[1][35] != ele[27][35];
    ele[1][35] != ele[28][35];
    ele[1][35] != ele[29][35];
    ele[1][35] != ele[3][30];
    ele[1][35] != ele[3][31];
    ele[1][35] != ele[3][32];
    ele[1][35] != ele[3][33];
    ele[1][35] != ele[3][34];
    ele[1][35] != ele[3][35];
    ele[1][35] != ele[30][35];
    ele[1][35] != ele[31][35];
    ele[1][35] != ele[32][35];
    ele[1][35] != ele[33][35];
    ele[1][35] != ele[34][35];
    ele[1][35] != ele[35][35];
    ele[1][35] != ele[4][30];
    ele[1][35] != ele[4][31];
    ele[1][35] != ele[4][32];
    ele[1][35] != ele[4][33];
    ele[1][35] != ele[4][34];
    ele[1][35] != ele[4][35];
    ele[1][35] != ele[5][30];
    ele[1][35] != ele[5][31];
    ele[1][35] != ele[5][32];
    ele[1][35] != ele[5][33];
    ele[1][35] != ele[5][34];
    ele[1][35] != ele[5][35];
    ele[1][35] != ele[6][35];
    ele[1][35] != ele[7][35];
    ele[1][35] != ele[8][35];
    ele[1][35] != ele[9][35];
    ele[1][4] != ele[1][10];
    ele[1][4] != ele[1][11];
    ele[1][4] != ele[1][12];
    ele[1][4] != ele[1][13];
    ele[1][4] != ele[1][14];
    ele[1][4] != ele[1][15];
    ele[1][4] != ele[1][16];
    ele[1][4] != ele[1][17];
    ele[1][4] != ele[1][18];
    ele[1][4] != ele[1][19];
    ele[1][4] != ele[1][20];
    ele[1][4] != ele[1][21];
    ele[1][4] != ele[1][22];
    ele[1][4] != ele[1][23];
    ele[1][4] != ele[1][24];
    ele[1][4] != ele[1][25];
    ele[1][4] != ele[1][26];
    ele[1][4] != ele[1][27];
    ele[1][4] != ele[1][28];
    ele[1][4] != ele[1][29];
    ele[1][4] != ele[1][30];
    ele[1][4] != ele[1][31];
    ele[1][4] != ele[1][32];
    ele[1][4] != ele[1][33];
    ele[1][4] != ele[1][34];
    ele[1][4] != ele[1][35];
    ele[1][4] != ele[1][5];
    ele[1][4] != ele[1][6];
    ele[1][4] != ele[1][7];
    ele[1][4] != ele[1][8];
    ele[1][4] != ele[1][9];
    ele[1][4] != ele[10][4];
    ele[1][4] != ele[11][4];
    ele[1][4] != ele[12][4];
    ele[1][4] != ele[13][4];
    ele[1][4] != ele[14][4];
    ele[1][4] != ele[15][4];
    ele[1][4] != ele[16][4];
    ele[1][4] != ele[17][4];
    ele[1][4] != ele[18][4];
    ele[1][4] != ele[19][4];
    ele[1][4] != ele[2][0];
    ele[1][4] != ele[2][1];
    ele[1][4] != ele[2][2];
    ele[1][4] != ele[2][3];
    ele[1][4] != ele[2][4];
    ele[1][4] != ele[2][5];
    ele[1][4] != ele[20][4];
    ele[1][4] != ele[21][4];
    ele[1][4] != ele[22][4];
    ele[1][4] != ele[23][4];
    ele[1][4] != ele[24][4];
    ele[1][4] != ele[25][4];
    ele[1][4] != ele[26][4];
    ele[1][4] != ele[27][4];
    ele[1][4] != ele[28][4];
    ele[1][4] != ele[29][4];
    ele[1][4] != ele[3][0];
    ele[1][4] != ele[3][1];
    ele[1][4] != ele[3][2];
    ele[1][4] != ele[3][3];
    ele[1][4] != ele[3][4];
    ele[1][4] != ele[3][5];
    ele[1][4] != ele[30][4];
    ele[1][4] != ele[31][4];
    ele[1][4] != ele[32][4];
    ele[1][4] != ele[33][4];
    ele[1][4] != ele[34][4];
    ele[1][4] != ele[35][4];
    ele[1][4] != ele[4][0];
    ele[1][4] != ele[4][1];
    ele[1][4] != ele[4][2];
    ele[1][4] != ele[4][3];
    ele[1][4] != ele[4][4];
    ele[1][4] != ele[4][5];
    ele[1][4] != ele[5][0];
    ele[1][4] != ele[5][1];
    ele[1][4] != ele[5][2];
    ele[1][4] != ele[5][3];
    ele[1][4] != ele[5][4];
    ele[1][4] != ele[5][5];
    ele[1][4] != ele[6][4];
    ele[1][4] != ele[7][4];
    ele[1][4] != ele[8][4];
    ele[1][4] != ele[9][4];
    ele[1][5] != ele[1][10];
    ele[1][5] != ele[1][11];
    ele[1][5] != ele[1][12];
    ele[1][5] != ele[1][13];
    ele[1][5] != ele[1][14];
    ele[1][5] != ele[1][15];
    ele[1][5] != ele[1][16];
    ele[1][5] != ele[1][17];
    ele[1][5] != ele[1][18];
    ele[1][5] != ele[1][19];
    ele[1][5] != ele[1][20];
    ele[1][5] != ele[1][21];
    ele[1][5] != ele[1][22];
    ele[1][5] != ele[1][23];
    ele[1][5] != ele[1][24];
    ele[1][5] != ele[1][25];
    ele[1][5] != ele[1][26];
    ele[1][5] != ele[1][27];
    ele[1][5] != ele[1][28];
    ele[1][5] != ele[1][29];
    ele[1][5] != ele[1][30];
    ele[1][5] != ele[1][31];
    ele[1][5] != ele[1][32];
    ele[1][5] != ele[1][33];
    ele[1][5] != ele[1][34];
    ele[1][5] != ele[1][35];
    ele[1][5] != ele[1][6];
    ele[1][5] != ele[1][7];
    ele[1][5] != ele[1][8];
    ele[1][5] != ele[1][9];
    ele[1][5] != ele[10][5];
    ele[1][5] != ele[11][5];
    ele[1][5] != ele[12][5];
    ele[1][5] != ele[13][5];
    ele[1][5] != ele[14][5];
    ele[1][5] != ele[15][5];
    ele[1][5] != ele[16][5];
    ele[1][5] != ele[17][5];
    ele[1][5] != ele[18][5];
    ele[1][5] != ele[19][5];
    ele[1][5] != ele[2][0];
    ele[1][5] != ele[2][1];
    ele[1][5] != ele[2][2];
    ele[1][5] != ele[2][3];
    ele[1][5] != ele[2][4];
    ele[1][5] != ele[2][5];
    ele[1][5] != ele[20][5];
    ele[1][5] != ele[21][5];
    ele[1][5] != ele[22][5];
    ele[1][5] != ele[23][5];
    ele[1][5] != ele[24][5];
    ele[1][5] != ele[25][5];
    ele[1][5] != ele[26][5];
    ele[1][5] != ele[27][5];
    ele[1][5] != ele[28][5];
    ele[1][5] != ele[29][5];
    ele[1][5] != ele[3][0];
    ele[1][5] != ele[3][1];
    ele[1][5] != ele[3][2];
    ele[1][5] != ele[3][3];
    ele[1][5] != ele[3][4];
    ele[1][5] != ele[3][5];
    ele[1][5] != ele[30][5];
    ele[1][5] != ele[31][5];
    ele[1][5] != ele[32][5];
    ele[1][5] != ele[33][5];
    ele[1][5] != ele[34][5];
    ele[1][5] != ele[35][5];
    ele[1][5] != ele[4][0];
    ele[1][5] != ele[4][1];
    ele[1][5] != ele[4][2];
    ele[1][5] != ele[4][3];
    ele[1][5] != ele[4][4];
    ele[1][5] != ele[4][5];
    ele[1][5] != ele[5][0];
    ele[1][5] != ele[5][1];
    ele[1][5] != ele[5][2];
    ele[1][5] != ele[5][3];
    ele[1][5] != ele[5][4];
    ele[1][5] != ele[5][5];
    ele[1][5] != ele[6][5];
    ele[1][5] != ele[7][5];
    ele[1][5] != ele[8][5];
    ele[1][5] != ele[9][5];
    ele[1][6] != ele[1][10];
    ele[1][6] != ele[1][11];
    ele[1][6] != ele[1][12];
    ele[1][6] != ele[1][13];
    ele[1][6] != ele[1][14];
    ele[1][6] != ele[1][15];
    ele[1][6] != ele[1][16];
    ele[1][6] != ele[1][17];
    ele[1][6] != ele[1][18];
    ele[1][6] != ele[1][19];
    ele[1][6] != ele[1][20];
    ele[1][6] != ele[1][21];
    ele[1][6] != ele[1][22];
    ele[1][6] != ele[1][23];
    ele[1][6] != ele[1][24];
    ele[1][6] != ele[1][25];
    ele[1][6] != ele[1][26];
    ele[1][6] != ele[1][27];
    ele[1][6] != ele[1][28];
    ele[1][6] != ele[1][29];
    ele[1][6] != ele[1][30];
    ele[1][6] != ele[1][31];
    ele[1][6] != ele[1][32];
    ele[1][6] != ele[1][33];
    ele[1][6] != ele[1][34];
    ele[1][6] != ele[1][35];
    ele[1][6] != ele[1][7];
    ele[1][6] != ele[1][8];
    ele[1][6] != ele[1][9];
    ele[1][6] != ele[10][6];
    ele[1][6] != ele[11][6];
    ele[1][6] != ele[12][6];
    ele[1][6] != ele[13][6];
    ele[1][6] != ele[14][6];
    ele[1][6] != ele[15][6];
    ele[1][6] != ele[16][6];
    ele[1][6] != ele[17][6];
    ele[1][6] != ele[18][6];
    ele[1][6] != ele[19][6];
    ele[1][6] != ele[2][10];
    ele[1][6] != ele[2][11];
    ele[1][6] != ele[2][6];
    ele[1][6] != ele[2][7];
    ele[1][6] != ele[2][8];
    ele[1][6] != ele[2][9];
    ele[1][6] != ele[20][6];
    ele[1][6] != ele[21][6];
    ele[1][6] != ele[22][6];
    ele[1][6] != ele[23][6];
    ele[1][6] != ele[24][6];
    ele[1][6] != ele[25][6];
    ele[1][6] != ele[26][6];
    ele[1][6] != ele[27][6];
    ele[1][6] != ele[28][6];
    ele[1][6] != ele[29][6];
    ele[1][6] != ele[3][10];
    ele[1][6] != ele[3][11];
    ele[1][6] != ele[3][6];
    ele[1][6] != ele[3][7];
    ele[1][6] != ele[3][8];
    ele[1][6] != ele[3][9];
    ele[1][6] != ele[30][6];
    ele[1][6] != ele[31][6];
    ele[1][6] != ele[32][6];
    ele[1][6] != ele[33][6];
    ele[1][6] != ele[34][6];
    ele[1][6] != ele[35][6];
    ele[1][6] != ele[4][10];
    ele[1][6] != ele[4][11];
    ele[1][6] != ele[4][6];
    ele[1][6] != ele[4][7];
    ele[1][6] != ele[4][8];
    ele[1][6] != ele[4][9];
    ele[1][6] != ele[5][10];
    ele[1][6] != ele[5][11];
    ele[1][6] != ele[5][6];
    ele[1][6] != ele[5][7];
    ele[1][6] != ele[5][8];
    ele[1][6] != ele[5][9];
    ele[1][6] != ele[6][6];
    ele[1][6] != ele[7][6];
    ele[1][6] != ele[8][6];
    ele[1][6] != ele[9][6];
    ele[1][7] != ele[1][10];
    ele[1][7] != ele[1][11];
    ele[1][7] != ele[1][12];
    ele[1][7] != ele[1][13];
    ele[1][7] != ele[1][14];
    ele[1][7] != ele[1][15];
    ele[1][7] != ele[1][16];
    ele[1][7] != ele[1][17];
    ele[1][7] != ele[1][18];
    ele[1][7] != ele[1][19];
    ele[1][7] != ele[1][20];
    ele[1][7] != ele[1][21];
    ele[1][7] != ele[1][22];
    ele[1][7] != ele[1][23];
    ele[1][7] != ele[1][24];
    ele[1][7] != ele[1][25];
    ele[1][7] != ele[1][26];
    ele[1][7] != ele[1][27];
    ele[1][7] != ele[1][28];
    ele[1][7] != ele[1][29];
    ele[1][7] != ele[1][30];
    ele[1][7] != ele[1][31];
    ele[1][7] != ele[1][32];
    ele[1][7] != ele[1][33];
    ele[1][7] != ele[1][34];
    ele[1][7] != ele[1][35];
    ele[1][7] != ele[1][8];
    ele[1][7] != ele[1][9];
    ele[1][7] != ele[10][7];
    ele[1][7] != ele[11][7];
    ele[1][7] != ele[12][7];
    ele[1][7] != ele[13][7];
    ele[1][7] != ele[14][7];
    ele[1][7] != ele[15][7];
    ele[1][7] != ele[16][7];
    ele[1][7] != ele[17][7];
    ele[1][7] != ele[18][7];
    ele[1][7] != ele[19][7];
    ele[1][7] != ele[2][10];
    ele[1][7] != ele[2][11];
    ele[1][7] != ele[2][6];
    ele[1][7] != ele[2][7];
    ele[1][7] != ele[2][8];
    ele[1][7] != ele[2][9];
    ele[1][7] != ele[20][7];
    ele[1][7] != ele[21][7];
    ele[1][7] != ele[22][7];
    ele[1][7] != ele[23][7];
    ele[1][7] != ele[24][7];
    ele[1][7] != ele[25][7];
    ele[1][7] != ele[26][7];
    ele[1][7] != ele[27][7];
    ele[1][7] != ele[28][7];
    ele[1][7] != ele[29][7];
    ele[1][7] != ele[3][10];
    ele[1][7] != ele[3][11];
    ele[1][7] != ele[3][6];
    ele[1][7] != ele[3][7];
    ele[1][7] != ele[3][8];
    ele[1][7] != ele[3][9];
    ele[1][7] != ele[30][7];
    ele[1][7] != ele[31][7];
    ele[1][7] != ele[32][7];
    ele[1][7] != ele[33][7];
    ele[1][7] != ele[34][7];
    ele[1][7] != ele[35][7];
    ele[1][7] != ele[4][10];
    ele[1][7] != ele[4][11];
    ele[1][7] != ele[4][6];
    ele[1][7] != ele[4][7];
    ele[1][7] != ele[4][8];
    ele[1][7] != ele[4][9];
    ele[1][7] != ele[5][10];
    ele[1][7] != ele[5][11];
    ele[1][7] != ele[5][6];
    ele[1][7] != ele[5][7];
    ele[1][7] != ele[5][8];
    ele[1][7] != ele[5][9];
    ele[1][7] != ele[6][7];
    ele[1][7] != ele[7][7];
    ele[1][7] != ele[8][7];
    ele[1][7] != ele[9][7];
    ele[1][8] != ele[1][10];
    ele[1][8] != ele[1][11];
    ele[1][8] != ele[1][12];
    ele[1][8] != ele[1][13];
    ele[1][8] != ele[1][14];
    ele[1][8] != ele[1][15];
    ele[1][8] != ele[1][16];
    ele[1][8] != ele[1][17];
    ele[1][8] != ele[1][18];
    ele[1][8] != ele[1][19];
    ele[1][8] != ele[1][20];
    ele[1][8] != ele[1][21];
    ele[1][8] != ele[1][22];
    ele[1][8] != ele[1][23];
    ele[1][8] != ele[1][24];
    ele[1][8] != ele[1][25];
    ele[1][8] != ele[1][26];
    ele[1][8] != ele[1][27];
    ele[1][8] != ele[1][28];
    ele[1][8] != ele[1][29];
    ele[1][8] != ele[1][30];
    ele[1][8] != ele[1][31];
    ele[1][8] != ele[1][32];
    ele[1][8] != ele[1][33];
    ele[1][8] != ele[1][34];
    ele[1][8] != ele[1][35];
    ele[1][8] != ele[1][9];
    ele[1][8] != ele[10][8];
    ele[1][8] != ele[11][8];
    ele[1][8] != ele[12][8];
    ele[1][8] != ele[13][8];
    ele[1][8] != ele[14][8];
    ele[1][8] != ele[15][8];
    ele[1][8] != ele[16][8];
    ele[1][8] != ele[17][8];
    ele[1][8] != ele[18][8];
    ele[1][8] != ele[19][8];
    ele[1][8] != ele[2][10];
    ele[1][8] != ele[2][11];
    ele[1][8] != ele[2][6];
    ele[1][8] != ele[2][7];
    ele[1][8] != ele[2][8];
    ele[1][8] != ele[2][9];
    ele[1][8] != ele[20][8];
    ele[1][8] != ele[21][8];
    ele[1][8] != ele[22][8];
    ele[1][8] != ele[23][8];
    ele[1][8] != ele[24][8];
    ele[1][8] != ele[25][8];
    ele[1][8] != ele[26][8];
    ele[1][8] != ele[27][8];
    ele[1][8] != ele[28][8];
    ele[1][8] != ele[29][8];
    ele[1][8] != ele[3][10];
    ele[1][8] != ele[3][11];
    ele[1][8] != ele[3][6];
    ele[1][8] != ele[3][7];
    ele[1][8] != ele[3][8];
    ele[1][8] != ele[3][9];
    ele[1][8] != ele[30][8];
    ele[1][8] != ele[31][8];
    ele[1][8] != ele[32][8];
    ele[1][8] != ele[33][8];
    ele[1][8] != ele[34][8];
    ele[1][8] != ele[35][8];
    ele[1][8] != ele[4][10];
    ele[1][8] != ele[4][11];
    ele[1][8] != ele[4][6];
    ele[1][8] != ele[4][7];
    ele[1][8] != ele[4][8];
    ele[1][8] != ele[4][9];
    ele[1][8] != ele[5][10];
    ele[1][8] != ele[5][11];
    ele[1][8] != ele[5][6];
    ele[1][8] != ele[5][7];
    ele[1][8] != ele[5][8];
    ele[1][8] != ele[5][9];
    ele[1][8] != ele[6][8];
    ele[1][8] != ele[7][8];
    ele[1][8] != ele[8][8];
    ele[1][8] != ele[9][8];
    ele[1][9] != ele[1][10];
    ele[1][9] != ele[1][11];
    ele[1][9] != ele[1][12];
    ele[1][9] != ele[1][13];
    ele[1][9] != ele[1][14];
    ele[1][9] != ele[1][15];
    ele[1][9] != ele[1][16];
    ele[1][9] != ele[1][17];
    ele[1][9] != ele[1][18];
    ele[1][9] != ele[1][19];
    ele[1][9] != ele[1][20];
    ele[1][9] != ele[1][21];
    ele[1][9] != ele[1][22];
    ele[1][9] != ele[1][23];
    ele[1][9] != ele[1][24];
    ele[1][9] != ele[1][25];
    ele[1][9] != ele[1][26];
    ele[1][9] != ele[1][27];
    ele[1][9] != ele[1][28];
    ele[1][9] != ele[1][29];
    ele[1][9] != ele[1][30];
    ele[1][9] != ele[1][31];
    ele[1][9] != ele[1][32];
    ele[1][9] != ele[1][33];
    ele[1][9] != ele[1][34];
    ele[1][9] != ele[1][35];
    ele[1][9] != ele[10][9];
    ele[1][9] != ele[11][9];
    ele[1][9] != ele[12][9];
    ele[1][9] != ele[13][9];
    ele[1][9] != ele[14][9];
    ele[1][9] != ele[15][9];
    ele[1][9] != ele[16][9];
    ele[1][9] != ele[17][9];
    ele[1][9] != ele[18][9];
    ele[1][9] != ele[19][9];
    ele[1][9] != ele[2][10];
    ele[1][9] != ele[2][11];
    ele[1][9] != ele[2][6];
    ele[1][9] != ele[2][7];
    ele[1][9] != ele[2][8];
    ele[1][9] != ele[2][9];
    ele[1][9] != ele[20][9];
    ele[1][9] != ele[21][9];
    ele[1][9] != ele[22][9];
    ele[1][9] != ele[23][9];
    ele[1][9] != ele[24][9];
    ele[1][9] != ele[25][9];
    ele[1][9] != ele[26][9];
    ele[1][9] != ele[27][9];
    ele[1][9] != ele[28][9];
    ele[1][9] != ele[29][9];
    ele[1][9] != ele[3][10];
    ele[1][9] != ele[3][11];
    ele[1][9] != ele[3][6];
    ele[1][9] != ele[3][7];
    ele[1][9] != ele[3][8];
    ele[1][9] != ele[3][9];
    ele[1][9] != ele[30][9];
    ele[1][9] != ele[31][9];
    ele[1][9] != ele[32][9];
    ele[1][9] != ele[33][9];
    ele[1][9] != ele[34][9];
    ele[1][9] != ele[35][9];
    ele[1][9] != ele[4][10];
    ele[1][9] != ele[4][11];
    ele[1][9] != ele[4][6];
    ele[1][9] != ele[4][7];
    ele[1][9] != ele[4][8];
    ele[1][9] != ele[4][9];
    ele[1][9] != ele[5][10];
    ele[1][9] != ele[5][11];
    ele[1][9] != ele[5][6];
    ele[1][9] != ele[5][7];
    ele[1][9] != ele[5][8];
    ele[1][9] != ele[5][9];
    ele[1][9] != ele[6][9];
    ele[1][9] != ele[7][9];
    ele[1][9] != ele[8][9];
    ele[1][9] != ele[9][9];
    ele[10][0] != ele[10][1];
    ele[10][0] != ele[10][10];
    ele[10][0] != ele[10][11];
    ele[10][0] != ele[10][12];
    ele[10][0] != ele[10][13];
    ele[10][0] != ele[10][14];
    ele[10][0] != ele[10][15];
    ele[10][0] != ele[10][16];
    ele[10][0] != ele[10][17];
    ele[10][0] != ele[10][18];
    ele[10][0] != ele[10][19];
    ele[10][0] != ele[10][2];
    ele[10][0] != ele[10][20];
    ele[10][0] != ele[10][21];
    ele[10][0] != ele[10][22];
    ele[10][0] != ele[10][23];
    ele[10][0] != ele[10][24];
    ele[10][0] != ele[10][25];
    ele[10][0] != ele[10][26];
    ele[10][0] != ele[10][27];
    ele[10][0] != ele[10][28];
    ele[10][0] != ele[10][29];
    ele[10][0] != ele[10][3];
    ele[10][0] != ele[10][30];
    ele[10][0] != ele[10][31];
    ele[10][0] != ele[10][32];
    ele[10][0] != ele[10][33];
    ele[10][0] != ele[10][34];
    ele[10][0] != ele[10][35];
    ele[10][0] != ele[10][4];
    ele[10][0] != ele[10][5];
    ele[10][0] != ele[10][6];
    ele[10][0] != ele[10][7];
    ele[10][0] != ele[10][8];
    ele[10][0] != ele[10][9];
    ele[10][0] != ele[11][0];
    ele[10][0] != ele[11][1];
    ele[10][0] != ele[11][2];
    ele[10][0] != ele[11][3];
    ele[10][0] != ele[11][4];
    ele[10][0] != ele[11][5];
    ele[10][0] != ele[12][0];
    ele[10][0] != ele[13][0];
    ele[10][0] != ele[14][0];
    ele[10][0] != ele[15][0];
    ele[10][0] != ele[16][0];
    ele[10][0] != ele[17][0];
    ele[10][0] != ele[18][0];
    ele[10][0] != ele[19][0];
    ele[10][0] != ele[20][0];
    ele[10][0] != ele[21][0];
    ele[10][0] != ele[22][0];
    ele[10][0] != ele[23][0];
    ele[10][0] != ele[24][0];
    ele[10][0] != ele[25][0];
    ele[10][0] != ele[26][0];
    ele[10][0] != ele[27][0];
    ele[10][0] != ele[28][0];
    ele[10][0] != ele[29][0];
    ele[10][0] != ele[30][0];
    ele[10][0] != ele[31][0];
    ele[10][0] != ele[32][0];
    ele[10][0] != ele[33][0];
    ele[10][0] != ele[34][0];
    ele[10][0] != ele[35][0];
    ele[10][1] != ele[10][10];
    ele[10][1] != ele[10][11];
    ele[10][1] != ele[10][12];
    ele[10][1] != ele[10][13];
    ele[10][1] != ele[10][14];
    ele[10][1] != ele[10][15];
    ele[10][1] != ele[10][16];
    ele[10][1] != ele[10][17];
    ele[10][1] != ele[10][18];
    ele[10][1] != ele[10][19];
    ele[10][1] != ele[10][2];
    ele[10][1] != ele[10][20];
    ele[10][1] != ele[10][21];
    ele[10][1] != ele[10][22];
    ele[10][1] != ele[10][23];
    ele[10][1] != ele[10][24];
    ele[10][1] != ele[10][25];
    ele[10][1] != ele[10][26];
    ele[10][1] != ele[10][27];
    ele[10][1] != ele[10][28];
    ele[10][1] != ele[10][29];
    ele[10][1] != ele[10][3];
    ele[10][1] != ele[10][30];
    ele[10][1] != ele[10][31];
    ele[10][1] != ele[10][32];
    ele[10][1] != ele[10][33];
    ele[10][1] != ele[10][34];
    ele[10][1] != ele[10][35];
    ele[10][1] != ele[10][4];
    ele[10][1] != ele[10][5];
    ele[10][1] != ele[10][6];
    ele[10][1] != ele[10][7];
    ele[10][1] != ele[10][8];
    ele[10][1] != ele[10][9];
    ele[10][1] != ele[11][0];
    ele[10][1] != ele[11][1];
    ele[10][1] != ele[11][2];
    ele[10][1] != ele[11][3];
    ele[10][1] != ele[11][4];
    ele[10][1] != ele[11][5];
    ele[10][1] != ele[12][1];
    ele[10][1] != ele[13][1];
    ele[10][1] != ele[14][1];
    ele[10][1] != ele[15][1];
    ele[10][1] != ele[16][1];
    ele[10][1] != ele[17][1];
    ele[10][1] != ele[18][1];
    ele[10][1] != ele[19][1];
    ele[10][1] != ele[20][1];
    ele[10][1] != ele[21][1];
    ele[10][1] != ele[22][1];
    ele[10][1] != ele[23][1];
    ele[10][1] != ele[24][1];
    ele[10][1] != ele[25][1];
    ele[10][1] != ele[26][1];
    ele[10][1] != ele[27][1];
    ele[10][1] != ele[28][1];
    ele[10][1] != ele[29][1];
    ele[10][1] != ele[30][1];
    ele[10][1] != ele[31][1];
    ele[10][1] != ele[32][1];
    ele[10][1] != ele[33][1];
    ele[10][1] != ele[34][1];
    ele[10][1] != ele[35][1];
    ele[10][10] != ele[10][11];
    ele[10][10] != ele[10][12];
    ele[10][10] != ele[10][13];
    ele[10][10] != ele[10][14];
    ele[10][10] != ele[10][15];
    ele[10][10] != ele[10][16];
    ele[10][10] != ele[10][17];
    ele[10][10] != ele[10][18];
    ele[10][10] != ele[10][19];
    ele[10][10] != ele[10][20];
    ele[10][10] != ele[10][21];
    ele[10][10] != ele[10][22];
    ele[10][10] != ele[10][23];
    ele[10][10] != ele[10][24];
    ele[10][10] != ele[10][25];
    ele[10][10] != ele[10][26];
    ele[10][10] != ele[10][27];
    ele[10][10] != ele[10][28];
    ele[10][10] != ele[10][29];
    ele[10][10] != ele[10][30];
    ele[10][10] != ele[10][31];
    ele[10][10] != ele[10][32];
    ele[10][10] != ele[10][33];
    ele[10][10] != ele[10][34];
    ele[10][10] != ele[10][35];
    ele[10][10] != ele[11][10];
    ele[10][10] != ele[11][11];
    ele[10][10] != ele[11][6];
    ele[10][10] != ele[11][7];
    ele[10][10] != ele[11][8];
    ele[10][10] != ele[11][9];
    ele[10][10] != ele[12][10];
    ele[10][10] != ele[13][10];
    ele[10][10] != ele[14][10];
    ele[10][10] != ele[15][10];
    ele[10][10] != ele[16][10];
    ele[10][10] != ele[17][10];
    ele[10][10] != ele[18][10];
    ele[10][10] != ele[19][10];
    ele[10][10] != ele[20][10];
    ele[10][10] != ele[21][10];
    ele[10][10] != ele[22][10];
    ele[10][10] != ele[23][10];
    ele[10][10] != ele[24][10];
    ele[10][10] != ele[25][10];
    ele[10][10] != ele[26][10];
    ele[10][10] != ele[27][10];
    ele[10][10] != ele[28][10];
    ele[10][10] != ele[29][10];
    ele[10][10] != ele[30][10];
    ele[10][10] != ele[31][10];
    ele[10][10] != ele[32][10];
    ele[10][10] != ele[33][10];
    ele[10][10] != ele[34][10];
    ele[10][10] != ele[35][10];
    ele[10][11] != ele[10][12];
    ele[10][11] != ele[10][13];
    ele[10][11] != ele[10][14];
    ele[10][11] != ele[10][15];
    ele[10][11] != ele[10][16];
    ele[10][11] != ele[10][17];
    ele[10][11] != ele[10][18];
    ele[10][11] != ele[10][19];
    ele[10][11] != ele[10][20];
    ele[10][11] != ele[10][21];
    ele[10][11] != ele[10][22];
    ele[10][11] != ele[10][23];
    ele[10][11] != ele[10][24];
    ele[10][11] != ele[10][25];
    ele[10][11] != ele[10][26];
    ele[10][11] != ele[10][27];
    ele[10][11] != ele[10][28];
    ele[10][11] != ele[10][29];
    ele[10][11] != ele[10][30];
    ele[10][11] != ele[10][31];
    ele[10][11] != ele[10][32];
    ele[10][11] != ele[10][33];
    ele[10][11] != ele[10][34];
    ele[10][11] != ele[10][35];
    ele[10][11] != ele[11][10];
    ele[10][11] != ele[11][11];
    ele[10][11] != ele[11][6];
    ele[10][11] != ele[11][7];
    ele[10][11] != ele[11][8];
    ele[10][11] != ele[11][9];
    ele[10][11] != ele[12][11];
    ele[10][11] != ele[13][11];
    ele[10][11] != ele[14][11];
    ele[10][11] != ele[15][11];
    ele[10][11] != ele[16][11];
    ele[10][11] != ele[17][11];
    ele[10][11] != ele[18][11];
    ele[10][11] != ele[19][11];
    ele[10][11] != ele[20][11];
    ele[10][11] != ele[21][11];
    ele[10][11] != ele[22][11];
    ele[10][11] != ele[23][11];
    ele[10][11] != ele[24][11];
    ele[10][11] != ele[25][11];
    ele[10][11] != ele[26][11];
    ele[10][11] != ele[27][11];
    ele[10][11] != ele[28][11];
    ele[10][11] != ele[29][11];
    ele[10][11] != ele[30][11];
    ele[10][11] != ele[31][11];
    ele[10][11] != ele[32][11];
    ele[10][11] != ele[33][11];
    ele[10][11] != ele[34][11];
    ele[10][11] != ele[35][11];
    ele[10][12] != ele[10][13];
    ele[10][12] != ele[10][14];
    ele[10][12] != ele[10][15];
    ele[10][12] != ele[10][16];
    ele[10][12] != ele[10][17];
    ele[10][12] != ele[10][18];
    ele[10][12] != ele[10][19];
    ele[10][12] != ele[10][20];
    ele[10][12] != ele[10][21];
    ele[10][12] != ele[10][22];
    ele[10][12] != ele[10][23];
    ele[10][12] != ele[10][24];
    ele[10][12] != ele[10][25];
    ele[10][12] != ele[10][26];
    ele[10][12] != ele[10][27];
    ele[10][12] != ele[10][28];
    ele[10][12] != ele[10][29];
    ele[10][12] != ele[10][30];
    ele[10][12] != ele[10][31];
    ele[10][12] != ele[10][32];
    ele[10][12] != ele[10][33];
    ele[10][12] != ele[10][34];
    ele[10][12] != ele[10][35];
    ele[10][12] != ele[11][12];
    ele[10][12] != ele[11][13];
    ele[10][12] != ele[11][14];
    ele[10][12] != ele[11][15];
    ele[10][12] != ele[11][16];
    ele[10][12] != ele[11][17];
    ele[10][12] != ele[12][12];
    ele[10][12] != ele[13][12];
    ele[10][12] != ele[14][12];
    ele[10][12] != ele[15][12];
    ele[10][12] != ele[16][12];
    ele[10][12] != ele[17][12];
    ele[10][12] != ele[18][12];
    ele[10][12] != ele[19][12];
    ele[10][12] != ele[20][12];
    ele[10][12] != ele[21][12];
    ele[10][12] != ele[22][12];
    ele[10][12] != ele[23][12];
    ele[10][12] != ele[24][12];
    ele[10][12] != ele[25][12];
    ele[10][12] != ele[26][12];
    ele[10][12] != ele[27][12];
    ele[10][12] != ele[28][12];
    ele[10][12] != ele[29][12];
    ele[10][12] != ele[30][12];
    ele[10][12] != ele[31][12];
    ele[10][12] != ele[32][12];
    ele[10][12] != ele[33][12];
    ele[10][12] != ele[34][12];
    ele[10][12] != ele[35][12];
    ele[10][13] != ele[10][14];
    ele[10][13] != ele[10][15];
    ele[10][13] != ele[10][16];
    ele[10][13] != ele[10][17];
    ele[10][13] != ele[10][18];
    ele[10][13] != ele[10][19];
    ele[10][13] != ele[10][20];
    ele[10][13] != ele[10][21];
    ele[10][13] != ele[10][22];
    ele[10][13] != ele[10][23];
    ele[10][13] != ele[10][24];
    ele[10][13] != ele[10][25];
    ele[10][13] != ele[10][26];
    ele[10][13] != ele[10][27];
    ele[10][13] != ele[10][28];
    ele[10][13] != ele[10][29];
    ele[10][13] != ele[10][30];
    ele[10][13] != ele[10][31];
    ele[10][13] != ele[10][32];
    ele[10][13] != ele[10][33];
    ele[10][13] != ele[10][34];
    ele[10][13] != ele[10][35];
    ele[10][13] != ele[11][12];
    ele[10][13] != ele[11][13];
    ele[10][13] != ele[11][14];
    ele[10][13] != ele[11][15];
    ele[10][13] != ele[11][16];
    ele[10][13] != ele[11][17];
    ele[10][13] != ele[12][13];
    ele[10][13] != ele[13][13];
    ele[10][13] != ele[14][13];
    ele[10][13] != ele[15][13];
    ele[10][13] != ele[16][13];
    ele[10][13] != ele[17][13];
    ele[10][13] != ele[18][13];
    ele[10][13] != ele[19][13];
    ele[10][13] != ele[20][13];
    ele[10][13] != ele[21][13];
    ele[10][13] != ele[22][13];
    ele[10][13] != ele[23][13];
    ele[10][13] != ele[24][13];
    ele[10][13] != ele[25][13];
    ele[10][13] != ele[26][13];
    ele[10][13] != ele[27][13];
    ele[10][13] != ele[28][13];
    ele[10][13] != ele[29][13];
    ele[10][13] != ele[30][13];
    ele[10][13] != ele[31][13];
    ele[10][13] != ele[32][13];
    ele[10][13] != ele[33][13];
    ele[10][13] != ele[34][13];
    ele[10][13] != ele[35][13];
    ele[10][14] != ele[10][15];
    ele[10][14] != ele[10][16];
    ele[10][14] != ele[10][17];
    ele[10][14] != ele[10][18];
    ele[10][14] != ele[10][19];
    ele[10][14] != ele[10][20];
    ele[10][14] != ele[10][21];
    ele[10][14] != ele[10][22];
    ele[10][14] != ele[10][23];
    ele[10][14] != ele[10][24];
    ele[10][14] != ele[10][25];
    ele[10][14] != ele[10][26];
    ele[10][14] != ele[10][27];
    ele[10][14] != ele[10][28];
    ele[10][14] != ele[10][29];
    ele[10][14] != ele[10][30];
    ele[10][14] != ele[10][31];
    ele[10][14] != ele[10][32];
    ele[10][14] != ele[10][33];
    ele[10][14] != ele[10][34];
    ele[10][14] != ele[10][35];
    ele[10][14] != ele[11][12];
    ele[10][14] != ele[11][13];
    ele[10][14] != ele[11][14];
    ele[10][14] != ele[11][15];
    ele[10][14] != ele[11][16];
    ele[10][14] != ele[11][17];
    ele[10][14] != ele[12][14];
    ele[10][14] != ele[13][14];
    ele[10][14] != ele[14][14];
    ele[10][14] != ele[15][14];
    ele[10][14] != ele[16][14];
    ele[10][14] != ele[17][14];
    ele[10][14] != ele[18][14];
    ele[10][14] != ele[19][14];
    ele[10][14] != ele[20][14];
    ele[10][14] != ele[21][14];
    ele[10][14] != ele[22][14];
    ele[10][14] != ele[23][14];
    ele[10][14] != ele[24][14];
    ele[10][14] != ele[25][14];
    ele[10][14] != ele[26][14];
    ele[10][14] != ele[27][14];
    ele[10][14] != ele[28][14];
    ele[10][14] != ele[29][14];
    ele[10][14] != ele[30][14];
    ele[10][14] != ele[31][14];
    ele[10][14] != ele[32][14];
    ele[10][14] != ele[33][14];
    ele[10][14] != ele[34][14];
    ele[10][14] != ele[35][14];
    ele[10][15] != ele[10][16];
    ele[10][15] != ele[10][17];
    ele[10][15] != ele[10][18];
    ele[10][15] != ele[10][19];
    ele[10][15] != ele[10][20];
    ele[10][15] != ele[10][21];
    ele[10][15] != ele[10][22];
    ele[10][15] != ele[10][23];
    ele[10][15] != ele[10][24];
    ele[10][15] != ele[10][25];
    ele[10][15] != ele[10][26];
    ele[10][15] != ele[10][27];
    ele[10][15] != ele[10][28];
    ele[10][15] != ele[10][29];
    ele[10][15] != ele[10][30];
    ele[10][15] != ele[10][31];
    ele[10][15] != ele[10][32];
    ele[10][15] != ele[10][33];
    ele[10][15] != ele[10][34];
    ele[10][15] != ele[10][35];
    ele[10][15] != ele[11][12];
    ele[10][15] != ele[11][13];
    ele[10][15] != ele[11][14];
    ele[10][15] != ele[11][15];
    ele[10][15] != ele[11][16];
    ele[10][15] != ele[11][17];
    ele[10][15] != ele[12][15];
    ele[10][15] != ele[13][15];
    ele[10][15] != ele[14][15];
    ele[10][15] != ele[15][15];
    ele[10][15] != ele[16][15];
    ele[10][15] != ele[17][15];
    ele[10][15] != ele[18][15];
    ele[10][15] != ele[19][15];
    ele[10][15] != ele[20][15];
    ele[10][15] != ele[21][15];
    ele[10][15] != ele[22][15];
    ele[10][15] != ele[23][15];
    ele[10][15] != ele[24][15];
    ele[10][15] != ele[25][15];
    ele[10][15] != ele[26][15];
    ele[10][15] != ele[27][15];
    ele[10][15] != ele[28][15];
    ele[10][15] != ele[29][15];
    ele[10][15] != ele[30][15];
    ele[10][15] != ele[31][15];
    ele[10][15] != ele[32][15];
    ele[10][15] != ele[33][15];
    ele[10][15] != ele[34][15];
    ele[10][15] != ele[35][15];
    ele[10][16] != ele[10][17];
    ele[10][16] != ele[10][18];
    ele[10][16] != ele[10][19];
    ele[10][16] != ele[10][20];
    ele[10][16] != ele[10][21];
    ele[10][16] != ele[10][22];
    ele[10][16] != ele[10][23];
    ele[10][16] != ele[10][24];
    ele[10][16] != ele[10][25];
    ele[10][16] != ele[10][26];
    ele[10][16] != ele[10][27];
    ele[10][16] != ele[10][28];
    ele[10][16] != ele[10][29];
    ele[10][16] != ele[10][30];
    ele[10][16] != ele[10][31];
    ele[10][16] != ele[10][32];
    ele[10][16] != ele[10][33];
    ele[10][16] != ele[10][34];
    ele[10][16] != ele[10][35];
    ele[10][16] != ele[11][12];
    ele[10][16] != ele[11][13];
    ele[10][16] != ele[11][14];
    ele[10][16] != ele[11][15];
    ele[10][16] != ele[11][16];
    ele[10][16] != ele[11][17];
    ele[10][16] != ele[12][16];
    ele[10][16] != ele[13][16];
    ele[10][16] != ele[14][16];
    ele[10][16] != ele[15][16];
    ele[10][16] != ele[16][16];
    ele[10][16] != ele[17][16];
    ele[10][16] != ele[18][16];
    ele[10][16] != ele[19][16];
    ele[10][16] != ele[20][16];
    ele[10][16] != ele[21][16];
    ele[10][16] != ele[22][16];
    ele[10][16] != ele[23][16];
    ele[10][16] != ele[24][16];
    ele[10][16] != ele[25][16];
    ele[10][16] != ele[26][16];
    ele[10][16] != ele[27][16];
    ele[10][16] != ele[28][16];
    ele[10][16] != ele[29][16];
    ele[10][16] != ele[30][16];
    ele[10][16] != ele[31][16];
    ele[10][16] != ele[32][16];
    ele[10][16] != ele[33][16];
    ele[10][16] != ele[34][16];
    ele[10][16] != ele[35][16];
    ele[10][17] != ele[10][18];
    ele[10][17] != ele[10][19];
    ele[10][17] != ele[10][20];
    ele[10][17] != ele[10][21];
    ele[10][17] != ele[10][22];
    ele[10][17] != ele[10][23];
    ele[10][17] != ele[10][24];
    ele[10][17] != ele[10][25];
    ele[10][17] != ele[10][26];
    ele[10][17] != ele[10][27];
    ele[10][17] != ele[10][28];
    ele[10][17] != ele[10][29];
    ele[10][17] != ele[10][30];
    ele[10][17] != ele[10][31];
    ele[10][17] != ele[10][32];
    ele[10][17] != ele[10][33];
    ele[10][17] != ele[10][34];
    ele[10][17] != ele[10][35];
    ele[10][17] != ele[11][12];
    ele[10][17] != ele[11][13];
    ele[10][17] != ele[11][14];
    ele[10][17] != ele[11][15];
    ele[10][17] != ele[11][16];
    ele[10][17] != ele[11][17];
    ele[10][17] != ele[12][17];
    ele[10][17] != ele[13][17];
    ele[10][17] != ele[14][17];
    ele[10][17] != ele[15][17];
    ele[10][17] != ele[16][17];
    ele[10][17] != ele[17][17];
    ele[10][17] != ele[18][17];
    ele[10][17] != ele[19][17];
    ele[10][17] != ele[20][17];
    ele[10][17] != ele[21][17];
    ele[10][17] != ele[22][17];
    ele[10][17] != ele[23][17];
    ele[10][17] != ele[24][17];
    ele[10][17] != ele[25][17];
    ele[10][17] != ele[26][17];
    ele[10][17] != ele[27][17];
    ele[10][17] != ele[28][17];
    ele[10][17] != ele[29][17];
    ele[10][17] != ele[30][17];
    ele[10][17] != ele[31][17];
    ele[10][17] != ele[32][17];
    ele[10][17] != ele[33][17];
    ele[10][17] != ele[34][17];
    ele[10][17] != ele[35][17];
    ele[10][18] != ele[10][19];
    ele[10][18] != ele[10][20];
    ele[10][18] != ele[10][21];
    ele[10][18] != ele[10][22];
    ele[10][18] != ele[10][23];
    ele[10][18] != ele[10][24];
    ele[10][18] != ele[10][25];
    ele[10][18] != ele[10][26];
    ele[10][18] != ele[10][27];
    ele[10][18] != ele[10][28];
    ele[10][18] != ele[10][29];
    ele[10][18] != ele[10][30];
    ele[10][18] != ele[10][31];
    ele[10][18] != ele[10][32];
    ele[10][18] != ele[10][33];
    ele[10][18] != ele[10][34];
    ele[10][18] != ele[10][35];
    ele[10][18] != ele[11][18];
    ele[10][18] != ele[11][19];
    ele[10][18] != ele[11][20];
    ele[10][18] != ele[11][21];
    ele[10][18] != ele[11][22];
    ele[10][18] != ele[11][23];
    ele[10][18] != ele[12][18];
    ele[10][18] != ele[13][18];
    ele[10][18] != ele[14][18];
    ele[10][18] != ele[15][18];
    ele[10][18] != ele[16][18];
    ele[10][18] != ele[17][18];
    ele[10][18] != ele[18][18];
    ele[10][18] != ele[19][18];
    ele[10][18] != ele[20][18];
    ele[10][18] != ele[21][18];
    ele[10][18] != ele[22][18];
    ele[10][18] != ele[23][18];
    ele[10][18] != ele[24][18];
    ele[10][18] != ele[25][18];
    ele[10][18] != ele[26][18];
    ele[10][18] != ele[27][18];
    ele[10][18] != ele[28][18];
    ele[10][18] != ele[29][18];
    ele[10][18] != ele[30][18];
    ele[10][18] != ele[31][18];
    ele[10][18] != ele[32][18];
    ele[10][18] != ele[33][18];
    ele[10][18] != ele[34][18];
    ele[10][18] != ele[35][18];
    ele[10][19] != ele[10][20];
    ele[10][19] != ele[10][21];
    ele[10][19] != ele[10][22];
    ele[10][19] != ele[10][23];
    ele[10][19] != ele[10][24];
    ele[10][19] != ele[10][25];
    ele[10][19] != ele[10][26];
    ele[10][19] != ele[10][27];
    ele[10][19] != ele[10][28];
    ele[10][19] != ele[10][29];
    ele[10][19] != ele[10][30];
    ele[10][19] != ele[10][31];
    ele[10][19] != ele[10][32];
    ele[10][19] != ele[10][33];
    ele[10][19] != ele[10][34];
    ele[10][19] != ele[10][35];
    ele[10][19] != ele[11][18];
    ele[10][19] != ele[11][19];
    ele[10][19] != ele[11][20];
    ele[10][19] != ele[11][21];
    ele[10][19] != ele[11][22];
    ele[10][19] != ele[11][23];
    ele[10][19] != ele[12][19];
    ele[10][19] != ele[13][19];
    ele[10][19] != ele[14][19];
    ele[10][19] != ele[15][19];
    ele[10][19] != ele[16][19];
    ele[10][19] != ele[17][19];
    ele[10][19] != ele[18][19];
    ele[10][19] != ele[19][19];
    ele[10][19] != ele[20][19];
    ele[10][19] != ele[21][19];
    ele[10][19] != ele[22][19];
    ele[10][19] != ele[23][19];
    ele[10][19] != ele[24][19];
    ele[10][19] != ele[25][19];
    ele[10][19] != ele[26][19];
    ele[10][19] != ele[27][19];
    ele[10][19] != ele[28][19];
    ele[10][19] != ele[29][19];
    ele[10][19] != ele[30][19];
    ele[10][19] != ele[31][19];
    ele[10][19] != ele[32][19];
    ele[10][19] != ele[33][19];
    ele[10][19] != ele[34][19];
    ele[10][19] != ele[35][19];
    ele[10][2] != ele[10][10];
    ele[10][2] != ele[10][11];
    ele[10][2] != ele[10][12];
    ele[10][2] != ele[10][13];
    ele[10][2] != ele[10][14];
    ele[10][2] != ele[10][15];
    ele[10][2] != ele[10][16];
    ele[10][2] != ele[10][17];
    ele[10][2] != ele[10][18];
    ele[10][2] != ele[10][19];
    ele[10][2] != ele[10][20];
    ele[10][2] != ele[10][21];
    ele[10][2] != ele[10][22];
    ele[10][2] != ele[10][23];
    ele[10][2] != ele[10][24];
    ele[10][2] != ele[10][25];
    ele[10][2] != ele[10][26];
    ele[10][2] != ele[10][27];
    ele[10][2] != ele[10][28];
    ele[10][2] != ele[10][29];
    ele[10][2] != ele[10][3];
    ele[10][2] != ele[10][30];
    ele[10][2] != ele[10][31];
    ele[10][2] != ele[10][32];
    ele[10][2] != ele[10][33];
    ele[10][2] != ele[10][34];
    ele[10][2] != ele[10][35];
    ele[10][2] != ele[10][4];
    ele[10][2] != ele[10][5];
    ele[10][2] != ele[10][6];
    ele[10][2] != ele[10][7];
    ele[10][2] != ele[10][8];
    ele[10][2] != ele[10][9];
    ele[10][2] != ele[11][0];
    ele[10][2] != ele[11][1];
    ele[10][2] != ele[11][2];
    ele[10][2] != ele[11][3];
    ele[10][2] != ele[11][4];
    ele[10][2] != ele[11][5];
    ele[10][2] != ele[12][2];
    ele[10][2] != ele[13][2];
    ele[10][2] != ele[14][2];
    ele[10][2] != ele[15][2];
    ele[10][2] != ele[16][2];
    ele[10][2] != ele[17][2];
    ele[10][2] != ele[18][2];
    ele[10][2] != ele[19][2];
    ele[10][2] != ele[20][2];
    ele[10][2] != ele[21][2];
    ele[10][2] != ele[22][2];
    ele[10][2] != ele[23][2];
    ele[10][2] != ele[24][2];
    ele[10][2] != ele[25][2];
    ele[10][2] != ele[26][2];
    ele[10][2] != ele[27][2];
    ele[10][2] != ele[28][2];
    ele[10][2] != ele[29][2];
    ele[10][2] != ele[30][2];
    ele[10][2] != ele[31][2];
    ele[10][2] != ele[32][2];
    ele[10][2] != ele[33][2];
    ele[10][2] != ele[34][2];
    ele[10][2] != ele[35][2];
    ele[10][20] != ele[10][21];
    ele[10][20] != ele[10][22];
    ele[10][20] != ele[10][23];
    ele[10][20] != ele[10][24];
    ele[10][20] != ele[10][25];
    ele[10][20] != ele[10][26];
    ele[10][20] != ele[10][27];
    ele[10][20] != ele[10][28];
    ele[10][20] != ele[10][29];
    ele[10][20] != ele[10][30];
    ele[10][20] != ele[10][31];
    ele[10][20] != ele[10][32];
    ele[10][20] != ele[10][33];
    ele[10][20] != ele[10][34];
    ele[10][20] != ele[10][35];
    ele[10][20] != ele[11][18];
    ele[10][20] != ele[11][19];
    ele[10][20] != ele[11][20];
    ele[10][20] != ele[11][21];
    ele[10][20] != ele[11][22];
    ele[10][20] != ele[11][23];
    ele[10][20] != ele[12][20];
    ele[10][20] != ele[13][20];
    ele[10][20] != ele[14][20];
    ele[10][20] != ele[15][20];
    ele[10][20] != ele[16][20];
    ele[10][20] != ele[17][20];
    ele[10][20] != ele[18][20];
    ele[10][20] != ele[19][20];
    ele[10][20] != ele[20][20];
    ele[10][20] != ele[21][20];
    ele[10][20] != ele[22][20];
    ele[10][20] != ele[23][20];
    ele[10][20] != ele[24][20];
    ele[10][20] != ele[25][20];
    ele[10][20] != ele[26][20];
    ele[10][20] != ele[27][20];
    ele[10][20] != ele[28][20];
    ele[10][20] != ele[29][20];
    ele[10][20] != ele[30][20];
    ele[10][20] != ele[31][20];
    ele[10][20] != ele[32][20];
    ele[10][20] != ele[33][20];
    ele[10][20] != ele[34][20];
    ele[10][20] != ele[35][20];
    ele[10][21] != ele[10][22];
    ele[10][21] != ele[10][23];
    ele[10][21] != ele[10][24];
    ele[10][21] != ele[10][25];
    ele[10][21] != ele[10][26];
    ele[10][21] != ele[10][27];
    ele[10][21] != ele[10][28];
    ele[10][21] != ele[10][29];
    ele[10][21] != ele[10][30];
    ele[10][21] != ele[10][31];
    ele[10][21] != ele[10][32];
    ele[10][21] != ele[10][33];
    ele[10][21] != ele[10][34];
    ele[10][21] != ele[10][35];
    ele[10][21] != ele[11][18];
    ele[10][21] != ele[11][19];
    ele[10][21] != ele[11][20];
    ele[10][21] != ele[11][21];
    ele[10][21] != ele[11][22];
    ele[10][21] != ele[11][23];
    ele[10][21] != ele[12][21];
    ele[10][21] != ele[13][21];
    ele[10][21] != ele[14][21];
    ele[10][21] != ele[15][21];
    ele[10][21] != ele[16][21];
    ele[10][21] != ele[17][21];
    ele[10][21] != ele[18][21];
    ele[10][21] != ele[19][21];
    ele[10][21] != ele[20][21];
    ele[10][21] != ele[21][21];
    ele[10][21] != ele[22][21];
    ele[10][21] != ele[23][21];
    ele[10][21] != ele[24][21];
    ele[10][21] != ele[25][21];
    ele[10][21] != ele[26][21];
    ele[10][21] != ele[27][21];
    ele[10][21] != ele[28][21];
    ele[10][21] != ele[29][21];
    ele[10][21] != ele[30][21];
    ele[10][21] != ele[31][21];
    ele[10][21] != ele[32][21];
    ele[10][21] != ele[33][21];
    ele[10][21] != ele[34][21];
    ele[10][21] != ele[35][21];
    ele[10][22] != ele[10][23];
    ele[10][22] != ele[10][24];
    ele[10][22] != ele[10][25];
    ele[10][22] != ele[10][26];
    ele[10][22] != ele[10][27];
    ele[10][22] != ele[10][28];
    ele[10][22] != ele[10][29];
    ele[10][22] != ele[10][30];
    ele[10][22] != ele[10][31];
    ele[10][22] != ele[10][32];
    ele[10][22] != ele[10][33];
    ele[10][22] != ele[10][34];
    ele[10][22] != ele[10][35];
    ele[10][22] != ele[11][18];
    ele[10][22] != ele[11][19];
    ele[10][22] != ele[11][20];
    ele[10][22] != ele[11][21];
    ele[10][22] != ele[11][22];
    ele[10][22] != ele[11][23];
    ele[10][22] != ele[12][22];
    ele[10][22] != ele[13][22];
    ele[10][22] != ele[14][22];
    ele[10][22] != ele[15][22];
    ele[10][22] != ele[16][22];
    ele[10][22] != ele[17][22];
    ele[10][22] != ele[18][22];
    ele[10][22] != ele[19][22];
    ele[10][22] != ele[20][22];
    ele[10][22] != ele[21][22];
    ele[10][22] != ele[22][22];
    ele[10][22] != ele[23][22];
    ele[10][22] != ele[24][22];
    ele[10][22] != ele[25][22];
    ele[10][22] != ele[26][22];
    ele[10][22] != ele[27][22];
    ele[10][22] != ele[28][22];
    ele[10][22] != ele[29][22];
    ele[10][22] != ele[30][22];
    ele[10][22] != ele[31][22];
    ele[10][22] != ele[32][22];
    ele[10][22] != ele[33][22];
    ele[10][22] != ele[34][22];
    ele[10][22] != ele[35][22];
    ele[10][23] != ele[10][24];
    ele[10][23] != ele[10][25];
    ele[10][23] != ele[10][26];
    ele[10][23] != ele[10][27];
    ele[10][23] != ele[10][28];
    ele[10][23] != ele[10][29];
    ele[10][23] != ele[10][30];
    ele[10][23] != ele[10][31];
    ele[10][23] != ele[10][32];
    ele[10][23] != ele[10][33];
    ele[10][23] != ele[10][34];
    ele[10][23] != ele[10][35];
    ele[10][23] != ele[11][18];
    ele[10][23] != ele[11][19];
    ele[10][23] != ele[11][20];
    ele[10][23] != ele[11][21];
    ele[10][23] != ele[11][22];
    ele[10][23] != ele[11][23];
    ele[10][23] != ele[12][23];
    ele[10][23] != ele[13][23];
    ele[10][23] != ele[14][23];
    ele[10][23] != ele[15][23];
    ele[10][23] != ele[16][23];
    ele[10][23] != ele[17][23];
    ele[10][23] != ele[18][23];
    ele[10][23] != ele[19][23];
    ele[10][23] != ele[20][23];
    ele[10][23] != ele[21][23];
    ele[10][23] != ele[22][23];
    ele[10][23] != ele[23][23];
    ele[10][23] != ele[24][23];
    ele[10][23] != ele[25][23];
    ele[10][23] != ele[26][23];
    ele[10][23] != ele[27][23];
    ele[10][23] != ele[28][23];
    ele[10][23] != ele[29][23];
    ele[10][23] != ele[30][23];
    ele[10][23] != ele[31][23];
    ele[10][23] != ele[32][23];
    ele[10][23] != ele[33][23];
    ele[10][23] != ele[34][23];
    ele[10][23] != ele[35][23];
    ele[10][24] != ele[10][25];
    ele[10][24] != ele[10][26];
    ele[10][24] != ele[10][27];
    ele[10][24] != ele[10][28];
    ele[10][24] != ele[10][29];
    ele[10][24] != ele[10][30];
    ele[10][24] != ele[10][31];
    ele[10][24] != ele[10][32];
    ele[10][24] != ele[10][33];
    ele[10][24] != ele[10][34];
    ele[10][24] != ele[10][35];
    ele[10][24] != ele[11][24];
    ele[10][24] != ele[11][25];
    ele[10][24] != ele[11][26];
    ele[10][24] != ele[11][27];
    ele[10][24] != ele[11][28];
    ele[10][24] != ele[11][29];
    ele[10][24] != ele[12][24];
    ele[10][24] != ele[13][24];
    ele[10][24] != ele[14][24];
    ele[10][24] != ele[15][24];
    ele[10][24] != ele[16][24];
    ele[10][24] != ele[17][24];
    ele[10][24] != ele[18][24];
    ele[10][24] != ele[19][24];
    ele[10][24] != ele[20][24];
    ele[10][24] != ele[21][24];
    ele[10][24] != ele[22][24];
    ele[10][24] != ele[23][24];
    ele[10][24] != ele[24][24];
    ele[10][24] != ele[25][24];
    ele[10][24] != ele[26][24];
    ele[10][24] != ele[27][24];
    ele[10][24] != ele[28][24];
    ele[10][24] != ele[29][24];
    ele[10][24] != ele[30][24];
    ele[10][24] != ele[31][24];
    ele[10][24] != ele[32][24];
    ele[10][24] != ele[33][24];
    ele[10][24] != ele[34][24];
    ele[10][24] != ele[35][24];
    ele[10][25] != ele[10][26];
    ele[10][25] != ele[10][27];
    ele[10][25] != ele[10][28];
    ele[10][25] != ele[10][29];
    ele[10][25] != ele[10][30];
    ele[10][25] != ele[10][31];
    ele[10][25] != ele[10][32];
    ele[10][25] != ele[10][33];
    ele[10][25] != ele[10][34];
    ele[10][25] != ele[10][35];
    ele[10][25] != ele[11][24];
    ele[10][25] != ele[11][25];
    ele[10][25] != ele[11][26];
    ele[10][25] != ele[11][27];
    ele[10][25] != ele[11][28];
    ele[10][25] != ele[11][29];
    ele[10][25] != ele[12][25];
    ele[10][25] != ele[13][25];
    ele[10][25] != ele[14][25];
    ele[10][25] != ele[15][25];
    ele[10][25] != ele[16][25];
    ele[10][25] != ele[17][25];
    ele[10][25] != ele[18][25];
    ele[10][25] != ele[19][25];
    ele[10][25] != ele[20][25];
    ele[10][25] != ele[21][25];
    ele[10][25] != ele[22][25];
    ele[10][25] != ele[23][25];
    ele[10][25] != ele[24][25];
    ele[10][25] != ele[25][25];
    ele[10][25] != ele[26][25];
    ele[10][25] != ele[27][25];
    ele[10][25] != ele[28][25];
    ele[10][25] != ele[29][25];
    ele[10][25] != ele[30][25];
    ele[10][25] != ele[31][25];
    ele[10][25] != ele[32][25];
    ele[10][25] != ele[33][25];
    ele[10][25] != ele[34][25];
    ele[10][25] != ele[35][25];
    ele[10][26] != ele[10][27];
    ele[10][26] != ele[10][28];
    ele[10][26] != ele[10][29];
    ele[10][26] != ele[10][30];
    ele[10][26] != ele[10][31];
    ele[10][26] != ele[10][32];
    ele[10][26] != ele[10][33];
    ele[10][26] != ele[10][34];
    ele[10][26] != ele[10][35];
    ele[10][26] != ele[11][24];
    ele[10][26] != ele[11][25];
    ele[10][26] != ele[11][26];
    ele[10][26] != ele[11][27];
    ele[10][26] != ele[11][28];
    ele[10][26] != ele[11][29];
    ele[10][26] != ele[12][26];
    ele[10][26] != ele[13][26];
    ele[10][26] != ele[14][26];
    ele[10][26] != ele[15][26];
    ele[10][26] != ele[16][26];
    ele[10][26] != ele[17][26];
    ele[10][26] != ele[18][26];
    ele[10][26] != ele[19][26];
    ele[10][26] != ele[20][26];
    ele[10][26] != ele[21][26];
    ele[10][26] != ele[22][26];
    ele[10][26] != ele[23][26];
    ele[10][26] != ele[24][26];
    ele[10][26] != ele[25][26];
    ele[10][26] != ele[26][26];
    ele[10][26] != ele[27][26];
    ele[10][26] != ele[28][26];
    ele[10][26] != ele[29][26];
    ele[10][26] != ele[30][26];
    ele[10][26] != ele[31][26];
    ele[10][26] != ele[32][26];
    ele[10][26] != ele[33][26];
    ele[10][26] != ele[34][26];
    ele[10][26] != ele[35][26];
    ele[10][27] != ele[10][28];
    ele[10][27] != ele[10][29];
    ele[10][27] != ele[10][30];
    ele[10][27] != ele[10][31];
    ele[10][27] != ele[10][32];
    ele[10][27] != ele[10][33];
    ele[10][27] != ele[10][34];
    ele[10][27] != ele[10][35];
    ele[10][27] != ele[11][24];
    ele[10][27] != ele[11][25];
    ele[10][27] != ele[11][26];
    ele[10][27] != ele[11][27];
    ele[10][27] != ele[11][28];
    ele[10][27] != ele[11][29];
    ele[10][27] != ele[12][27];
    ele[10][27] != ele[13][27];
    ele[10][27] != ele[14][27];
    ele[10][27] != ele[15][27];
    ele[10][27] != ele[16][27];
    ele[10][27] != ele[17][27];
    ele[10][27] != ele[18][27];
    ele[10][27] != ele[19][27];
    ele[10][27] != ele[20][27];
    ele[10][27] != ele[21][27];
    ele[10][27] != ele[22][27];
    ele[10][27] != ele[23][27];
    ele[10][27] != ele[24][27];
    ele[10][27] != ele[25][27];
    ele[10][27] != ele[26][27];
    ele[10][27] != ele[27][27];
    ele[10][27] != ele[28][27];
    ele[10][27] != ele[29][27];
    ele[10][27] != ele[30][27];
    ele[10][27] != ele[31][27];
    ele[10][27] != ele[32][27];
    ele[10][27] != ele[33][27];
    ele[10][27] != ele[34][27];
    ele[10][27] != ele[35][27];
    ele[10][28] != ele[10][29];
    ele[10][28] != ele[10][30];
    ele[10][28] != ele[10][31];
    ele[10][28] != ele[10][32];
    ele[10][28] != ele[10][33];
    ele[10][28] != ele[10][34];
    ele[10][28] != ele[10][35];
    ele[10][28] != ele[11][24];
    ele[10][28] != ele[11][25];
    ele[10][28] != ele[11][26];
    ele[10][28] != ele[11][27];
    ele[10][28] != ele[11][28];
    ele[10][28] != ele[11][29];
    ele[10][28] != ele[12][28];
    ele[10][28] != ele[13][28];
    ele[10][28] != ele[14][28];
    ele[10][28] != ele[15][28];
    ele[10][28] != ele[16][28];
    ele[10][28] != ele[17][28];
    ele[10][28] != ele[18][28];
    ele[10][28] != ele[19][28];
    ele[10][28] != ele[20][28];
    ele[10][28] != ele[21][28];
    ele[10][28] != ele[22][28];
    ele[10][28] != ele[23][28];
    ele[10][28] != ele[24][28];
    ele[10][28] != ele[25][28];
    ele[10][28] != ele[26][28];
    ele[10][28] != ele[27][28];
    ele[10][28] != ele[28][28];
    ele[10][28] != ele[29][28];
    ele[10][28] != ele[30][28];
    ele[10][28] != ele[31][28];
    ele[10][28] != ele[32][28];
    ele[10][28] != ele[33][28];
    ele[10][28] != ele[34][28];
    ele[10][28] != ele[35][28];
    ele[10][29] != ele[10][30];
    ele[10][29] != ele[10][31];
    ele[10][29] != ele[10][32];
    ele[10][29] != ele[10][33];
    ele[10][29] != ele[10][34];
    ele[10][29] != ele[10][35];
    ele[10][29] != ele[11][24];
    ele[10][29] != ele[11][25];
    ele[10][29] != ele[11][26];
    ele[10][29] != ele[11][27];
    ele[10][29] != ele[11][28];
    ele[10][29] != ele[11][29];
    ele[10][29] != ele[12][29];
    ele[10][29] != ele[13][29];
    ele[10][29] != ele[14][29];
    ele[10][29] != ele[15][29];
    ele[10][29] != ele[16][29];
    ele[10][29] != ele[17][29];
    ele[10][29] != ele[18][29];
    ele[10][29] != ele[19][29];
    ele[10][29] != ele[20][29];
    ele[10][29] != ele[21][29];
    ele[10][29] != ele[22][29];
    ele[10][29] != ele[23][29];
    ele[10][29] != ele[24][29];
    ele[10][29] != ele[25][29];
    ele[10][29] != ele[26][29];
    ele[10][29] != ele[27][29];
    ele[10][29] != ele[28][29];
    ele[10][29] != ele[29][29];
    ele[10][29] != ele[30][29];
    ele[10][29] != ele[31][29];
    ele[10][29] != ele[32][29];
    ele[10][29] != ele[33][29];
    ele[10][29] != ele[34][29];
    ele[10][29] != ele[35][29];
    ele[10][3] != ele[10][10];
    ele[10][3] != ele[10][11];
    ele[10][3] != ele[10][12];
    ele[10][3] != ele[10][13];
    ele[10][3] != ele[10][14];
    ele[10][3] != ele[10][15];
    ele[10][3] != ele[10][16];
    ele[10][3] != ele[10][17];
    ele[10][3] != ele[10][18];
    ele[10][3] != ele[10][19];
    ele[10][3] != ele[10][20];
    ele[10][3] != ele[10][21];
    ele[10][3] != ele[10][22];
    ele[10][3] != ele[10][23];
    ele[10][3] != ele[10][24];
    ele[10][3] != ele[10][25];
    ele[10][3] != ele[10][26];
    ele[10][3] != ele[10][27];
    ele[10][3] != ele[10][28];
    ele[10][3] != ele[10][29];
    ele[10][3] != ele[10][30];
    ele[10][3] != ele[10][31];
    ele[10][3] != ele[10][32];
    ele[10][3] != ele[10][33];
    ele[10][3] != ele[10][34];
    ele[10][3] != ele[10][35];
    ele[10][3] != ele[10][4];
    ele[10][3] != ele[10][5];
    ele[10][3] != ele[10][6];
    ele[10][3] != ele[10][7];
    ele[10][3] != ele[10][8];
    ele[10][3] != ele[10][9];
    ele[10][3] != ele[11][0];
    ele[10][3] != ele[11][1];
    ele[10][3] != ele[11][2];
    ele[10][3] != ele[11][3];
    ele[10][3] != ele[11][4];
    ele[10][3] != ele[11][5];
    ele[10][3] != ele[12][3];
    ele[10][3] != ele[13][3];
    ele[10][3] != ele[14][3];
    ele[10][3] != ele[15][3];
    ele[10][3] != ele[16][3];
    ele[10][3] != ele[17][3];
    ele[10][3] != ele[18][3];
    ele[10][3] != ele[19][3];
    ele[10][3] != ele[20][3];
    ele[10][3] != ele[21][3];
    ele[10][3] != ele[22][3];
    ele[10][3] != ele[23][3];
    ele[10][3] != ele[24][3];
    ele[10][3] != ele[25][3];
    ele[10][3] != ele[26][3];
    ele[10][3] != ele[27][3];
    ele[10][3] != ele[28][3];
    ele[10][3] != ele[29][3];
    ele[10][3] != ele[30][3];
    ele[10][3] != ele[31][3];
    ele[10][3] != ele[32][3];
    ele[10][3] != ele[33][3];
    ele[10][3] != ele[34][3];
    ele[10][3] != ele[35][3];
    ele[10][30] != ele[10][31];
    ele[10][30] != ele[10][32];
    ele[10][30] != ele[10][33];
    ele[10][30] != ele[10][34];
    ele[10][30] != ele[10][35];
    ele[10][30] != ele[11][30];
    ele[10][30] != ele[11][31];
    ele[10][30] != ele[11][32];
    ele[10][30] != ele[11][33];
    ele[10][30] != ele[11][34];
    ele[10][30] != ele[11][35];
    ele[10][30] != ele[12][30];
    ele[10][30] != ele[13][30];
    ele[10][30] != ele[14][30];
    ele[10][30] != ele[15][30];
    ele[10][30] != ele[16][30];
    ele[10][30] != ele[17][30];
    ele[10][30] != ele[18][30];
    ele[10][30] != ele[19][30];
    ele[10][30] != ele[20][30];
    ele[10][30] != ele[21][30];
    ele[10][30] != ele[22][30];
    ele[10][30] != ele[23][30];
    ele[10][30] != ele[24][30];
    ele[10][30] != ele[25][30];
    ele[10][30] != ele[26][30];
    ele[10][30] != ele[27][30];
    ele[10][30] != ele[28][30];
    ele[10][30] != ele[29][30];
    ele[10][30] != ele[30][30];
    ele[10][30] != ele[31][30];
    ele[10][30] != ele[32][30];
    ele[10][30] != ele[33][30];
    ele[10][30] != ele[34][30];
    ele[10][30] != ele[35][30];
    ele[10][31] != ele[10][32];
    ele[10][31] != ele[10][33];
    ele[10][31] != ele[10][34];
    ele[10][31] != ele[10][35];
    ele[10][31] != ele[11][30];
    ele[10][31] != ele[11][31];
    ele[10][31] != ele[11][32];
    ele[10][31] != ele[11][33];
    ele[10][31] != ele[11][34];
    ele[10][31] != ele[11][35];
    ele[10][31] != ele[12][31];
    ele[10][31] != ele[13][31];
    ele[10][31] != ele[14][31];
    ele[10][31] != ele[15][31];
    ele[10][31] != ele[16][31];
    ele[10][31] != ele[17][31];
    ele[10][31] != ele[18][31];
    ele[10][31] != ele[19][31];
    ele[10][31] != ele[20][31];
    ele[10][31] != ele[21][31];
    ele[10][31] != ele[22][31];
    ele[10][31] != ele[23][31];
    ele[10][31] != ele[24][31];
    ele[10][31] != ele[25][31];
    ele[10][31] != ele[26][31];
    ele[10][31] != ele[27][31];
    ele[10][31] != ele[28][31];
    ele[10][31] != ele[29][31];
    ele[10][31] != ele[30][31];
    ele[10][31] != ele[31][31];
    ele[10][31] != ele[32][31];
    ele[10][31] != ele[33][31];
    ele[10][31] != ele[34][31];
    ele[10][31] != ele[35][31];
    ele[10][32] != ele[10][33];
    ele[10][32] != ele[10][34];
    ele[10][32] != ele[10][35];
    ele[10][32] != ele[11][30];
    ele[10][32] != ele[11][31];
    ele[10][32] != ele[11][32];
    ele[10][32] != ele[11][33];
    ele[10][32] != ele[11][34];
    ele[10][32] != ele[11][35];
    ele[10][32] != ele[12][32];
    ele[10][32] != ele[13][32];
    ele[10][32] != ele[14][32];
    ele[10][32] != ele[15][32];
    ele[10][32] != ele[16][32];
    ele[10][32] != ele[17][32];
    ele[10][32] != ele[18][32];
    ele[10][32] != ele[19][32];
    ele[10][32] != ele[20][32];
    ele[10][32] != ele[21][32];
    ele[10][32] != ele[22][32];
    ele[10][32] != ele[23][32];
    ele[10][32] != ele[24][32];
    ele[10][32] != ele[25][32];
    ele[10][32] != ele[26][32];
    ele[10][32] != ele[27][32];
    ele[10][32] != ele[28][32];
    ele[10][32] != ele[29][32];
    ele[10][32] != ele[30][32];
    ele[10][32] != ele[31][32];
    ele[10][32] != ele[32][32];
    ele[10][32] != ele[33][32];
    ele[10][32] != ele[34][32];
    ele[10][32] != ele[35][32];
    ele[10][33] != ele[10][34];
    ele[10][33] != ele[10][35];
    ele[10][33] != ele[11][30];
    ele[10][33] != ele[11][31];
    ele[10][33] != ele[11][32];
    ele[10][33] != ele[11][33];
    ele[10][33] != ele[11][34];
    ele[10][33] != ele[11][35];
    ele[10][33] != ele[12][33];
    ele[10][33] != ele[13][33];
    ele[10][33] != ele[14][33];
    ele[10][33] != ele[15][33];
    ele[10][33] != ele[16][33];
    ele[10][33] != ele[17][33];
    ele[10][33] != ele[18][33];
    ele[10][33] != ele[19][33];
    ele[10][33] != ele[20][33];
    ele[10][33] != ele[21][33];
    ele[10][33] != ele[22][33];
    ele[10][33] != ele[23][33];
    ele[10][33] != ele[24][33];
    ele[10][33] != ele[25][33];
    ele[10][33] != ele[26][33];
    ele[10][33] != ele[27][33];
    ele[10][33] != ele[28][33];
    ele[10][33] != ele[29][33];
    ele[10][33] != ele[30][33];
    ele[10][33] != ele[31][33];
    ele[10][33] != ele[32][33];
    ele[10][33] != ele[33][33];
    ele[10][33] != ele[34][33];
    ele[10][33] != ele[35][33];
    ele[10][34] != ele[10][35];
    ele[10][34] != ele[11][30];
    ele[10][34] != ele[11][31];
    ele[10][34] != ele[11][32];
    ele[10][34] != ele[11][33];
    ele[10][34] != ele[11][34];
    ele[10][34] != ele[11][35];
    ele[10][34] != ele[12][34];
    ele[10][34] != ele[13][34];
    ele[10][34] != ele[14][34];
    ele[10][34] != ele[15][34];
    ele[10][34] != ele[16][34];
    ele[10][34] != ele[17][34];
    ele[10][34] != ele[18][34];
    ele[10][34] != ele[19][34];
    ele[10][34] != ele[20][34];
    ele[10][34] != ele[21][34];
    ele[10][34] != ele[22][34];
    ele[10][34] != ele[23][34];
    ele[10][34] != ele[24][34];
    ele[10][34] != ele[25][34];
    ele[10][34] != ele[26][34];
    ele[10][34] != ele[27][34];
    ele[10][34] != ele[28][34];
    ele[10][34] != ele[29][34];
    ele[10][34] != ele[30][34];
    ele[10][34] != ele[31][34];
    ele[10][34] != ele[32][34];
    ele[10][34] != ele[33][34];
    ele[10][34] != ele[34][34];
    ele[10][34] != ele[35][34];
    ele[10][35] != ele[11][30];
    ele[10][35] != ele[11][31];
    ele[10][35] != ele[11][32];
    ele[10][35] != ele[11][33];
    ele[10][35] != ele[11][34];
    ele[10][35] != ele[11][35];
    ele[10][35] != ele[12][35];
    ele[10][35] != ele[13][35];
    ele[10][35] != ele[14][35];
    ele[10][35] != ele[15][35];
    ele[10][35] != ele[16][35];
    ele[10][35] != ele[17][35];
    ele[10][35] != ele[18][35];
    ele[10][35] != ele[19][35];
    ele[10][35] != ele[20][35];
    ele[10][35] != ele[21][35];
    ele[10][35] != ele[22][35];
    ele[10][35] != ele[23][35];
    ele[10][35] != ele[24][35];
    ele[10][35] != ele[25][35];
    ele[10][35] != ele[26][35];
    ele[10][35] != ele[27][35];
    ele[10][35] != ele[28][35];
    ele[10][35] != ele[29][35];
    ele[10][35] != ele[30][35];
    ele[10][35] != ele[31][35];
    ele[10][35] != ele[32][35];
    ele[10][35] != ele[33][35];
    ele[10][35] != ele[34][35];
    ele[10][35] != ele[35][35];
    ele[10][4] != ele[10][10];
    ele[10][4] != ele[10][11];
    ele[10][4] != ele[10][12];
    ele[10][4] != ele[10][13];
    ele[10][4] != ele[10][14];
    ele[10][4] != ele[10][15];
    ele[10][4] != ele[10][16];
    ele[10][4] != ele[10][17];
    ele[10][4] != ele[10][18];
    ele[10][4] != ele[10][19];
    ele[10][4] != ele[10][20];
    ele[10][4] != ele[10][21];
    ele[10][4] != ele[10][22];
    ele[10][4] != ele[10][23];
    ele[10][4] != ele[10][24];
    ele[10][4] != ele[10][25];
    ele[10][4] != ele[10][26];
    ele[10][4] != ele[10][27];
    ele[10][4] != ele[10][28];
    ele[10][4] != ele[10][29];
    ele[10][4] != ele[10][30];
    ele[10][4] != ele[10][31];
    ele[10][4] != ele[10][32];
    ele[10][4] != ele[10][33];
    ele[10][4] != ele[10][34];
    ele[10][4] != ele[10][35];
    ele[10][4] != ele[10][5];
    ele[10][4] != ele[10][6];
    ele[10][4] != ele[10][7];
    ele[10][4] != ele[10][8];
    ele[10][4] != ele[10][9];
    ele[10][4] != ele[11][0];
    ele[10][4] != ele[11][1];
    ele[10][4] != ele[11][2];
    ele[10][4] != ele[11][3];
    ele[10][4] != ele[11][4];
    ele[10][4] != ele[11][5];
    ele[10][4] != ele[12][4];
    ele[10][4] != ele[13][4];
    ele[10][4] != ele[14][4];
    ele[10][4] != ele[15][4];
    ele[10][4] != ele[16][4];
    ele[10][4] != ele[17][4];
    ele[10][4] != ele[18][4];
    ele[10][4] != ele[19][4];
    ele[10][4] != ele[20][4];
    ele[10][4] != ele[21][4];
    ele[10][4] != ele[22][4];
    ele[10][4] != ele[23][4];
    ele[10][4] != ele[24][4];
    ele[10][4] != ele[25][4];
    ele[10][4] != ele[26][4];
    ele[10][4] != ele[27][4];
    ele[10][4] != ele[28][4];
    ele[10][4] != ele[29][4];
    ele[10][4] != ele[30][4];
    ele[10][4] != ele[31][4];
    ele[10][4] != ele[32][4];
    ele[10][4] != ele[33][4];
    ele[10][4] != ele[34][4];
    ele[10][4] != ele[35][4];
    ele[10][5] != ele[10][10];
    ele[10][5] != ele[10][11];
    ele[10][5] != ele[10][12];
    ele[10][5] != ele[10][13];
    ele[10][5] != ele[10][14];
    ele[10][5] != ele[10][15];
    ele[10][5] != ele[10][16];
    ele[10][5] != ele[10][17];
    ele[10][5] != ele[10][18];
    ele[10][5] != ele[10][19];
    ele[10][5] != ele[10][20];
    ele[10][5] != ele[10][21];
    ele[10][5] != ele[10][22];
    ele[10][5] != ele[10][23];
    ele[10][5] != ele[10][24];
    ele[10][5] != ele[10][25];
    ele[10][5] != ele[10][26];
    ele[10][5] != ele[10][27];
    ele[10][5] != ele[10][28];
    ele[10][5] != ele[10][29];
    ele[10][5] != ele[10][30];
    ele[10][5] != ele[10][31];
    ele[10][5] != ele[10][32];
    ele[10][5] != ele[10][33];
    ele[10][5] != ele[10][34];
    ele[10][5] != ele[10][35];
    ele[10][5] != ele[10][6];
    ele[10][5] != ele[10][7];
    ele[10][5] != ele[10][8];
    ele[10][5] != ele[10][9];
    ele[10][5] != ele[11][0];
    ele[10][5] != ele[11][1];
    ele[10][5] != ele[11][2];
    ele[10][5] != ele[11][3];
    ele[10][5] != ele[11][4];
    ele[10][5] != ele[11][5];
    ele[10][5] != ele[12][5];
    ele[10][5] != ele[13][5];
    ele[10][5] != ele[14][5];
    ele[10][5] != ele[15][5];
    ele[10][5] != ele[16][5];
    ele[10][5] != ele[17][5];
    ele[10][5] != ele[18][5];
    ele[10][5] != ele[19][5];
    ele[10][5] != ele[20][5];
    ele[10][5] != ele[21][5];
    ele[10][5] != ele[22][5];
    ele[10][5] != ele[23][5];
    ele[10][5] != ele[24][5];
    ele[10][5] != ele[25][5];
    ele[10][5] != ele[26][5];
    ele[10][5] != ele[27][5];
    ele[10][5] != ele[28][5];
    ele[10][5] != ele[29][5];
    ele[10][5] != ele[30][5];
    ele[10][5] != ele[31][5];
    ele[10][5] != ele[32][5];
    ele[10][5] != ele[33][5];
    ele[10][5] != ele[34][5];
    ele[10][5] != ele[35][5];
    ele[10][6] != ele[10][10];
    ele[10][6] != ele[10][11];
    ele[10][6] != ele[10][12];
    ele[10][6] != ele[10][13];
    ele[10][6] != ele[10][14];
    ele[10][6] != ele[10][15];
    ele[10][6] != ele[10][16];
    ele[10][6] != ele[10][17];
    ele[10][6] != ele[10][18];
    ele[10][6] != ele[10][19];
    ele[10][6] != ele[10][20];
    ele[10][6] != ele[10][21];
    ele[10][6] != ele[10][22];
    ele[10][6] != ele[10][23];
    ele[10][6] != ele[10][24];
    ele[10][6] != ele[10][25];
    ele[10][6] != ele[10][26];
    ele[10][6] != ele[10][27];
    ele[10][6] != ele[10][28];
    ele[10][6] != ele[10][29];
    ele[10][6] != ele[10][30];
    ele[10][6] != ele[10][31];
    ele[10][6] != ele[10][32];
    ele[10][6] != ele[10][33];
    ele[10][6] != ele[10][34];
    ele[10][6] != ele[10][35];
    ele[10][6] != ele[10][7];
    ele[10][6] != ele[10][8];
    ele[10][6] != ele[10][9];
    ele[10][6] != ele[11][10];
    ele[10][6] != ele[11][11];
    ele[10][6] != ele[11][6];
    ele[10][6] != ele[11][7];
    ele[10][6] != ele[11][8];
    ele[10][6] != ele[11][9];
    ele[10][6] != ele[12][6];
    ele[10][6] != ele[13][6];
    ele[10][6] != ele[14][6];
    ele[10][6] != ele[15][6];
    ele[10][6] != ele[16][6];
    ele[10][6] != ele[17][6];
    ele[10][6] != ele[18][6];
    ele[10][6] != ele[19][6];
    ele[10][6] != ele[20][6];
    ele[10][6] != ele[21][6];
    ele[10][6] != ele[22][6];
    ele[10][6] != ele[23][6];
    ele[10][6] != ele[24][6];
    ele[10][6] != ele[25][6];
    ele[10][6] != ele[26][6];
    ele[10][6] != ele[27][6];
    ele[10][6] != ele[28][6];
    ele[10][6] != ele[29][6];
    ele[10][6] != ele[30][6];
    ele[10][6] != ele[31][6];
    ele[10][6] != ele[32][6];
    ele[10][6] != ele[33][6];
    ele[10][6] != ele[34][6];
    ele[10][6] != ele[35][6];
    ele[10][7] != ele[10][10];
    ele[10][7] != ele[10][11];
    ele[10][7] != ele[10][12];
    ele[10][7] != ele[10][13];
    ele[10][7] != ele[10][14];
    ele[10][7] != ele[10][15];
    ele[10][7] != ele[10][16];
    ele[10][7] != ele[10][17];
    ele[10][7] != ele[10][18];
    ele[10][7] != ele[10][19];
    ele[10][7] != ele[10][20];
    ele[10][7] != ele[10][21];
    ele[10][7] != ele[10][22];
    ele[10][7] != ele[10][23];
    ele[10][7] != ele[10][24];
    ele[10][7] != ele[10][25];
    ele[10][7] != ele[10][26];
    ele[10][7] != ele[10][27];
    ele[10][7] != ele[10][28];
    ele[10][7] != ele[10][29];
    ele[10][7] != ele[10][30];
    ele[10][7] != ele[10][31];
    ele[10][7] != ele[10][32];
    ele[10][7] != ele[10][33];
    ele[10][7] != ele[10][34];
    ele[10][7] != ele[10][35];
    ele[10][7] != ele[10][8];
    ele[10][7] != ele[10][9];
    ele[10][7] != ele[11][10];
    ele[10][7] != ele[11][11];
    ele[10][7] != ele[11][6];
    ele[10][7] != ele[11][7];
    ele[10][7] != ele[11][8];
    ele[10][7] != ele[11][9];
    ele[10][7] != ele[12][7];
    ele[10][7] != ele[13][7];
    ele[10][7] != ele[14][7];
    ele[10][7] != ele[15][7];
    ele[10][7] != ele[16][7];
    ele[10][7] != ele[17][7];
    ele[10][7] != ele[18][7];
    ele[10][7] != ele[19][7];
    ele[10][7] != ele[20][7];
    ele[10][7] != ele[21][7];
    ele[10][7] != ele[22][7];
    ele[10][7] != ele[23][7];
    ele[10][7] != ele[24][7];
    ele[10][7] != ele[25][7];
    ele[10][7] != ele[26][7];
    ele[10][7] != ele[27][7];
    ele[10][7] != ele[28][7];
    ele[10][7] != ele[29][7];
    ele[10][7] != ele[30][7];
    ele[10][7] != ele[31][7];
    ele[10][7] != ele[32][7];
    ele[10][7] != ele[33][7];
    ele[10][7] != ele[34][7];
    ele[10][7] != ele[35][7];
    ele[10][8] != ele[10][10];
    ele[10][8] != ele[10][11];
    ele[10][8] != ele[10][12];
    ele[10][8] != ele[10][13];
    ele[10][8] != ele[10][14];
    ele[10][8] != ele[10][15];
    ele[10][8] != ele[10][16];
    ele[10][8] != ele[10][17];
    ele[10][8] != ele[10][18];
    ele[10][8] != ele[10][19];
    ele[10][8] != ele[10][20];
    ele[10][8] != ele[10][21];
    ele[10][8] != ele[10][22];
    ele[10][8] != ele[10][23];
    ele[10][8] != ele[10][24];
    ele[10][8] != ele[10][25];
    ele[10][8] != ele[10][26];
    ele[10][8] != ele[10][27];
    ele[10][8] != ele[10][28];
    ele[10][8] != ele[10][29];
    ele[10][8] != ele[10][30];
    ele[10][8] != ele[10][31];
    ele[10][8] != ele[10][32];
    ele[10][8] != ele[10][33];
    ele[10][8] != ele[10][34];
    ele[10][8] != ele[10][35];
    ele[10][8] != ele[10][9];
    ele[10][8] != ele[11][10];
    ele[10][8] != ele[11][11];
    ele[10][8] != ele[11][6];
    ele[10][8] != ele[11][7];
    ele[10][8] != ele[11][8];
    ele[10][8] != ele[11][9];
    ele[10][8] != ele[12][8];
    ele[10][8] != ele[13][8];
    ele[10][8] != ele[14][8];
    ele[10][8] != ele[15][8];
    ele[10][8] != ele[16][8];
    ele[10][8] != ele[17][8];
    ele[10][8] != ele[18][8];
    ele[10][8] != ele[19][8];
    ele[10][8] != ele[20][8];
    ele[10][8] != ele[21][8];
    ele[10][8] != ele[22][8];
    ele[10][8] != ele[23][8];
    ele[10][8] != ele[24][8];
    ele[10][8] != ele[25][8];
    ele[10][8] != ele[26][8];
    ele[10][8] != ele[27][8];
    ele[10][8] != ele[28][8];
    ele[10][8] != ele[29][8];
    ele[10][8] != ele[30][8];
    ele[10][8] != ele[31][8];
    ele[10][8] != ele[32][8];
    ele[10][8] != ele[33][8];
    ele[10][8] != ele[34][8];
    ele[10][8] != ele[35][8];
    ele[10][9] != ele[10][10];
    ele[10][9] != ele[10][11];
    ele[10][9] != ele[10][12];
    ele[10][9] != ele[10][13];
    ele[10][9] != ele[10][14];
    ele[10][9] != ele[10][15];
    ele[10][9] != ele[10][16];
    ele[10][9] != ele[10][17];
    ele[10][9] != ele[10][18];
    ele[10][9] != ele[10][19];
    ele[10][9] != ele[10][20];
    ele[10][9] != ele[10][21];
    ele[10][9] != ele[10][22];
    ele[10][9] != ele[10][23];
    ele[10][9] != ele[10][24];
    ele[10][9] != ele[10][25];
    ele[10][9] != ele[10][26];
    ele[10][9] != ele[10][27];
    ele[10][9] != ele[10][28];
    ele[10][9] != ele[10][29];
    ele[10][9] != ele[10][30];
    ele[10][9] != ele[10][31];
    ele[10][9] != ele[10][32];
    ele[10][9] != ele[10][33];
    ele[10][9] != ele[10][34];
    ele[10][9] != ele[10][35];
    ele[10][9] != ele[11][10];
    ele[10][9] != ele[11][11];
    ele[10][9] != ele[11][6];
    ele[10][9] != ele[11][7];
    ele[10][9] != ele[11][8];
    ele[10][9] != ele[11][9];
    ele[10][9] != ele[12][9];
    ele[10][9] != ele[13][9];
    ele[10][9] != ele[14][9];
    ele[10][9] != ele[15][9];
    ele[10][9] != ele[16][9];
    ele[10][9] != ele[17][9];
    ele[10][9] != ele[18][9];
    ele[10][9] != ele[19][9];
    ele[10][9] != ele[20][9];
    ele[10][9] != ele[21][9];
    ele[10][9] != ele[22][9];
    ele[10][9] != ele[23][9];
    ele[10][9] != ele[24][9];
    ele[10][9] != ele[25][9];
    ele[10][9] != ele[26][9];
    ele[10][9] != ele[27][9];
    ele[10][9] != ele[28][9];
    ele[10][9] != ele[29][9];
    ele[10][9] != ele[30][9];
    ele[10][9] != ele[31][9];
    ele[10][9] != ele[32][9];
    ele[10][9] != ele[33][9];
    ele[10][9] != ele[34][9];
    ele[10][9] != ele[35][9];
    ele[11][0] != ele[11][1];
    ele[11][0] != ele[11][10];
    ele[11][0] != ele[11][11];
    ele[11][0] != ele[11][12];
    ele[11][0] != ele[11][13];
    ele[11][0] != ele[11][14];
    ele[11][0] != ele[11][15];
    ele[11][0] != ele[11][16];
    ele[11][0] != ele[11][17];
    ele[11][0] != ele[11][18];
    ele[11][0] != ele[11][19];
    ele[11][0] != ele[11][2];
    ele[11][0] != ele[11][20];
    ele[11][0] != ele[11][21];
    ele[11][0] != ele[11][22];
    ele[11][0] != ele[11][23];
    ele[11][0] != ele[11][24];
    ele[11][0] != ele[11][25];
    ele[11][0] != ele[11][26];
    ele[11][0] != ele[11][27];
    ele[11][0] != ele[11][28];
    ele[11][0] != ele[11][29];
    ele[11][0] != ele[11][3];
    ele[11][0] != ele[11][30];
    ele[11][0] != ele[11][31];
    ele[11][0] != ele[11][32];
    ele[11][0] != ele[11][33];
    ele[11][0] != ele[11][34];
    ele[11][0] != ele[11][35];
    ele[11][0] != ele[11][4];
    ele[11][0] != ele[11][5];
    ele[11][0] != ele[11][6];
    ele[11][0] != ele[11][7];
    ele[11][0] != ele[11][8];
    ele[11][0] != ele[11][9];
    ele[11][0] != ele[12][0];
    ele[11][0] != ele[13][0];
    ele[11][0] != ele[14][0];
    ele[11][0] != ele[15][0];
    ele[11][0] != ele[16][0];
    ele[11][0] != ele[17][0];
    ele[11][0] != ele[18][0];
    ele[11][0] != ele[19][0];
    ele[11][0] != ele[20][0];
    ele[11][0] != ele[21][0];
    ele[11][0] != ele[22][0];
    ele[11][0] != ele[23][0];
    ele[11][0] != ele[24][0];
    ele[11][0] != ele[25][0];
    ele[11][0] != ele[26][0];
    ele[11][0] != ele[27][0];
    ele[11][0] != ele[28][0];
    ele[11][0] != ele[29][0];
    ele[11][0] != ele[30][0];
    ele[11][0] != ele[31][0];
    ele[11][0] != ele[32][0];
    ele[11][0] != ele[33][0];
    ele[11][0] != ele[34][0];
    ele[11][0] != ele[35][0];
    ele[11][1] != ele[11][10];
    ele[11][1] != ele[11][11];
    ele[11][1] != ele[11][12];
    ele[11][1] != ele[11][13];
    ele[11][1] != ele[11][14];
    ele[11][1] != ele[11][15];
    ele[11][1] != ele[11][16];
    ele[11][1] != ele[11][17];
    ele[11][1] != ele[11][18];
    ele[11][1] != ele[11][19];
    ele[11][1] != ele[11][2];
    ele[11][1] != ele[11][20];
    ele[11][1] != ele[11][21];
    ele[11][1] != ele[11][22];
    ele[11][1] != ele[11][23];
    ele[11][1] != ele[11][24];
    ele[11][1] != ele[11][25];
    ele[11][1] != ele[11][26];
    ele[11][1] != ele[11][27];
    ele[11][1] != ele[11][28];
    ele[11][1] != ele[11][29];
    ele[11][1] != ele[11][3];
    ele[11][1] != ele[11][30];
    ele[11][1] != ele[11][31];
    ele[11][1] != ele[11][32];
    ele[11][1] != ele[11][33];
    ele[11][1] != ele[11][34];
    ele[11][1] != ele[11][35];
    ele[11][1] != ele[11][4];
    ele[11][1] != ele[11][5];
    ele[11][1] != ele[11][6];
    ele[11][1] != ele[11][7];
    ele[11][1] != ele[11][8];
    ele[11][1] != ele[11][9];
    ele[11][1] != ele[12][1];
    ele[11][1] != ele[13][1];
    ele[11][1] != ele[14][1];
    ele[11][1] != ele[15][1];
    ele[11][1] != ele[16][1];
    ele[11][1] != ele[17][1];
    ele[11][1] != ele[18][1];
    ele[11][1] != ele[19][1];
    ele[11][1] != ele[20][1];
    ele[11][1] != ele[21][1];
    ele[11][1] != ele[22][1];
    ele[11][1] != ele[23][1];
    ele[11][1] != ele[24][1];
    ele[11][1] != ele[25][1];
    ele[11][1] != ele[26][1];
    ele[11][1] != ele[27][1];
    ele[11][1] != ele[28][1];
    ele[11][1] != ele[29][1];
    ele[11][1] != ele[30][1];
    ele[11][1] != ele[31][1];
    ele[11][1] != ele[32][1];
    ele[11][1] != ele[33][1];
    ele[11][1] != ele[34][1];
    ele[11][1] != ele[35][1];
    ele[11][10] != ele[11][11];
    ele[11][10] != ele[11][12];
    ele[11][10] != ele[11][13];
    ele[11][10] != ele[11][14];
    ele[11][10] != ele[11][15];
    ele[11][10] != ele[11][16];
    ele[11][10] != ele[11][17];
    ele[11][10] != ele[11][18];
    ele[11][10] != ele[11][19];
    ele[11][10] != ele[11][20];
    ele[11][10] != ele[11][21];
    ele[11][10] != ele[11][22];
    ele[11][10] != ele[11][23];
    ele[11][10] != ele[11][24];
    ele[11][10] != ele[11][25];
    ele[11][10] != ele[11][26];
    ele[11][10] != ele[11][27];
    ele[11][10] != ele[11][28];
    ele[11][10] != ele[11][29];
    ele[11][10] != ele[11][30];
    ele[11][10] != ele[11][31];
    ele[11][10] != ele[11][32];
    ele[11][10] != ele[11][33];
    ele[11][10] != ele[11][34];
    ele[11][10] != ele[11][35];
    ele[11][10] != ele[12][10];
    ele[11][10] != ele[13][10];
    ele[11][10] != ele[14][10];
    ele[11][10] != ele[15][10];
    ele[11][10] != ele[16][10];
    ele[11][10] != ele[17][10];
    ele[11][10] != ele[18][10];
    ele[11][10] != ele[19][10];
    ele[11][10] != ele[20][10];
    ele[11][10] != ele[21][10];
    ele[11][10] != ele[22][10];
    ele[11][10] != ele[23][10];
    ele[11][10] != ele[24][10];
    ele[11][10] != ele[25][10];
    ele[11][10] != ele[26][10];
    ele[11][10] != ele[27][10];
    ele[11][10] != ele[28][10];
    ele[11][10] != ele[29][10];
    ele[11][10] != ele[30][10];
    ele[11][10] != ele[31][10];
    ele[11][10] != ele[32][10];
    ele[11][10] != ele[33][10];
    ele[11][10] != ele[34][10];
    ele[11][10] != ele[35][10];
    ele[11][11] != ele[11][12];
    ele[11][11] != ele[11][13];
    ele[11][11] != ele[11][14];
    ele[11][11] != ele[11][15];
    ele[11][11] != ele[11][16];
    ele[11][11] != ele[11][17];
    ele[11][11] != ele[11][18];
    ele[11][11] != ele[11][19];
    ele[11][11] != ele[11][20];
    ele[11][11] != ele[11][21];
    ele[11][11] != ele[11][22];
    ele[11][11] != ele[11][23];
    ele[11][11] != ele[11][24];
    ele[11][11] != ele[11][25];
    ele[11][11] != ele[11][26];
    ele[11][11] != ele[11][27];
    ele[11][11] != ele[11][28];
    ele[11][11] != ele[11][29];
    ele[11][11] != ele[11][30];
    ele[11][11] != ele[11][31];
    ele[11][11] != ele[11][32];
    ele[11][11] != ele[11][33];
    ele[11][11] != ele[11][34];
    ele[11][11] != ele[11][35];
    ele[11][11] != ele[12][11];
    ele[11][11] != ele[13][11];
    ele[11][11] != ele[14][11];
    ele[11][11] != ele[15][11];
    ele[11][11] != ele[16][11];
    ele[11][11] != ele[17][11];
    ele[11][11] != ele[18][11];
    ele[11][11] != ele[19][11];
    ele[11][11] != ele[20][11];
    ele[11][11] != ele[21][11];
    ele[11][11] != ele[22][11];
    ele[11][11] != ele[23][11];
    ele[11][11] != ele[24][11];
    ele[11][11] != ele[25][11];
    ele[11][11] != ele[26][11];
    ele[11][11] != ele[27][11];
    ele[11][11] != ele[28][11];
    ele[11][11] != ele[29][11];
    ele[11][11] != ele[30][11];
    ele[11][11] != ele[31][11];
    ele[11][11] != ele[32][11];
    ele[11][11] != ele[33][11];
    ele[11][11] != ele[34][11];
    ele[11][11] != ele[35][11];
    ele[11][12] != ele[11][13];
    ele[11][12] != ele[11][14];
    ele[11][12] != ele[11][15];
    ele[11][12] != ele[11][16];
    ele[11][12] != ele[11][17];
    ele[11][12] != ele[11][18];
    ele[11][12] != ele[11][19];
    ele[11][12] != ele[11][20];
    ele[11][12] != ele[11][21];
    ele[11][12] != ele[11][22];
    ele[11][12] != ele[11][23];
    ele[11][12] != ele[11][24];
    ele[11][12] != ele[11][25];
    ele[11][12] != ele[11][26];
    ele[11][12] != ele[11][27];
    ele[11][12] != ele[11][28];
    ele[11][12] != ele[11][29];
    ele[11][12] != ele[11][30];
    ele[11][12] != ele[11][31];
    ele[11][12] != ele[11][32];
    ele[11][12] != ele[11][33];
    ele[11][12] != ele[11][34];
    ele[11][12] != ele[11][35];
    ele[11][12] != ele[12][12];
    ele[11][12] != ele[13][12];
    ele[11][12] != ele[14][12];
    ele[11][12] != ele[15][12];
    ele[11][12] != ele[16][12];
    ele[11][12] != ele[17][12];
    ele[11][12] != ele[18][12];
    ele[11][12] != ele[19][12];
    ele[11][12] != ele[20][12];
    ele[11][12] != ele[21][12];
    ele[11][12] != ele[22][12];
    ele[11][12] != ele[23][12];
    ele[11][12] != ele[24][12];
    ele[11][12] != ele[25][12];
    ele[11][12] != ele[26][12];
    ele[11][12] != ele[27][12];
    ele[11][12] != ele[28][12];
    ele[11][12] != ele[29][12];
    ele[11][12] != ele[30][12];
    ele[11][12] != ele[31][12];
    ele[11][12] != ele[32][12];
    ele[11][12] != ele[33][12];
    ele[11][12] != ele[34][12];
    ele[11][12] != ele[35][12];
    ele[11][13] != ele[11][14];
    ele[11][13] != ele[11][15];
    ele[11][13] != ele[11][16];
    ele[11][13] != ele[11][17];
    ele[11][13] != ele[11][18];
    ele[11][13] != ele[11][19];
    ele[11][13] != ele[11][20];
    ele[11][13] != ele[11][21];
    ele[11][13] != ele[11][22];
    ele[11][13] != ele[11][23];
    ele[11][13] != ele[11][24];
    ele[11][13] != ele[11][25];
    ele[11][13] != ele[11][26];
    ele[11][13] != ele[11][27];
    ele[11][13] != ele[11][28];
    ele[11][13] != ele[11][29];
    ele[11][13] != ele[11][30];
    ele[11][13] != ele[11][31];
    ele[11][13] != ele[11][32];
    ele[11][13] != ele[11][33];
    ele[11][13] != ele[11][34];
    ele[11][13] != ele[11][35];
    ele[11][13] != ele[12][13];
    ele[11][13] != ele[13][13];
    ele[11][13] != ele[14][13];
    ele[11][13] != ele[15][13];
    ele[11][13] != ele[16][13];
    ele[11][13] != ele[17][13];
    ele[11][13] != ele[18][13];
    ele[11][13] != ele[19][13];
    ele[11][13] != ele[20][13];
    ele[11][13] != ele[21][13];
    ele[11][13] != ele[22][13];
    ele[11][13] != ele[23][13];
    ele[11][13] != ele[24][13];
    ele[11][13] != ele[25][13];
    ele[11][13] != ele[26][13];
    ele[11][13] != ele[27][13];
    ele[11][13] != ele[28][13];
    ele[11][13] != ele[29][13];
    ele[11][13] != ele[30][13];
    ele[11][13] != ele[31][13];
    ele[11][13] != ele[32][13];
    ele[11][13] != ele[33][13];
    ele[11][13] != ele[34][13];
    ele[11][13] != ele[35][13];
    ele[11][14] != ele[11][15];
    ele[11][14] != ele[11][16];
    ele[11][14] != ele[11][17];
    ele[11][14] != ele[11][18];
    ele[11][14] != ele[11][19];
    ele[11][14] != ele[11][20];
    ele[11][14] != ele[11][21];
    ele[11][14] != ele[11][22];
    ele[11][14] != ele[11][23];
    ele[11][14] != ele[11][24];
    ele[11][14] != ele[11][25];
    ele[11][14] != ele[11][26];
    ele[11][14] != ele[11][27];
    ele[11][14] != ele[11][28];
    ele[11][14] != ele[11][29];
    ele[11][14] != ele[11][30];
    ele[11][14] != ele[11][31];
    ele[11][14] != ele[11][32];
    ele[11][14] != ele[11][33];
    ele[11][14] != ele[11][34];
    ele[11][14] != ele[11][35];
    ele[11][14] != ele[12][14];
    ele[11][14] != ele[13][14];
    ele[11][14] != ele[14][14];
    ele[11][14] != ele[15][14];
    ele[11][14] != ele[16][14];
    ele[11][14] != ele[17][14];
    ele[11][14] != ele[18][14];
    ele[11][14] != ele[19][14];
    ele[11][14] != ele[20][14];
    ele[11][14] != ele[21][14];
    ele[11][14] != ele[22][14];
    ele[11][14] != ele[23][14];
    ele[11][14] != ele[24][14];
    ele[11][14] != ele[25][14];
    ele[11][14] != ele[26][14];
    ele[11][14] != ele[27][14];
    ele[11][14] != ele[28][14];
    ele[11][14] != ele[29][14];
    ele[11][14] != ele[30][14];
    ele[11][14] != ele[31][14];
    ele[11][14] != ele[32][14];
    ele[11][14] != ele[33][14];
    ele[11][14] != ele[34][14];
    ele[11][14] != ele[35][14];
    ele[11][15] != ele[11][16];
    ele[11][15] != ele[11][17];
    ele[11][15] != ele[11][18];
    ele[11][15] != ele[11][19];
    ele[11][15] != ele[11][20];
    ele[11][15] != ele[11][21];
    ele[11][15] != ele[11][22];
    ele[11][15] != ele[11][23];
    ele[11][15] != ele[11][24];
    ele[11][15] != ele[11][25];
    ele[11][15] != ele[11][26];
    ele[11][15] != ele[11][27];
    ele[11][15] != ele[11][28];
    ele[11][15] != ele[11][29];
    ele[11][15] != ele[11][30];
    ele[11][15] != ele[11][31];
    ele[11][15] != ele[11][32];
    ele[11][15] != ele[11][33];
    ele[11][15] != ele[11][34];
    ele[11][15] != ele[11][35];
    ele[11][15] != ele[12][15];
    ele[11][15] != ele[13][15];
    ele[11][15] != ele[14][15];
    ele[11][15] != ele[15][15];
    ele[11][15] != ele[16][15];
    ele[11][15] != ele[17][15];
    ele[11][15] != ele[18][15];
    ele[11][15] != ele[19][15];
    ele[11][15] != ele[20][15];
    ele[11][15] != ele[21][15];
    ele[11][15] != ele[22][15];
    ele[11][15] != ele[23][15];
    ele[11][15] != ele[24][15];
    ele[11][15] != ele[25][15];
    ele[11][15] != ele[26][15];
    ele[11][15] != ele[27][15];
    ele[11][15] != ele[28][15];
    ele[11][15] != ele[29][15];
    ele[11][15] != ele[30][15];
    ele[11][15] != ele[31][15];
    ele[11][15] != ele[32][15];
    ele[11][15] != ele[33][15];
    ele[11][15] != ele[34][15];
    ele[11][15] != ele[35][15];
    ele[11][16] != ele[11][17];
    ele[11][16] != ele[11][18];
    ele[11][16] != ele[11][19];
    ele[11][16] != ele[11][20];
    ele[11][16] != ele[11][21];
    ele[11][16] != ele[11][22];
    ele[11][16] != ele[11][23];
    ele[11][16] != ele[11][24];
    ele[11][16] != ele[11][25];
    ele[11][16] != ele[11][26];
    ele[11][16] != ele[11][27];
    ele[11][16] != ele[11][28];
    ele[11][16] != ele[11][29];
    ele[11][16] != ele[11][30];
    ele[11][16] != ele[11][31];
    ele[11][16] != ele[11][32];
    ele[11][16] != ele[11][33];
    ele[11][16] != ele[11][34];
    ele[11][16] != ele[11][35];
    ele[11][16] != ele[12][16];
    ele[11][16] != ele[13][16];
    ele[11][16] != ele[14][16];
    ele[11][16] != ele[15][16];
    ele[11][16] != ele[16][16];
    ele[11][16] != ele[17][16];
    ele[11][16] != ele[18][16];
    ele[11][16] != ele[19][16];
    ele[11][16] != ele[20][16];
    ele[11][16] != ele[21][16];
    ele[11][16] != ele[22][16];
    ele[11][16] != ele[23][16];
    ele[11][16] != ele[24][16];
    ele[11][16] != ele[25][16];
    ele[11][16] != ele[26][16];
    ele[11][16] != ele[27][16];
    ele[11][16] != ele[28][16];
    ele[11][16] != ele[29][16];
    ele[11][16] != ele[30][16];
    ele[11][16] != ele[31][16];
    ele[11][16] != ele[32][16];
    ele[11][16] != ele[33][16];
    ele[11][16] != ele[34][16];
    ele[11][16] != ele[35][16];
    ele[11][17] != ele[11][18];
    ele[11][17] != ele[11][19];
    ele[11][17] != ele[11][20];
    ele[11][17] != ele[11][21];
    ele[11][17] != ele[11][22];
    ele[11][17] != ele[11][23];
    ele[11][17] != ele[11][24];
    ele[11][17] != ele[11][25];
    ele[11][17] != ele[11][26];
    ele[11][17] != ele[11][27];
    ele[11][17] != ele[11][28];
    ele[11][17] != ele[11][29];
    ele[11][17] != ele[11][30];
    ele[11][17] != ele[11][31];
    ele[11][17] != ele[11][32];
    ele[11][17] != ele[11][33];
    ele[11][17] != ele[11][34];
    ele[11][17] != ele[11][35];
    ele[11][17] != ele[12][17];
    ele[11][17] != ele[13][17];
    ele[11][17] != ele[14][17];
    ele[11][17] != ele[15][17];
    ele[11][17] != ele[16][17];
    ele[11][17] != ele[17][17];
    ele[11][17] != ele[18][17];
    ele[11][17] != ele[19][17];
    ele[11][17] != ele[20][17];
    ele[11][17] != ele[21][17];
    ele[11][17] != ele[22][17];
    ele[11][17] != ele[23][17];
    ele[11][17] != ele[24][17];
    ele[11][17] != ele[25][17];
    ele[11][17] != ele[26][17];
    ele[11][17] != ele[27][17];
    ele[11][17] != ele[28][17];
    ele[11][17] != ele[29][17];
    ele[11][17] != ele[30][17];
    ele[11][17] != ele[31][17];
    ele[11][17] != ele[32][17];
    ele[11][17] != ele[33][17];
    ele[11][17] != ele[34][17];
    ele[11][17] != ele[35][17];
    ele[11][18] != ele[11][19];
    ele[11][18] != ele[11][20];
    ele[11][18] != ele[11][21];
    ele[11][18] != ele[11][22];
    ele[11][18] != ele[11][23];
    ele[11][18] != ele[11][24];
    ele[11][18] != ele[11][25];
    ele[11][18] != ele[11][26];
    ele[11][18] != ele[11][27];
    ele[11][18] != ele[11][28];
    ele[11][18] != ele[11][29];
    ele[11][18] != ele[11][30];
    ele[11][18] != ele[11][31];
    ele[11][18] != ele[11][32];
    ele[11][18] != ele[11][33];
    ele[11][18] != ele[11][34];
    ele[11][18] != ele[11][35];
    ele[11][18] != ele[12][18];
    ele[11][18] != ele[13][18];
    ele[11][18] != ele[14][18];
    ele[11][18] != ele[15][18];
    ele[11][18] != ele[16][18];
    ele[11][18] != ele[17][18];
    ele[11][18] != ele[18][18];
    ele[11][18] != ele[19][18];
    ele[11][18] != ele[20][18];
    ele[11][18] != ele[21][18];
    ele[11][18] != ele[22][18];
    ele[11][18] != ele[23][18];
    ele[11][18] != ele[24][18];
    ele[11][18] != ele[25][18];
    ele[11][18] != ele[26][18];
    ele[11][18] != ele[27][18];
    ele[11][18] != ele[28][18];
    ele[11][18] != ele[29][18];
    ele[11][18] != ele[30][18];
    ele[11][18] != ele[31][18];
    ele[11][18] != ele[32][18];
    ele[11][18] != ele[33][18];
    ele[11][18] != ele[34][18];
    ele[11][18] != ele[35][18];
    ele[11][19] != ele[11][20];
    ele[11][19] != ele[11][21];
    ele[11][19] != ele[11][22];
    ele[11][19] != ele[11][23];
    ele[11][19] != ele[11][24];
    ele[11][19] != ele[11][25];
    ele[11][19] != ele[11][26];
    ele[11][19] != ele[11][27];
    ele[11][19] != ele[11][28];
    ele[11][19] != ele[11][29];
    ele[11][19] != ele[11][30];
    ele[11][19] != ele[11][31];
    ele[11][19] != ele[11][32];
    ele[11][19] != ele[11][33];
    ele[11][19] != ele[11][34];
    ele[11][19] != ele[11][35];
    ele[11][19] != ele[12][19];
    ele[11][19] != ele[13][19];
    ele[11][19] != ele[14][19];
    ele[11][19] != ele[15][19];
    ele[11][19] != ele[16][19];
    ele[11][19] != ele[17][19];
    ele[11][19] != ele[18][19];
    ele[11][19] != ele[19][19];
    ele[11][19] != ele[20][19];
    ele[11][19] != ele[21][19];
    ele[11][19] != ele[22][19];
    ele[11][19] != ele[23][19];
    ele[11][19] != ele[24][19];
    ele[11][19] != ele[25][19];
    ele[11][19] != ele[26][19];
    ele[11][19] != ele[27][19];
    ele[11][19] != ele[28][19];
    ele[11][19] != ele[29][19];
    ele[11][19] != ele[30][19];
    ele[11][19] != ele[31][19];
    ele[11][19] != ele[32][19];
    ele[11][19] != ele[33][19];
    ele[11][19] != ele[34][19];
    ele[11][19] != ele[35][19];
    ele[11][2] != ele[11][10];
    ele[11][2] != ele[11][11];
    ele[11][2] != ele[11][12];
    ele[11][2] != ele[11][13];
    ele[11][2] != ele[11][14];
    ele[11][2] != ele[11][15];
    ele[11][2] != ele[11][16];
    ele[11][2] != ele[11][17];
    ele[11][2] != ele[11][18];
    ele[11][2] != ele[11][19];
    ele[11][2] != ele[11][20];
    ele[11][2] != ele[11][21];
    ele[11][2] != ele[11][22];
    ele[11][2] != ele[11][23];
    ele[11][2] != ele[11][24];
    ele[11][2] != ele[11][25];
    ele[11][2] != ele[11][26];
    ele[11][2] != ele[11][27];
    ele[11][2] != ele[11][28];
    ele[11][2] != ele[11][29];
    ele[11][2] != ele[11][3];
    ele[11][2] != ele[11][30];
    ele[11][2] != ele[11][31];
    ele[11][2] != ele[11][32];
    ele[11][2] != ele[11][33];
    ele[11][2] != ele[11][34];
    ele[11][2] != ele[11][35];
    ele[11][2] != ele[11][4];
    ele[11][2] != ele[11][5];
    ele[11][2] != ele[11][6];
    ele[11][2] != ele[11][7];
    ele[11][2] != ele[11][8];
    ele[11][2] != ele[11][9];
    ele[11][2] != ele[12][2];
    ele[11][2] != ele[13][2];
    ele[11][2] != ele[14][2];
    ele[11][2] != ele[15][2];
    ele[11][2] != ele[16][2];
    ele[11][2] != ele[17][2];
    ele[11][2] != ele[18][2];
    ele[11][2] != ele[19][2];
    ele[11][2] != ele[20][2];
    ele[11][2] != ele[21][2];
    ele[11][2] != ele[22][2];
    ele[11][2] != ele[23][2];
    ele[11][2] != ele[24][2];
    ele[11][2] != ele[25][2];
    ele[11][2] != ele[26][2];
    ele[11][2] != ele[27][2];
    ele[11][2] != ele[28][2];
    ele[11][2] != ele[29][2];
    ele[11][2] != ele[30][2];
    ele[11][2] != ele[31][2];
    ele[11][2] != ele[32][2];
    ele[11][2] != ele[33][2];
    ele[11][2] != ele[34][2];
    ele[11][2] != ele[35][2];
    ele[11][20] != ele[11][21];
    ele[11][20] != ele[11][22];
    ele[11][20] != ele[11][23];
    ele[11][20] != ele[11][24];
    ele[11][20] != ele[11][25];
    ele[11][20] != ele[11][26];
    ele[11][20] != ele[11][27];
    ele[11][20] != ele[11][28];
    ele[11][20] != ele[11][29];
    ele[11][20] != ele[11][30];
    ele[11][20] != ele[11][31];
    ele[11][20] != ele[11][32];
    ele[11][20] != ele[11][33];
    ele[11][20] != ele[11][34];
    ele[11][20] != ele[11][35];
    ele[11][20] != ele[12][20];
    ele[11][20] != ele[13][20];
    ele[11][20] != ele[14][20];
    ele[11][20] != ele[15][20];
    ele[11][20] != ele[16][20];
    ele[11][20] != ele[17][20];
    ele[11][20] != ele[18][20];
    ele[11][20] != ele[19][20];
    ele[11][20] != ele[20][20];
    ele[11][20] != ele[21][20];
    ele[11][20] != ele[22][20];
    ele[11][20] != ele[23][20];
    ele[11][20] != ele[24][20];
    ele[11][20] != ele[25][20];
    ele[11][20] != ele[26][20];
    ele[11][20] != ele[27][20];
    ele[11][20] != ele[28][20];
    ele[11][20] != ele[29][20];
    ele[11][20] != ele[30][20];
    ele[11][20] != ele[31][20];
    ele[11][20] != ele[32][20];
    ele[11][20] != ele[33][20];
    ele[11][20] != ele[34][20];
    ele[11][20] != ele[35][20];
    ele[11][21] != ele[11][22];
    ele[11][21] != ele[11][23];
    ele[11][21] != ele[11][24];
    ele[11][21] != ele[11][25];
    ele[11][21] != ele[11][26];
    ele[11][21] != ele[11][27];
    ele[11][21] != ele[11][28];
    ele[11][21] != ele[11][29];
    ele[11][21] != ele[11][30];
    ele[11][21] != ele[11][31];
    ele[11][21] != ele[11][32];
    ele[11][21] != ele[11][33];
    ele[11][21] != ele[11][34];
    ele[11][21] != ele[11][35];
    ele[11][21] != ele[12][21];
    ele[11][21] != ele[13][21];
    ele[11][21] != ele[14][21];
    ele[11][21] != ele[15][21];
    ele[11][21] != ele[16][21];
    ele[11][21] != ele[17][21];
    ele[11][21] != ele[18][21];
    ele[11][21] != ele[19][21];
    ele[11][21] != ele[20][21];
    ele[11][21] != ele[21][21];
    ele[11][21] != ele[22][21];
    ele[11][21] != ele[23][21];
    ele[11][21] != ele[24][21];
    ele[11][21] != ele[25][21];
    ele[11][21] != ele[26][21];
    ele[11][21] != ele[27][21];
    ele[11][21] != ele[28][21];
    ele[11][21] != ele[29][21];
    ele[11][21] != ele[30][21];
    ele[11][21] != ele[31][21];
    ele[11][21] != ele[32][21];
    ele[11][21] != ele[33][21];
    ele[11][21] != ele[34][21];
    ele[11][21] != ele[35][21];
    ele[11][22] != ele[11][23];
    ele[11][22] != ele[11][24];
    ele[11][22] != ele[11][25];
    ele[11][22] != ele[11][26];
    ele[11][22] != ele[11][27];
    ele[11][22] != ele[11][28];
    ele[11][22] != ele[11][29];
    ele[11][22] != ele[11][30];
    ele[11][22] != ele[11][31];
    ele[11][22] != ele[11][32];
    ele[11][22] != ele[11][33];
    ele[11][22] != ele[11][34];
    ele[11][22] != ele[11][35];
    ele[11][22] != ele[12][22];
    ele[11][22] != ele[13][22];
    ele[11][22] != ele[14][22];
    ele[11][22] != ele[15][22];
    ele[11][22] != ele[16][22];
    ele[11][22] != ele[17][22];
    ele[11][22] != ele[18][22];
    ele[11][22] != ele[19][22];
    ele[11][22] != ele[20][22];
    ele[11][22] != ele[21][22];
    ele[11][22] != ele[22][22];
    ele[11][22] != ele[23][22];
    ele[11][22] != ele[24][22];
    ele[11][22] != ele[25][22];
    ele[11][22] != ele[26][22];
    ele[11][22] != ele[27][22];
    ele[11][22] != ele[28][22];
    ele[11][22] != ele[29][22];
    ele[11][22] != ele[30][22];
    ele[11][22] != ele[31][22];
    ele[11][22] != ele[32][22];
    ele[11][22] != ele[33][22];
    ele[11][22] != ele[34][22];
    ele[11][22] != ele[35][22];
    ele[11][23] != ele[11][24];
    ele[11][23] != ele[11][25];
    ele[11][23] != ele[11][26];
    ele[11][23] != ele[11][27];
    ele[11][23] != ele[11][28];
    ele[11][23] != ele[11][29];
    ele[11][23] != ele[11][30];
    ele[11][23] != ele[11][31];
    ele[11][23] != ele[11][32];
    ele[11][23] != ele[11][33];
    ele[11][23] != ele[11][34];
    ele[11][23] != ele[11][35];
    ele[11][23] != ele[12][23];
    ele[11][23] != ele[13][23];
    ele[11][23] != ele[14][23];
    ele[11][23] != ele[15][23];
    ele[11][23] != ele[16][23];
    ele[11][23] != ele[17][23];
    ele[11][23] != ele[18][23];
    ele[11][23] != ele[19][23];
    ele[11][23] != ele[20][23];
    ele[11][23] != ele[21][23];
    ele[11][23] != ele[22][23];
    ele[11][23] != ele[23][23];
    ele[11][23] != ele[24][23];
    ele[11][23] != ele[25][23];
    ele[11][23] != ele[26][23];
    ele[11][23] != ele[27][23];
    ele[11][23] != ele[28][23];
    ele[11][23] != ele[29][23];
    ele[11][23] != ele[30][23];
    ele[11][23] != ele[31][23];
    ele[11][23] != ele[32][23];
    ele[11][23] != ele[33][23];
    ele[11][23] != ele[34][23];
    ele[11][23] != ele[35][23];
    ele[11][24] != ele[11][25];
    ele[11][24] != ele[11][26];
    ele[11][24] != ele[11][27];
    ele[11][24] != ele[11][28];
    ele[11][24] != ele[11][29];
    ele[11][24] != ele[11][30];
    ele[11][24] != ele[11][31];
    ele[11][24] != ele[11][32];
    ele[11][24] != ele[11][33];
    ele[11][24] != ele[11][34];
    ele[11][24] != ele[11][35];
    ele[11][24] != ele[12][24];
    ele[11][24] != ele[13][24];
    ele[11][24] != ele[14][24];
    ele[11][24] != ele[15][24];
    ele[11][24] != ele[16][24];
    ele[11][24] != ele[17][24];
    ele[11][24] != ele[18][24];
    ele[11][24] != ele[19][24];
    ele[11][24] != ele[20][24];
    ele[11][24] != ele[21][24];
    ele[11][24] != ele[22][24];
    ele[11][24] != ele[23][24];
    ele[11][24] != ele[24][24];
    ele[11][24] != ele[25][24];
    ele[11][24] != ele[26][24];
    ele[11][24] != ele[27][24];
    ele[11][24] != ele[28][24];
    ele[11][24] != ele[29][24];
    ele[11][24] != ele[30][24];
    ele[11][24] != ele[31][24];
    ele[11][24] != ele[32][24];
    ele[11][24] != ele[33][24];
    ele[11][24] != ele[34][24];
    ele[11][24] != ele[35][24];
    ele[11][25] != ele[11][26];
    ele[11][25] != ele[11][27];
    ele[11][25] != ele[11][28];
    ele[11][25] != ele[11][29];
    ele[11][25] != ele[11][30];
    ele[11][25] != ele[11][31];
    ele[11][25] != ele[11][32];
    ele[11][25] != ele[11][33];
    ele[11][25] != ele[11][34];
    ele[11][25] != ele[11][35];
    ele[11][25] != ele[12][25];
    ele[11][25] != ele[13][25];
    ele[11][25] != ele[14][25];
    ele[11][25] != ele[15][25];
    ele[11][25] != ele[16][25];
    ele[11][25] != ele[17][25];
    ele[11][25] != ele[18][25];
    ele[11][25] != ele[19][25];
    ele[11][25] != ele[20][25];
    ele[11][25] != ele[21][25];
    ele[11][25] != ele[22][25];
    ele[11][25] != ele[23][25];
    ele[11][25] != ele[24][25];
    ele[11][25] != ele[25][25];
    ele[11][25] != ele[26][25];
    ele[11][25] != ele[27][25];
    ele[11][25] != ele[28][25];
    ele[11][25] != ele[29][25];
    ele[11][25] != ele[30][25];
    ele[11][25] != ele[31][25];
    ele[11][25] != ele[32][25];
    ele[11][25] != ele[33][25];
    ele[11][25] != ele[34][25];
    ele[11][25] != ele[35][25];
    ele[11][26] != ele[11][27];
    ele[11][26] != ele[11][28];
    ele[11][26] != ele[11][29];
    ele[11][26] != ele[11][30];
    ele[11][26] != ele[11][31];
    ele[11][26] != ele[11][32];
    ele[11][26] != ele[11][33];
    ele[11][26] != ele[11][34];
    ele[11][26] != ele[11][35];
    ele[11][26] != ele[12][26];
    ele[11][26] != ele[13][26];
    ele[11][26] != ele[14][26];
    ele[11][26] != ele[15][26];
    ele[11][26] != ele[16][26];
    ele[11][26] != ele[17][26];
    ele[11][26] != ele[18][26];
    ele[11][26] != ele[19][26];
    ele[11][26] != ele[20][26];
    ele[11][26] != ele[21][26];
    ele[11][26] != ele[22][26];
    ele[11][26] != ele[23][26];
    ele[11][26] != ele[24][26];
    ele[11][26] != ele[25][26];
    ele[11][26] != ele[26][26];
    ele[11][26] != ele[27][26];
    ele[11][26] != ele[28][26];
    ele[11][26] != ele[29][26];
    ele[11][26] != ele[30][26];
    ele[11][26] != ele[31][26];
    ele[11][26] != ele[32][26];
    ele[11][26] != ele[33][26];
    ele[11][26] != ele[34][26];
    ele[11][26] != ele[35][26];
    ele[11][27] != ele[11][28];
    ele[11][27] != ele[11][29];
    ele[11][27] != ele[11][30];
    ele[11][27] != ele[11][31];
    ele[11][27] != ele[11][32];
    ele[11][27] != ele[11][33];
    ele[11][27] != ele[11][34];
    ele[11][27] != ele[11][35];
    ele[11][27] != ele[12][27];
    ele[11][27] != ele[13][27];
    ele[11][27] != ele[14][27];
    ele[11][27] != ele[15][27];
    ele[11][27] != ele[16][27];
    ele[11][27] != ele[17][27];
    ele[11][27] != ele[18][27];
    ele[11][27] != ele[19][27];
    ele[11][27] != ele[20][27];
    ele[11][27] != ele[21][27];
    ele[11][27] != ele[22][27];
    ele[11][27] != ele[23][27];
    ele[11][27] != ele[24][27];
    ele[11][27] != ele[25][27];
    ele[11][27] != ele[26][27];
    ele[11][27] != ele[27][27];
    ele[11][27] != ele[28][27];
    ele[11][27] != ele[29][27];
    ele[11][27] != ele[30][27];
    ele[11][27] != ele[31][27];
    ele[11][27] != ele[32][27];
    ele[11][27] != ele[33][27];
    ele[11][27] != ele[34][27];
    ele[11][27] != ele[35][27];
    ele[11][28] != ele[11][29];
    ele[11][28] != ele[11][30];
    ele[11][28] != ele[11][31];
    ele[11][28] != ele[11][32];
    ele[11][28] != ele[11][33];
    ele[11][28] != ele[11][34];
    ele[11][28] != ele[11][35];
    ele[11][28] != ele[12][28];
    ele[11][28] != ele[13][28];
    ele[11][28] != ele[14][28];
    ele[11][28] != ele[15][28];
    ele[11][28] != ele[16][28];
    ele[11][28] != ele[17][28];
    ele[11][28] != ele[18][28];
    ele[11][28] != ele[19][28];
    ele[11][28] != ele[20][28];
    ele[11][28] != ele[21][28];
    ele[11][28] != ele[22][28];
    ele[11][28] != ele[23][28];
    ele[11][28] != ele[24][28];
    ele[11][28] != ele[25][28];
    ele[11][28] != ele[26][28];
    ele[11][28] != ele[27][28];
    ele[11][28] != ele[28][28];
    ele[11][28] != ele[29][28];
    ele[11][28] != ele[30][28];
    ele[11][28] != ele[31][28];
    ele[11][28] != ele[32][28];
    ele[11][28] != ele[33][28];
    ele[11][28] != ele[34][28];
    ele[11][28] != ele[35][28];
    ele[11][29] != ele[11][30];
    ele[11][29] != ele[11][31];
    ele[11][29] != ele[11][32];
    ele[11][29] != ele[11][33];
    ele[11][29] != ele[11][34];
    ele[11][29] != ele[11][35];
    ele[11][29] != ele[12][29];
    ele[11][29] != ele[13][29];
    ele[11][29] != ele[14][29];
    ele[11][29] != ele[15][29];
    ele[11][29] != ele[16][29];
    ele[11][29] != ele[17][29];
    ele[11][29] != ele[18][29];
    ele[11][29] != ele[19][29];
    ele[11][29] != ele[20][29];
    ele[11][29] != ele[21][29];
    ele[11][29] != ele[22][29];
    ele[11][29] != ele[23][29];
    ele[11][29] != ele[24][29];
    ele[11][29] != ele[25][29];
    ele[11][29] != ele[26][29];
    ele[11][29] != ele[27][29];
    ele[11][29] != ele[28][29];
    ele[11][29] != ele[29][29];
    ele[11][29] != ele[30][29];
    ele[11][29] != ele[31][29];
    ele[11][29] != ele[32][29];
    ele[11][29] != ele[33][29];
    ele[11][29] != ele[34][29];
    ele[11][29] != ele[35][29];
    ele[11][3] != ele[11][10];
    ele[11][3] != ele[11][11];
    ele[11][3] != ele[11][12];
    ele[11][3] != ele[11][13];
    ele[11][3] != ele[11][14];
    ele[11][3] != ele[11][15];
    ele[11][3] != ele[11][16];
    ele[11][3] != ele[11][17];
    ele[11][3] != ele[11][18];
    ele[11][3] != ele[11][19];
    ele[11][3] != ele[11][20];
    ele[11][3] != ele[11][21];
    ele[11][3] != ele[11][22];
    ele[11][3] != ele[11][23];
    ele[11][3] != ele[11][24];
    ele[11][3] != ele[11][25];
    ele[11][3] != ele[11][26];
    ele[11][3] != ele[11][27];
    ele[11][3] != ele[11][28];
    ele[11][3] != ele[11][29];
    ele[11][3] != ele[11][30];
    ele[11][3] != ele[11][31];
    ele[11][3] != ele[11][32];
    ele[11][3] != ele[11][33];
    ele[11][3] != ele[11][34];
    ele[11][3] != ele[11][35];
    ele[11][3] != ele[11][4];
    ele[11][3] != ele[11][5];
    ele[11][3] != ele[11][6];
    ele[11][3] != ele[11][7];
    ele[11][3] != ele[11][8];
    ele[11][3] != ele[11][9];
    ele[11][3] != ele[12][3];
    ele[11][3] != ele[13][3];
    ele[11][3] != ele[14][3];
    ele[11][3] != ele[15][3];
    ele[11][3] != ele[16][3];
    ele[11][3] != ele[17][3];
    ele[11][3] != ele[18][3];
    ele[11][3] != ele[19][3];
    ele[11][3] != ele[20][3];
    ele[11][3] != ele[21][3];
    ele[11][3] != ele[22][3];
    ele[11][3] != ele[23][3];
    ele[11][3] != ele[24][3];
    ele[11][3] != ele[25][3];
    ele[11][3] != ele[26][3];
    ele[11][3] != ele[27][3];
    ele[11][3] != ele[28][3];
    ele[11][3] != ele[29][3];
    ele[11][3] != ele[30][3];
    ele[11][3] != ele[31][3];
    ele[11][3] != ele[32][3];
    ele[11][3] != ele[33][3];
    ele[11][3] != ele[34][3];
    ele[11][3] != ele[35][3];
    ele[11][30] != ele[11][31];
    ele[11][30] != ele[11][32];
    ele[11][30] != ele[11][33];
    ele[11][30] != ele[11][34];
    ele[11][30] != ele[11][35];
    ele[11][30] != ele[12][30];
    ele[11][30] != ele[13][30];
    ele[11][30] != ele[14][30];
    ele[11][30] != ele[15][30];
    ele[11][30] != ele[16][30];
    ele[11][30] != ele[17][30];
    ele[11][30] != ele[18][30];
    ele[11][30] != ele[19][30];
    ele[11][30] != ele[20][30];
    ele[11][30] != ele[21][30];
    ele[11][30] != ele[22][30];
    ele[11][30] != ele[23][30];
    ele[11][30] != ele[24][30];
    ele[11][30] != ele[25][30];
    ele[11][30] != ele[26][30];
    ele[11][30] != ele[27][30];
    ele[11][30] != ele[28][30];
    ele[11][30] != ele[29][30];
    ele[11][30] != ele[30][30];
    ele[11][30] != ele[31][30];
    ele[11][30] != ele[32][30];
    ele[11][30] != ele[33][30];
    ele[11][30] != ele[34][30];
    ele[11][30] != ele[35][30];
    ele[11][31] != ele[11][32];
    ele[11][31] != ele[11][33];
    ele[11][31] != ele[11][34];
    ele[11][31] != ele[11][35];
    ele[11][31] != ele[12][31];
    ele[11][31] != ele[13][31];
    ele[11][31] != ele[14][31];
    ele[11][31] != ele[15][31];
    ele[11][31] != ele[16][31];
    ele[11][31] != ele[17][31];
    ele[11][31] != ele[18][31];
    ele[11][31] != ele[19][31];
    ele[11][31] != ele[20][31];
    ele[11][31] != ele[21][31];
    ele[11][31] != ele[22][31];
    ele[11][31] != ele[23][31];
    ele[11][31] != ele[24][31];
    ele[11][31] != ele[25][31];
    ele[11][31] != ele[26][31];
    ele[11][31] != ele[27][31];
    ele[11][31] != ele[28][31];
    ele[11][31] != ele[29][31];
    ele[11][31] != ele[30][31];
    ele[11][31] != ele[31][31];
    ele[11][31] != ele[32][31];
    ele[11][31] != ele[33][31];
    ele[11][31] != ele[34][31];
    ele[11][31] != ele[35][31];
    ele[11][32] != ele[11][33];
    ele[11][32] != ele[11][34];
    ele[11][32] != ele[11][35];
    ele[11][32] != ele[12][32];
    ele[11][32] != ele[13][32];
    ele[11][32] != ele[14][32];
    ele[11][32] != ele[15][32];
    ele[11][32] != ele[16][32];
    ele[11][32] != ele[17][32];
    ele[11][32] != ele[18][32];
    ele[11][32] != ele[19][32];
    ele[11][32] != ele[20][32];
    ele[11][32] != ele[21][32];
    ele[11][32] != ele[22][32];
    ele[11][32] != ele[23][32];
    ele[11][32] != ele[24][32];
    ele[11][32] != ele[25][32];
    ele[11][32] != ele[26][32];
    ele[11][32] != ele[27][32];
    ele[11][32] != ele[28][32];
    ele[11][32] != ele[29][32];
    ele[11][32] != ele[30][32];
    ele[11][32] != ele[31][32];
    ele[11][32] != ele[32][32];
    ele[11][32] != ele[33][32];
    ele[11][32] != ele[34][32];
    ele[11][32] != ele[35][32];
    ele[11][33] != ele[11][34];
    ele[11][33] != ele[11][35];
    ele[11][33] != ele[12][33];
    ele[11][33] != ele[13][33];
    ele[11][33] != ele[14][33];
    ele[11][33] != ele[15][33];
    ele[11][33] != ele[16][33];
    ele[11][33] != ele[17][33];
    ele[11][33] != ele[18][33];
    ele[11][33] != ele[19][33];
    ele[11][33] != ele[20][33];
    ele[11][33] != ele[21][33];
    ele[11][33] != ele[22][33];
    ele[11][33] != ele[23][33];
    ele[11][33] != ele[24][33];
    ele[11][33] != ele[25][33];
    ele[11][33] != ele[26][33];
    ele[11][33] != ele[27][33];
    ele[11][33] != ele[28][33];
    ele[11][33] != ele[29][33];
    ele[11][33] != ele[30][33];
    ele[11][33] != ele[31][33];
    ele[11][33] != ele[32][33];
    ele[11][33] != ele[33][33];
    ele[11][33] != ele[34][33];
    ele[11][33] != ele[35][33];
    ele[11][34] != ele[11][35];
    ele[11][34] != ele[12][34];
    ele[11][34] != ele[13][34];
    ele[11][34] != ele[14][34];
    ele[11][34] != ele[15][34];
    ele[11][34] != ele[16][34];
    ele[11][34] != ele[17][34];
    ele[11][34] != ele[18][34];
    ele[11][34] != ele[19][34];
    ele[11][34] != ele[20][34];
    ele[11][34] != ele[21][34];
    ele[11][34] != ele[22][34];
    ele[11][34] != ele[23][34];
    ele[11][34] != ele[24][34];
    ele[11][34] != ele[25][34];
    ele[11][34] != ele[26][34];
    ele[11][34] != ele[27][34];
    ele[11][34] != ele[28][34];
    ele[11][34] != ele[29][34];
    ele[11][34] != ele[30][34];
    ele[11][34] != ele[31][34];
    ele[11][34] != ele[32][34];
    ele[11][34] != ele[33][34];
    ele[11][34] != ele[34][34];
    ele[11][34] != ele[35][34];
    ele[11][35] != ele[12][35];
    ele[11][35] != ele[13][35];
    ele[11][35] != ele[14][35];
    ele[11][35] != ele[15][35];
    ele[11][35] != ele[16][35];
    ele[11][35] != ele[17][35];
    ele[11][35] != ele[18][35];
    ele[11][35] != ele[19][35];
    ele[11][35] != ele[20][35];
    ele[11][35] != ele[21][35];
    ele[11][35] != ele[22][35];
    ele[11][35] != ele[23][35];
    ele[11][35] != ele[24][35];
    ele[11][35] != ele[25][35];
    ele[11][35] != ele[26][35];
    ele[11][35] != ele[27][35];
    ele[11][35] != ele[28][35];
    ele[11][35] != ele[29][35];
    ele[11][35] != ele[30][35];
    ele[11][35] != ele[31][35];
    ele[11][35] != ele[32][35];
    ele[11][35] != ele[33][35];
    ele[11][35] != ele[34][35];
    ele[11][35] != ele[35][35];
    ele[11][4] != ele[11][10];
    ele[11][4] != ele[11][11];
    ele[11][4] != ele[11][12];
    ele[11][4] != ele[11][13];
    ele[11][4] != ele[11][14];
    ele[11][4] != ele[11][15];
    ele[11][4] != ele[11][16];
    ele[11][4] != ele[11][17];
    ele[11][4] != ele[11][18];
    ele[11][4] != ele[11][19];
    ele[11][4] != ele[11][20];
    ele[11][4] != ele[11][21];
    ele[11][4] != ele[11][22];
    ele[11][4] != ele[11][23];
    ele[11][4] != ele[11][24];
    ele[11][4] != ele[11][25];
    ele[11][4] != ele[11][26];
    ele[11][4] != ele[11][27];
    ele[11][4] != ele[11][28];
    ele[11][4] != ele[11][29];
    ele[11][4] != ele[11][30];
    ele[11][4] != ele[11][31];
    ele[11][4] != ele[11][32];
    ele[11][4] != ele[11][33];
    ele[11][4] != ele[11][34];
    ele[11][4] != ele[11][35];
    ele[11][4] != ele[11][5];
    ele[11][4] != ele[11][6];
    ele[11][4] != ele[11][7];
    ele[11][4] != ele[11][8];
    ele[11][4] != ele[11][9];
    ele[11][4] != ele[12][4];
    ele[11][4] != ele[13][4];
    ele[11][4] != ele[14][4];
    ele[11][4] != ele[15][4];
    ele[11][4] != ele[16][4];
    ele[11][4] != ele[17][4];
    ele[11][4] != ele[18][4];
    ele[11][4] != ele[19][4];
    ele[11][4] != ele[20][4];
    ele[11][4] != ele[21][4];
    ele[11][4] != ele[22][4];
    ele[11][4] != ele[23][4];
    ele[11][4] != ele[24][4];
    ele[11][4] != ele[25][4];
    ele[11][4] != ele[26][4];
    ele[11][4] != ele[27][4];
    ele[11][4] != ele[28][4];
    ele[11][4] != ele[29][4];
    ele[11][4] != ele[30][4];
    ele[11][4] != ele[31][4];
    ele[11][4] != ele[32][4];
    ele[11][4] != ele[33][4];
    ele[11][4] != ele[34][4];
    ele[11][4] != ele[35][4];
    ele[11][5] != ele[11][10];
    ele[11][5] != ele[11][11];
    ele[11][5] != ele[11][12];
    ele[11][5] != ele[11][13];
    ele[11][5] != ele[11][14];
    ele[11][5] != ele[11][15];
    ele[11][5] != ele[11][16];
    ele[11][5] != ele[11][17];
    ele[11][5] != ele[11][18];
    ele[11][5] != ele[11][19];
    ele[11][5] != ele[11][20];
    ele[11][5] != ele[11][21];
    ele[11][5] != ele[11][22];
    ele[11][5] != ele[11][23];
    ele[11][5] != ele[11][24];
    ele[11][5] != ele[11][25];
    ele[11][5] != ele[11][26];
    ele[11][5] != ele[11][27];
    ele[11][5] != ele[11][28];
    ele[11][5] != ele[11][29];
    ele[11][5] != ele[11][30];
    ele[11][5] != ele[11][31];
    ele[11][5] != ele[11][32];
    ele[11][5] != ele[11][33];
    ele[11][5] != ele[11][34];
    ele[11][5] != ele[11][35];
    ele[11][5] != ele[11][6];
    ele[11][5] != ele[11][7];
    ele[11][5] != ele[11][8];
    ele[11][5] != ele[11][9];
    ele[11][5] != ele[12][5];
    ele[11][5] != ele[13][5];
    ele[11][5] != ele[14][5];
    ele[11][5] != ele[15][5];
    ele[11][5] != ele[16][5];
    ele[11][5] != ele[17][5];
    ele[11][5] != ele[18][5];
    ele[11][5] != ele[19][5];
    ele[11][5] != ele[20][5];
    ele[11][5] != ele[21][5];
    ele[11][5] != ele[22][5];
    ele[11][5] != ele[23][5];
    ele[11][5] != ele[24][5];
    ele[11][5] != ele[25][5];
    ele[11][5] != ele[26][5];
    ele[11][5] != ele[27][5];
    ele[11][5] != ele[28][5];
    ele[11][5] != ele[29][5];
    ele[11][5] != ele[30][5];
    ele[11][5] != ele[31][5];
    ele[11][5] != ele[32][5];
    ele[11][5] != ele[33][5];
    ele[11][5] != ele[34][5];
    ele[11][5] != ele[35][5];
    ele[11][6] != ele[11][10];
    ele[11][6] != ele[11][11];
    ele[11][6] != ele[11][12];
    ele[11][6] != ele[11][13];
    ele[11][6] != ele[11][14];
    ele[11][6] != ele[11][15];
    ele[11][6] != ele[11][16];
    ele[11][6] != ele[11][17];
    ele[11][6] != ele[11][18];
    ele[11][6] != ele[11][19];
    ele[11][6] != ele[11][20];
    ele[11][6] != ele[11][21];
    ele[11][6] != ele[11][22];
    ele[11][6] != ele[11][23];
    ele[11][6] != ele[11][24];
    ele[11][6] != ele[11][25];
    ele[11][6] != ele[11][26];
    ele[11][6] != ele[11][27];
    ele[11][6] != ele[11][28];
    ele[11][6] != ele[11][29];
    ele[11][6] != ele[11][30];
    ele[11][6] != ele[11][31];
    ele[11][6] != ele[11][32];
    ele[11][6] != ele[11][33];
    ele[11][6] != ele[11][34];
    ele[11][6] != ele[11][35];
    ele[11][6] != ele[11][7];
    ele[11][6] != ele[11][8];
    ele[11][6] != ele[11][9];
    ele[11][6] != ele[12][6];
    ele[11][6] != ele[13][6];
    ele[11][6] != ele[14][6];
    ele[11][6] != ele[15][6];
    ele[11][6] != ele[16][6];
    ele[11][6] != ele[17][6];
    ele[11][6] != ele[18][6];
    ele[11][6] != ele[19][6];
    ele[11][6] != ele[20][6];
    ele[11][6] != ele[21][6];
    ele[11][6] != ele[22][6];
    ele[11][6] != ele[23][6];
    ele[11][6] != ele[24][6];
    ele[11][6] != ele[25][6];
    ele[11][6] != ele[26][6];
    ele[11][6] != ele[27][6];
    ele[11][6] != ele[28][6];
    ele[11][6] != ele[29][6];
    ele[11][6] != ele[30][6];
    ele[11][6] != ele[31][6];
    ele[11][6] != ele[32][6];
    ele[11][6] != ele[33][6];
    ele[11][6] != ele[34][6];
    ele[11][6] != ele[35][6];
    ele[11][7] != ele[11][10];
    ele[11][7] != ele[11][11];
    ele[11][7] != ele[11][12];
    ele[11][7] != ele[11][13];
    ele[11][7] != ele[11][14];
    ele[11][7] != ele[11][15];
    ele[11][7] != ele[11][16];
    ele[11][7] != ele[11][17];
    ele[11][7] != ele[11][18];
    ele[11][7] != ele[11][19];
    ele[11][7] != ele[11][20];
    ele[11][7] != ele[11][21];
    ele[11][7] != ele[11][22];
    ele[11][7] != ele[11][23];
    ele[11][7] != ele[11][24];
    ele[11][7] != ele[11][25];
    ele[11][7] != ele[11][26];
    ele[11][7] != ele[11][27];
    ele[11][7] != ele[11][28];
    ele[11][7] != ele[11][29];
    ele[11][7] != ele[11][30];
    ele[11][7] != ele[11][31];
    ele[11][7] != ele[11][32];
    ele[11][7] != ele[11][33];
    ele[11][7] != ele[11][34];
    ele[11][7] != ele[11][35];
    ele[11][7] != ele[11][8];
    ele[11][7] != ele[11][9];
    ele[11][7] != ele[12][7];
    ele[11][7] != ele[13][7];
    ele[11][7] != ele[14][7];
    ele[11][7] != ele[15][7];
    ele[11][7] != ele[16][7];
    ele[11][7] != ele[17][7];
    ele[11][7] != ele[18][7];
    ele[11][7] != ele[19][7];
    ele[11][7] != ele[20][7];
    ele[11][7] != ele[21][7];
    ele[11][7] != ele[22][7];
    ele[11][7] != ele[23][7];
    ele[11][7] != ele[24][7];
    ele[11][7] != ele[25][7];
    ele[11][7] != ele[26][7];
    ele[11][7] != ele[27][7];
    ele[11][7] != ele[28][7];
    ele[11][7] != ele[29][7];
    ele[11][7] != ele[30][7];
    ele[11][7] != ele[31][7];
    ele[11][7] != ele[32][7];
    ele[11][7] != ele[33][7];
    ele[11][7] != ele[34][7];
    ele[11][7] != ele[35][7];
    ele[11][8] != ele[11][10];
    ele[11][8] != ele[11][11];
    ele[11][8] != ele[11][12];
    ele[11][8] != ele[11][13];
    ele[11][8] != ele[11][14];
    ele[11][8] != ele[11][15];
    ele[11][8] != ele[11][16];
    ele[11][8] != ele[11][17];
    ele[11][8] != ele[11][18];
    ele[11][8] != ele[11][19];
    ele[11][8] != ele[11][20];
    ele[11][8] != ele[11][21];
    ele[11][8] != ele[11][22];
    ele[11][8] != ele[11][23];
    ele[11][8] != ele[11][24];
    ele[11][8] != ele[11][25];
    ele[11][8] != ele[11][26];
    ele[11][8] != ele[11][27];
    ele[11][8] != ele[11][28];
    ele[11][8] != ele[11][29];
    ele[11][8] != ele[11][30];
    ele[11][8] != ele[11][31];
    ele[11][8] != ele[11][32];
    ele[11][8] != ele[11][33];
    ele[11][8] != ele[11][34];
    ele[11][8] != ele[11][35];
    ele[11][8] != ele[11][9];
    ele[11][8] != ele[12][8];
    ele[11][8] != ele[13][8];
    ele[11][8] != ele[14][8];
    ele[11][8] != ele[15][8];
    ele[11][8] != ele[16][8];
    ele[11][8] != ele[17][8];
    ele[11][8] != ele[18][8];
    ele[11][8] != ele[19][8];
    ele[11][8] != ele[20][8];
    ele[11][8] != ele[21][8];
    ele[11][8] != ele[22][8];
    ele[11][8] != ele[23][8];
    ele[11][8] != ele[24][8];
    ele[11][8] != ele[25][8];
    ele[11][8] != ele[26][8];
    ele[11][8] != ele[27][8];
    ele[11][8] != ele[28][8];
    ele[11][8] != ele[29][8];
    ele[11][8] != ele[30][8];
    ele[11][8] != ele[31][8];
    ele[11][8] != ele[32][8];
    ele[11][8] != ele[33][8];
    ele[11][8] != ele[34][8];
    ele[11][8] != ele[35][8];
    ele[11][9] != ele[11][10];
    ele[11][9] != ele[11][11];
    ele[11][9] != ele[11][12];
    ele[11][9] != ele[11][13];
    ele[11][9] != ele[11][14];
    ele[11][9] != ele[11][15];
    ele[11][9] != ele[11][16];
    ele[11][9] != ele[11][17];
    ele[11][9] != ele[11][18];
    ele[11][9] != ele[11][19];
    ele[11][9] != ele[11][20];
    ele[11][9] != ele[11][21];
    ele[11][9] != ele[11][22];
    ele[11][9] != ele[11][23];
    ele[11][9] != ele[11][24];
    ele[11][9] != ele[11][25];
    ele[11][9] != ele[11][26];
    ele[11][9] != ele[11][27];
    ele[11][9] != ele[11][28];
    ele[11][9] != ele[11][29];
    ele[11][9] != ele[11][30];
    ele[11][9] != ele[11][31];
    ele[11][9] != ele[11][32];
    ele[11][9] != ele[11][33];
    ele[11][9] != ele[11][34];
    ele[11][9] != ele[11][35];
    ele[11][9] != ele[12][9];
    ele[11][9] != ele[13][9];
    ele[11][9] != ele[14][9];
    ele[11][9] != ele[15][9];
    ele[11][9] != ele[16][9];
    ele[11][9] != ele[17][9];
    ele[11][9] != ele[18][9];
    ele[11][9] != ele[19][9];
    ele[11][9] != ele[20][9];
    ele[11][9] != ele[21][9];
    ele[11][9] != ele[22][9];
    ele[11][9] != ele[23][9];
    ele[11][9] != ele[24][9];
    ele[11][9] != ele[25][9];
    ele[11][9] != ele[26][9];
    ele[11][9] != ele[27][9];
    ele[11][9] != ele[28][9];
    ele[11][9] != ele[29][9];
    ele[11][9] != ele[30][9];
    ele[11][9] != ele[31][9];
    ele[11][9] != ele[32][9];
    ele[11][9] != ele[33][9];
    ele[11][9] != ele[34][9];
    ele[11][9] != ele[35][9];
    ele[12][0] != ele[12][1];
    ele[12][0] != ele[12][10];
    ele[12][0] != ele[12][11];
    ele[12][0] != ele[12][12];
    ele[12][0] != ele[12][13];
    ele[12][0] != ele[12][14];
    ele[12][0] != ele[12][15];
    ele[12][0] != ele[12][16];
    ele[12][0] != ele[12][17];
    ele[12][0] != ele[12][18];
    ele[12][0] != ele[12][19];
    ele[12][0] != ele[12][2];
    ele[12][0] != ele[12][20];
    ele[12][0] != ele[12][21];
    ele[12][0] != ele[12][22];
    ele[12][0] != ele[12][23];
    ele[12][0] != ele[12][24];
    ele[12][0] != ele[12][25];
    ele[12][0] != ele[12][26];
    ele[12][0] != ele[12][27];
    ele[12][0] != ele[12][28];
    ele[12][0] != ele[12][29];
    ele[12][0] != ele[12][3];
    ele[12][0] != ele[12][30];
    ele[12][0] != ele[12][31];
    ele[12][0] != ele[12][32];
    ele[12][0] != ele[12][33];
    ele[12][0] != ele[12][34];
    ele[12][0] != ele[12][35];
    ele[12][0] != ele[12][4];
    ele[12][0] != ele[12][5];
    ele[12][0] != ele[12][6];
    ele[12][0] != ele[12][7];
    ele[12][0] != ele[12][8];
    ele[12][0] != ele[12][9];
    ele[12][0] != ele[13][0];
    ele[12][0] != ele[13][1];
    ele[12][0] != ele[13][2];
    ele[12][0] != ele[13][3];
    ele[12][0] != ele[13][4];
    ele[12][0] != ele[13][5];
    ele[12][0] != ele[14][0];
    ele[12][0] != ele[14][1];
    ele[12][0] != ele[14][2];
    ele[12][0] != ele[14][3];
    ele[12][0] != ele[14][4];
    ele[12][0] != ele[14][5];
    ele[12][0] != ele[15][0];
    ele[12][0] != ele[15][1];
    ele[12][0] != ele[15][2];
    ele[12][0] != ele[15][3];
    ele[12][0] != ele[15][4];
    ele[12][0] != ele[15][5];
    ele[12][0] != ele[16][0];
    ele[12][0] != ele[16][1];
    ele[12][0] != ele[16][2];
    ele[12][0] != ele[16][3];
    ele[12][0] != ele[16][4];
    ele[12][0] != ele[16][5];
    ele[12][0] != ele[17][0];
    ele[12][0] != ele[17][1];
    ele[12][0] != ele[17][2];
    ele[12][0] != ele[17][3];
    ele[12][0] != ele[17][4];
    ele[12][0] != ele[17][5];
    ele[12][0] != ele[18][0];
    ele[12][0] != ele[19][0];
    ele[12][0] != ele[20][0];
    ele[12][0] != ele[21][0];
    ele[12][0] != ele[22][0];
    ele[12][0] != ele[23][0];
    ele[12][0] != ele[24][0];
    ele[12][0] != ele[25][0];
    ele[12][0] != ele[26][0];
    ele[12][0] != ele[27][0];
    ele[12][0] != ele[28][0];
    ele[12][0] != ele[29][0];
    ele[12][0] != ele[30][0];
    ele[12][0] != ele[31][0];
    ele[12][0] != ele[32][0];
    ele[12][0] != ele[33][0];
    ele[12][0] != ele[34][0];
    ele[12][0] != ele[35][0];
    ele[12][1] != ele[12][10];
    ele[12][1] != ele[12][11];
    ele[12][1] != ele[12][12];
    ele[12][1] != ele[12][13];
    ele[12][1] != ele[12][14];
    ele[12][1] != ele[12][15];
    ele[12][1] != ele[12][16];
    ele[12][1] != ele[12][17];
    ele[12][1] != ele[12][18];
    ele[12][1] != ele[12][19];
    ele[12][1] != ele[12][2];
    ele[12][1] != ele[12][20];
    ele[12][1] != ele[12][21];
    ele[12][1] != ele[12][22];
    ele[12][1] != ele[12][23];
    ele[12][1] != ele[12][24];
    ele[12][1] != ele[12][25];
    ele[12][1] != ele[12][26];
    ele[12][1] != ele[12][27];
    ele[12][1] != ele[12][28];
    ele[12][1] != ele[12][29];
    ele[12][1] != ele[12][3];
    ele[12][1] != ele[12][30];
    ele[12][1] != ele[12][31];
    ele[12][1] != ele[12][32];
    ele[12][1] != ele[12][33];
    ele[12][1] != ele[12][34];
    ele[12][1] != ele[12][35];
    ele[12][1] != ele[12][4];
    ele[12][1] != ele[12][5];
    ele[12][1] != ele[12][6];
    ele[12][1] != ele[12][7];
    ele[12][1] != ele[12][8];
    ele[12][1] != ele[12][9];
    ele[12][1] != ele[13][0];
    ele[12][1] != ele[13][1];
    ele[12][1] != ele[13][2];
    ele[12][1] != ele[13][3];
    ele[12][1] != ele[13][4];
    ele[12][1] != ele[13][5];
    ele[12][1] != ele[14][0];
    ele[12][1] != ele[14][1];
    ele[12][1] != ele[14][2];
    ele[12][1] != ele[14][3];
    ele[12][1] != ele[14][4];
    ele[12][1] != ele[14][5];
    ele[12][1] != ele[15][0];
    ele[12][1] != ele[15][1];
    ele[12][1] != ele[15][2];
    ele[12][1] != ele[15][3];
    ele[12][1] != ele[15][4];
    ele[12][1] != ele[15][5];
    ele[12][1] != ele[16][0];
    ele[12][1] != ele[16][1];
    ele[12][1] != ele[16][2];
    ele[12][1] != ele[16][3];
    ele[12][1] != ele[16][4];
    ele[12][1] != ele[16][5];
    ele[12][1] != ele[17][0];
    ele[12][1] != ele[17][1];
    ele[12][1] != ele[17][2];
    ele[12][1] != ele[17][3];
    ele[12][1] != ele[17][4];
    ele[12][1] != ele[17][5];
    ele[12][1] != ele[18][1];
    ele[12][1] != ele[19][1];
    ele[12][1] != ele[20][1];
    ele[12][1] != ele[21][1];
    ele[12][1] != ele[22][1];
    ele[12][1] != ele[23][1];
    ele[12][1] != ele[24][1];
    ele[12][1] != ele[25][1];
    ele[12][1] != ele[26][1];
    ele[12][1] != ele[27][1];
    ele[12][1] != ele[28][1];
    ele[12][1] != ele[29][1];
    ele[12][1] != ele[30][1];
    ele[12][1] != ele[31][1];
    ele[12][1] != ele[32][1];
    ele[12][1] != ele[33][1];
    ele[12][1] != ele[34][1];
    ele[12][1] != ele[35][1];
    ele[12][10] != ele[12][11];
    ele[12][10] != ele[12][12];
    ele[12][10] != ele[12][13];
    ele[12][10] != ele[12][14];
    ele[12][10] != ele[12][15];
    ele[12][10] != ele[12][16];
    ele[12][10] != ele[12][17];
    ele[12][10] != ele[12][18];
    ele[12][10] != ele[12][19];
    ele[12][10] != ele[12][20];
    ele[12][10] != ele[12][21];
    ele[12][10] != ele[12][22];
    ele[12][10] != ele[12][23];
    ele[12][10] != ele[12][24];
    ele[12][10] != ele[12][25];
    ele[12][10] != ele[12][26];
    ele[12][10] != ele[12][27];
    ele[12][10] != ele[12][28];
    ele[12][10] != ele[12][29];
    ele[12][10] != ele[12][30];
    ele[12][10] != ele[12][31];
    ele[12][10] != ele[12][32];
    ele[12][10] != ele[12][33];
    ele[12][10] != ele[12][34];
    ele[12][10] != ele[12][35];
    ele[12][10] != ele[13][10];
    ele[12][10] != ele[13][11];
    ele[12][10] != ele[13][6];
    ele[12][10] != ele[13][7];
    ele[12][10] != ele[13][8];
    ele[12][10] != ele[13][9];
    ele[12][10] != ele[14][10];
    ele[12][10] != ele[14][11];
    ele[12][10] != ele[14][6];
    ele[12][10] != ele[14][7];
    ele[12][10] != ele[14][8];
    ele[12][10] != ele[14][9];
    ele[12][10] != ele[15][10];
    ele[12][10] != ele[15][11];
    ele[12][10] != ele[15][6];
    ele[12][10] != ele[15][7];
    ele[12][10] != ele[15][8];
    ele[12][10] != ele[15][9];
    ele[12][10] != ele[16][10];
    ele[12][10] != ele[16][11];
    ele[12][10] != ele[16][6];
    ele[12][10] != ele[16][7];
    ele[12][10] != ele[16][8];
    ele[12][10] != ele[16][9];
    ele[12][10] != ele[17][10];
    ele[12][10] != ele[17][11];
    ele[12][10] != ele[17][6];
    ele[12][10] != ele[17][7];
    ele[12][10] != ele[17][8];
    ele[12][10] != ele[17][9];
    ele[12][10] != ele[18][10];
    ele[12][10] != ele[19][10];
    ele[12][10] != ele[20][10];
    ele[12][10] != ele[21][10];
    ele[12][10] != ele[22][10];
    ele[12][10] != ele[23][10];
    ele[12][10] != ele[24][10];
    ele[12][10] != ele[25][10];
    ele[12][10] != ele[26][10];
    ele[12][10] != ele[27][10];
    ele[12][10] != ele[28][10];
    ele[12][10] != ele[29][10];
    ele[12][10] != ele[30][10];
    ele[12][10] != ele[31][10];
    ele[12][10] != ele[32][10];
    ele[12][10] != ele[33][10];
    ele[12][10] != ele[34][10];
    ele[12][10] != ele[35][10];
    ele[12][11] != ele[12][12];
    ele[12][11] != ele[12][13];
    ele[12][11] != ele[12][14];
    ele[12][11] != ele[12][15];
    ele[12][11] != ele[12][16];
    ele[12][11] != ele[12][17];
    ele[12][11] != ele[12][18];
    ele[12][11] != ele[12][19];
    ele[12][11] != ele[12][20];
    ele[12][11] != ele[12][21];
    ele[12][11] != ele[12][22];
    ele[12][11] != ele[12][23];
    ele[12][11] != ele[12][24];
    ele[12][11] != ele[12][25];
    ele[12][11] != ele[12][26];
    ele[12][11] != ele[12][27];
    ele[12][11] != ele[12][28];
    ele[12][11] != ele[12][29];
    ele[12][11] != ele[12][30];
    ele[12][11] != ele[12][31];
    ele[12][11] != ele[12][32];
    ele[12][11] != ele[12][33];
    ele[12][11] != ele[12][34];
    ele[12][11] != ele[12][35];
    ele[12][11] != ele[13][10];
    ele[12][11] != ele[13][11];
    ele[12][11] != ele[13][6];
    ele[12][11] != ele[13][7];
    ele[12][11] != ele[13][8];
    ele[12][11] != ele[13][9];
    ele[12][11] != ele[14][10];
    ele[12][11] != ele[14][11];
    ele[12][11] != ele[14][6];
    ele[12][11] != ele[14][7];
    ele[12][11] != ele[14][8];
    ele[12][11] != ele[14][9];
    ele[12][11] != ele[15][10];
    ele[12][11] != ele[15][11];
    ele[12][11] != ele[15][6];
    ele[12][11] != ele[15][7];
    ele[12][11] != ele[15][8];
    ele[12][11] != ele[15][9];
    ele[12][11] != ele[16][10];
    ele[12][11] != ele[16][11];
    ele[12][11] != ele[16][6];
    ele[12][11] != ele[16][7];
    ele[12][11] != ele[16][8];
    ele[12][11] != ele[16][9];
    ele[12][11] != ele[17][10];
    ele[12][11] != ele[17][11];
    ele[12][11] != ele[17][6];
    ele[12][11] != ele[17][7];
    ele[12][11] != ele[17][8];
    ele[12][11] != ele[17][9];
    ele[12][11] != ele[18][11];
    ele[12][11] != ele[19][11];
    ele[12][11] != ele[20][11];
    ele[12][11] != ele[21][11];
    ele[12][11] != ele[22][11];
    ele[12][11] != ele[23][11];
    ele[12][11] != ele[24][11];
    ele[12][11] != ele[25][11];
    ele[12][11] != ele[26][11];
    ele[12][11] != ele[27][11];
    ele[12][11] != ele[28][11];
    ele[12][11] != ele[29][11];
    ele[12][11] != ele[30][11];
    ele[12][11] != ele[31][11];
    ele[12][11] != ele[32][11];
    ele[12][11] != ele[33][11];
    ele[12][11] != ele[34][11];
    ele[12][11] != ele[35][11];
    ele[12][12] != ele[12][13];
    ele[12][12] != ele[12][14];
    ele[12][12] != ele[12][15];
    ele[12][12] != ele[12][16];
    ele[12][12] != ele[12][17];
    ele[12][12] != ele[12][18];
    ele[12][12] != ele[12][19];
    ele[12][12] != ele[12][20];
    ele[12][12] != ele[12][21];
    ele[12][12] != ele[12][22];
    ele[12][12] != ele[12][23];
    ele[12][12] != ele[12][24];
    ele[12][12] != ele[12][25];
    ele[12][12] != ele[12][26];
    ele[12][12] != ele[12][27];
    ele[12][12] != ele[12][28];
    ele[12][12] != ele[12][29];
    ele[12][12] != ele[12][30];
    ele[12][12] != ele[12][31];
    ele[12][12] != ele[12][32];
    ele[12][12] != ele[12][33];
    ele[12][12] != ele[12][34];
    ele[12][12] != ele[12][35];
    ele[12][12] != ele[13][12];
    ele[12][12] != ele[13][13];
    ele[12][12] != ele[13][14];
    ele[12][12] != ele[13][15];
    ele[12][12] != ele[13][16];
    ele[12][12] != ele[13][17];
    ele[12][12] != ele[14][12];
    ele[12][12] != ele[14][13];
    ele[12][12] != ele[14][14];
    ele[12][12] != ele[14][15];
    ele[12][12] != ele[14][16];
    ele[12][12] != ele[14][17];
    ele[12][12] != ele[15][12];
    ele[12][12] != ele[15][13];
    ele[12][12] != ele[15][14];
    ele[12][12] != ele[15][15];
    ele[12][12] != ele[15][16];
    ele[12][12] != ele[15][17];
    ele[12][12] != ele[16][12];
    ele[12][12] != ele[16][13];
    ele[12][12] != ele[16][14];
    ele[12][12] != ele[16][15];
    ele[12][12] != ele[16][16];
    ele[12][12] != ele[16][17];
    ele[12][12] != ele[17][12];
    ele[12][12] != ele[17][13];
    ele[12][12] != ele[17][14];
    ele[12][12] != ele[17][15];
    ele[12][12] != ele[17][16];
    ele[12][12] != ele[17][17];
    ele[12][12] != ele[18][12];
    ele[12][12] != ele[19][12];
    ele[12][12] != ele[20][12];
    ele[12][12] != ele[21][12];
    ele[12][12] != ele[22][12];
    ele[12][12] != ele[23][12];
    ele[12][12] != ele[24][12];
    ele[12][12] != ele[25][12];
    ele[12][12] != ele[26][12];
    ele[12][12] != ele[27][12];
    ele[12][12] != ele[28][12];
    ele[12][12] != ele[29][12];
    ele[12][12] != ele[30][12];
    ele[12][12] != ele[31][12];
    ele[12][12] != ele[32][12];
    ele[12][12] != ele[33][12];
    ele[12][12] != ele[34][12];
    ele[12][12] != ele[35][12];
    ele[12][13] != ele[12][14];
    ele[12][13] != ele[12][15];
    ele[12][13] != ele[12][16];
    ele[12][13] != ele[12][17];
    ele[12][13] != ele[12][18];
    ele[12][13] != ele[12][19];
    ele[12][13] != ele[12][20];
    ele[12][13] != ele[12][21];
    ele[12][13] != ele[12][22];
    ele[12][13] != ele[12][23];
    ele[12][13] != ele[12][24];
    ele[12][13] != ele[12][25];
    ele[12][13] != ele[12][26];
    ele[12][13] != ele[12][27];
    ele[12][13] != ele[12][28];
    ele[12][13] != ele[12][29];
    ele[12][13] != ele[12][30];
    ele[12][13] != ele[12][31];
    ele[12][13] != ele[12][32];
    ele[12][13] != ele[12][33];
    ele[12][13] != ele[12][34];
    ele[12][13] != ele[12][35];
    ele[12][13] != ele[13][12];
    ele[12][13] != ele[13][13];
    ele[12][13] != ele[13][14];
    ele[12][13] != ele[13][15];
    ele[12][13] != ele[13][16];
    ele[12][13] != ele[13][17];
    ele[12][13] != ele[14][12];
    ele[12][13] != ele[14][13];
    ele[12][13] != ele[14][14];
    ele[12][13] != ele[14][15];
    ele[12][13] != ele[14][16];
    ele[12][13] != ele[14][17];
    ele[12][13] != ele[15][12];
    ele[12][13] != ele[15][13];
    ele[12][13] != ele[15][14];
    ele[12][13] != ele[15][15];
    ele[12][13] != ele[15][16];
    ele[12][13] != ele[15][17];
    ele[12][13] != ele[16][12];
    ele[12][13] != ele[16][13];
    ele[12][13] != ele[16][14];
    ele[12][13] != ele[16][15];
    ele[12][13] != ele[16][16];
    ele[12][13] != ele[16][17];
    ele[12][13] != ele[17][12];
    ele[12][13] != ele[17][13];
    ele[12][13] != ele[17][14];
    ele[12][13] != ele[17][15];
    ele[12][13] != ele[17][16];
    ele[12][13] != ele[17][17];
    ele[12][13] != ele[18][13];
    ele[12][13] != ele[19][13];
    ele[12][13] != ele[20][13];
    ele[12][13] != ele[21][13];
    ele[12][13] != ele[22][13];
    ele[12][13] != ele[23][13];
    ele[12][13] != ele[24][13];
    ele[12][13] != ele[25][13];
    ele[12][13] != ele[26][13];
    ele[12][13] != ele[27][13];
    ele[12][13] != ele[28][13];
    ele[12][13] != ele[29][13];
    ele[12][13] != ele[30][13];
    ele[12][13] != ele[31][13];
    ele[12][13] != ele[32][13];
    ele[12][13] != ele[33][13];
    ele[12][13] != ele[34][13];
    ele[12][13] != ele[35][13];
    ele[12][14] != ele[12][15];
    ele[12][14] != ele[12][16];
    ele[12][14] != ele[12][17];
    ele[12][14] != ele[12][18];
    ele[12][14] != ele[12][19];
    ele[12][14] != ele[12][20];
    ele[12][14] != ele[12][21];
    ele[12][14] != ele[12][22];
    ele[12][14] != ele[12][23];
    ele[12][14] != ele[12][24];
    ele[12][14] != ele[12][25];
    ele[12][14] != ele[12][26];
    ele[12][14] != ele[12][27];
    ele[12][14] != ele[12][28];
    ele[12][14] != ele[12][29];
    ele[12][14] != ele[12][30];
    ele[12][14] != ele[12][31];
    ele[12][14] != ele[12][32];
    ele[12][14] != ele[12][33];
    ele[12][14] != ele[12][34];
    ele[12][14] != ele[12][35];
    ele[12][14] != ele[13][12];
    ele[12][14] != ele[13][13];
    ele[12][14] != ele[13][14];
    ele[12][14] != ele[13][15];
    ele[12][14] != ele[13][16];
    ele[12][14] != ele[13][17];
    ele[12][14] != ele[14][12];
    ele[12][14] != ele[14][13];
    ele[12][14] != ele[14][14];
    ele[12][14] != ele[14][15];
    ele[12][14] != ele[14][16];
    ele[12][14] != ele[14][17];
    ele[12][14] != ele[15][12];
    ele[12][14] != ele[15][13];
    ele[12][14] != ele[15][14];
    ele[12][14] != ele[15][15];
    ele[12][14] != ele[15][16];
    ele[12][14] != ele[15][17];
    ele[12][14] != ele[16][12];
    ele[12][14] != ele[16][13];
    ele[12][14] != ele[16][14];
    ele[12][14] != ele[16][15];
    ele[12][14] != ele[16][16];
    ele[12][14] != ele[16][17];
    ele[12][14] != ele[17][12];
    ele[12][14] != ele[17][13];
    ele[12][14] != ele[17][14];
    ele[12][14] != ele[17][15];
    ele[12][14] != ele[17][16];
    ele[12][14] != ele[17][17];
    ele[12][14] != ele[18][14];
    ele[12][14] != ele[19][14];
    ele[12][14] != ele[20][14];
    ele[12][14] != ele[21][14];
    ele[12][14] != ele[22][14];
    ele[12][14] != ele[23][14];
    ele[12][14] != ele[24][14];
    ele[12][14] != ele[25][14];
    ele[12][14] != ele[26][14];
    ele[12][14] != ele[27][14];
    ele[12][14] != ele[28][14];
    ele[12][14] != ele[29][14];
    ele[12][14] != ele[30][14];
    ele[12][14] != ele[31][14];
    ele[12][14] != ele[32][14];
    ele[12][14] != ele[33][14];
    ele[12][14] != ele[34][14];
    ele[12][14] != ele[35][14];
    ele[12][15] != ele[12][16];
    ele[12][15] != ele[12][17];
    ele[12][15] != ele[12][18];
    ele[12][15] != ele[12][19];
    ele[12][15] != ele[12][20];
    ele[12][15] != ele[12][21];
    ele[12][15] != ele[12][22];
    ele[12][15] != ele[12][23];
    ele[12][15] != ele[12][24];
    ele[12][15] != ele[12][25];
    ele[12][15] != ele[12][26];
    ele[12][15] != ele[12][27];
    ele[12][15] != ele[12][28];
    ele[12][15] != ele[12][29];
    ele[12][15] != ele[12][30];
    ele[12][15] != ele[12][31];
    ele[12][15] != ele[12][32];
    ele[12][15] != ele[12][33];
    ele[12][15] != ele[12][34];
    ele[12][15] != ele[12][35];
    ele[12][15] != ele[13][12];
    ele[12][15] != ele[13][13];
    ele[12][15] != ele[13][14];
    ele[12][15] != ele[13][15];
    ele[12][15] != ele[13][16];
    ele[12][15] != ele[13][17];
    ele[12][15] != ele[14][12];
    ele[12][15] != ele[14][13];
    ele[12][15] != ele[14][14];
    ele[12][15] != ele[14][15];
    ele[12][15] != ele[14][16];
    ele[12][15] != ele[14][17];
    ele[12][15] != ele[15][12];
    ele[12][15] != ele[15][13];
    ele[12][15] != ele[15][14];
    ele[12][15] != ele[15][15];
    ele[12][15] != ele[15][16];
    ele[12][15] != ele[15][17];
    ele[12][15] != ele[16][12];
    ele[12][15] != ele[16][13];
    ele[12][15] != ele[16][14];
    ele[12][15] != ele[16][15];
    ele[12][15] != ele[16][16];
    ele[12][15] != ele[16][17];
    ele[12][15] != ele[17][12];
    ele[12][15] != ele[17][13];
    ele[12][15] != ele[17][14];
    ele[12][15] != ele[17][15];
    ele[12][15] != ele[17][16];
    ele[12][15] != ele[17][17];
    ele[12][15] != ele[18][15];
    ele[12][15] != ele[19][15];
    ele[12][15] != ele[20][15];
    ele[12][15] != ele[21][15];
    ele[12][15] != ele[22][15];
    ele[12][15] != ele[23][15];
    ele[12][15] != ele[24][15];
    ele[12][15] != ele[25][15];
    ele[12][15] != ele[26][15];
    ele[12][15] != ele[27][15];
    ele[12][15] != ele[28][15];
    ele[12][15] != ele[29][15];
    ele[12][15] != ele[30][15];
    ele[12][15] != ele[31][15];
    ele[12][15] != ele[32][15];
    ele[12][15] != ele[33][15];
    ele[12][15] != ele[34][15];
    ele[12][15] != ele[35][15];
    ele[12][16] != ele[12][17];
    ele[12][16] != ele[12][18];
    ele[12][16] != ele[12][19];
    ele[12][16] != ele[12][20];
    ele[12][16] != ele[12][21];
    ele[12][16] != ele[12][22];
    ele[12][16] != ele[12][23];
    ele[12][16] != ele[12][24];
    ele[12][16] != ele[12][25];
    ele[12][16] != ele[12][26];
    ele[12][16] != ele[12][27];
    ele[12][16] != ele[12][28];
    ele[12][16] != ele[12][29];
    ele[12][16] != ele[12][30];
    ele[12][16] != ele[12][31];
    ele[12][16] != ele[12][32];
    ele[12][16] != ele[12][33];
    ele[12][16] != ele[12][34];
    ele[12][16] != ele[12][35];
    ele[12][16] != ele[13][12];
    ele[12][16] != ele[13][13];
    ele[12][16] != ele[13][14];
    ele[12][16] != ele[13][15];
    ele[12][16] != ele[13][16];
    ele[12][16] != ele[13][17];
    ele[12][16] != ele[14][12];
    ele[12][16] != ele[14][13];
    ele[12][16] != ele[14][14];
    ele[12][16] != ele[14][15];
    ele[12][16] != ele[14][16];
    ele[12][16] != ele[14][17];
    ele[12][16] != ele[15][12];
    ele[12][16] != ele[15][13];
    ele[12][16] != ele[15][14];
    ele[12][16] != ele[15][15];
    ele[12][16] != ele[15][16];
    ele[12][16] != ele[15][17];
    ele[12][16] != ele[16][12];
    ele[12][16] != ele[16][13];
    ele[12][16] != ele[16][14];
    ele[12][16] != ele[16][15];
    ele[12][16] != ele[16][16];
    ele[12][16] != ele[16][17];
    ele[12][16] != ele[17][12];
    ele[12][16] != ele[17][13];
    ele[12][16] != ele[17][14];
    ele[12][16] != ele[17][15];
    ele[12][16] != ele[17][16];
    ele[12][16] != ele[17][17];
    ele[12][16] != ele[18][16];
    ele[12][16] != ele[19][16];
    ele[12][16] != ele[20][16];
    ele[12][16] != ele[21][16];
    ele[12][16] != ele[22][16];
    ele[12][16] != ele[23][16];
    ele[12][16] != ele[24][16];
    ele[12][16] != ele[25][16];
    ele[12][16] != ele[26][16];
    ele[12][16] != ele[27][16];
    ele[12][16] != ele[28][16];
    ele[12][16] != ele[29][16];
    ele[12][16] != ele[30][16];
    ele[12][16] != ele[31][16];
    ele[12][16] != ele[32][16];
    ele[12][16] != ele[33][16];
    ele[12][16] != ele[34][16];
    ele[12][16] != ele[35][16];
    ele[12][17] != ele[12][18];
    ele[12][17] != ele[12][19];
    ele[12][17] != ele[12][20];
    ele[12][17] != ele[12][21];
    ele[12][17] != ele[12][22];
    ele[12][17] != ele[12][23];
    ele[12][17] != ele[12][24];
    ele[12][17] != ele[12][25];
    ele[12][17] != ele[12][26];
    ele[12][17] != ele[12][27];
    ele[12][17] != ele[12][28];
    ele[12][17] != ele[12][29];
    ele[12][17] != ele[12][30];
    ele[12][17] != ele[12][31];
    ele[12][17] != ele[12][32];
    ele[12][17] != ele[12][33];
    ele[12][17] != ele[12][34];
    ele[12][17] != ele[12][35];
    ele[12][17] != ele[13][12];
    ele[12][17] != ele[13][13];
    ele[12][17] != ele[13][14];
    ele[12][17] != ele[13][15];
    ele[12][17] != ele[13][16];
    ele[12][17] != ele[13][17];
    ele[12][17] != ele[14][12];
    ele[12][17] != ele[14][13];
    ele[12][17] != ele[14][14];
    ele[12][17] != ele[14][15];
    ele[12][17] != ele[14][16];
    ele[12][17] != ele[14][17];
    ele[12][17] != ele[15][12];
    ele[12][17] != ele[15][13];
    ele[12][17] != ele[15][14];
    ele[12][17] != ele[15][15];
    ele[12][17] != ele[15][16];
    ele[12][17] != ele[15][17];
    ele[12][17] != ele[16][12];
    ele[12][17] != ele[16][13];
    ele[12][17] != ele[16][14];
    ele[12][17] != ele[16][15];
    ele[12][17] != ele[16][16];
    ele[12][17] != ele[16][17];
    ele[12][17] != ele[17][12];
    ele[12][17] != ele[17][13];
    ele[12][17] != ele[17][14];
    ele[12][17] != ele[17][15];
    ele[12][17] != ele[17][16];
    ele[12][17] != ele[17][17];
    ele[12][17] != ele[18][17];
    ele[12][17] != ele[19][17];
    ele[12][17] != ele[20][17];
    ele[12][17] != ele[21][17];
    ele[12][17] != ele[22][17];
    ele[12][17] != ele[23][17];
    ele[12][17] != ele[24][17];
    ele[12][17] != ele[25][17];
    ele[12][17] != ele[26][17];
    ele[12][17] != ele[27][17];
    ele[12][17] != ele[28][17];
    ele[12][17] != ele[29][17];
    ele[12][17] != ele[30][17];
    ele[12][17] != ele[31][17];
    ele[12][17] != ele[32][17];
    ele[12][17] != ele[33][17];
    ele[12][17] != ele[34][17];
    ele[12][17] != ele[35][17];
    ele[12][18] != ele[12][19];
    ele[12][18] != ele[12][20];
    ele[12][18] != ele[12][21];
    ele[12][18] != ele[12][22];
    ele[12][18] != ele[12][23];
    ele[12][18] != ele[12][24];
    ele[12][18] != ele[12][25];
    ele[12][18] != ele[12][26];
    ele[12][18] != ele[12][27];
    ele[12][18] != ele[12][28];
    ele[12][18] != ele[12][29];
    ele[12][18] != ele[12][30];
    ele[12][18] != ele[12][31];
    ele[12][18] != ele[12][32];
    ele[12][18] != ele[12][33];
    ele[12][18] != ele[12][34];
    ele[12][18] != ele[12][35];
    ele[12][18] != ele[13][18];
    ele[12][18] != ele[13][19];
    ele[12][18] != ele[13][20];
    ele[12][18] != ele[13][21];
    ele[12][18] != ele[13][22];
    ele[12][18] != ele[13][23];
    ele[12][18] != ele[14][18];
    ele[12][18] != ele[14][19];
    ele[12][18] != ele[14][20];
    ele[12][18] != ele[14][21];
    ele[12][18] != ele[14][22];
    ele[12][18] != ele[14][23];
    ele[12][18] != ele[15][18];
    ele[12][18] != ele[15][19];
    ele[12][18] != ele[15][20];
    ele[12][18] != ele[15][21];
    ele[12][18] != ele[15][22];
    ele[12][18] != ele[15][23];
    ele[12][18] != ele[16][18];
    ele[12][18] != ele[16][19];
    ele[12][18] != ele[16][20];
    ele[12][18] != ele[16][21];
    ele[12][18] != ele[16][22];
    ele[12][18] != ele[16][23];
    ele[12][18] != ele[17][18];
    ele[12][18] != ele[17][19];
    ele[12][18] != ele[17][20];
    ele[12][18] != ele[17][21];
    ele[12][18] != ele[17][22];
    ele[12][18] != ele[17][23];
    ele[12][18] != ele[18][18];
    ele[12][18] != ele[19][18];
    ele[12][18] != ele[20][18];
    ele[12][18] != ele[21][18];
    ele[12][18] != ele[22][18];
    ele[12][18] != ele[23][18];
    ele[12][18] != ele[24][18];
    ele[12][18] != ele[25][18];
    ele[12][18] != ele[26][18];
    ele[12][18] != ele[27][18];
    ele[12][18] != ele[28][18];
    ele[12][18] != ele[29][18];
    ele[12][18] != ele[30][18];
    ele[12][18] != ele[31][18];
    ele[12][18] != ele[32][18];
    ele[12][18] != ele[33][18];
    ele[12][18] != ele[34][18];
    ele[12][18] != ele[35][18];
    ele[12][19] != ele[12][20];
    ele[12][19] != ele[12][21];
    ele[12][19] != ele[12][22];
    ele[12][19] != ele[12][23];
    ele[12][19] != ele[12][24];
    ele[12][19] != ele[12][25];
    ele[12][19] != ele[12][26];
    ele[12][19] != ele[12][27];
    ele[12][19] != ele[12][28];
    ele[12][19] != ele[12][29];
    ele[12][19] != ele[12][30];
    ele[12][19] != ele[12][31];
    ele[12][19] != ele[12][32];
    ele[12][19] != ele[12][33];
    ele[12][19] != ele[12][34];
    ele[12][19] != ele[12][35];
    ele[12][19] != ele[13][18];
    ele[12][19] != ele[13][19];
    ele[12][19] != ele[13][20];
    ele[12][19] != ele[13][21];
    ele[12][19] != ele[13][22];
    ele[12][19] != ele[13][23];
    ele[12][19] != ele[14][18];
    ele[12][19] != ele[14][19];
    ele[12][19] != ele[14][20];
    ele[12][19] != ele[14][21];
    ele[12][19] != ele[14][22];
    ele[12][19] != ele[14][23];
    ele[12][19] != ele[15][18];
    ele[12][19] != ele[15][19];
    ele[12][19] != ele[15][20];
    ele[12][19] != ele[15][21];
    ele[12][19] != ele[15][22];
    ele[12][19] != ele[15][23];
    ele[12][19] != ele[16][18];
    ele[12][19] != ele[16][19];
    ele[12][19] != ele[16][20];
    ele[12][19] != ele[16][21];
    ele[12][19] != ele[16][22];
    ele[12][19] != ele[16][23];
    ele[12][19] != ele[17][18];
    ele[12][19] != ele[17][19];
    ele[12][19] != ele[17][20];
    ele[12][19] != ele[17][21];
    ele[12][19] != ele[17][22];
    ele[12][19] != ele[17][23];
    ele[12][19] != ele[18][19];
    ele[12][19] != ele[19][19];
    ele[12][19] != ele[20][19];
    ele[12][19] != ele[21][19];
    ele[12][19] != ele[22][19];
    ele[12][19] != ele[23][19];
    ele[12][19] != ele[24][19];
    ele[12][19] != ele[25][19];
    ele[12][19] != ele[26][19];
    ele[12][19] != ele[27][19];
    ele[12][19] != ele[28][19];
    ele[12][19] != ele[29][19];
    ele[12][19] != ele[30][19];
    ele[12][19] != ele[31][19];
    ele[12][19] != ele[32][19];
    ele[12][19] != ele[33][19];
    ele[12][19] != ele[34][19];
    ele[12][19] != ele[35][19];
    ele[12][2] != ele[12][10];
    ele[12][2] != ele[12][11];
    ele[12][2] != ele[12][12];
    ele[12][2] != ele[12][13];
    ele[12][2] != ele[12][14];
    ele[12][2] != ele[12][15];
    ele[12][2] != ele[12][16];
    ele[12][2] != ele[12][17];
    ele[12][2] != ele[12][18];
    ele[12][2] != ele[12][19];
    ele[12][2] != ele[12][20];
    ele[12][2] != ele[12][21];
    ele[12][2] != ele[12][22];
    ele[12][2] != ele[12][23];
    ele[12][2] != ele[12][24];
    ele[12][2] != ele[12][25];
    ele[12][2] != ele[12][26];
    ele[12][2] != ele[12][27];
    ele[12][2] != ele[12][28];
    ele[12][2] != ele[12][29];
    ele[12][2] != ele[12][3];
    ele[12][2] != ele[12][30];
    ele[12][2] != ele[12][31];
    ele[12][2] != ele[12][32];
    ele[12][2] != ele[12][33];
    ele[12][2] != ele[12][34];
    ele[12][2] != ele[12][35];
    ele[12][2] != ele[12][4];
    ele[12][2] != ele[12][5];
    ele[12][2] != ele[12][6];
    ele[12][2] != ele[12][7];
    ele[12][2] != ele[12][8];
    ele[12][2] != ele[12][9];
    ele[12][2] != ele[13][0];
    ele[12][2] != ele[13][1];
    ele[12][2] != ele[13][2];
    ele[12][2] != ele[13][3];
    ele[12][2] != ele[13][4];
    ele[12][2] != ele[13][5];
    ele[12][2] != ele[14][0];
    ele[12][2] != ele[14][1];
    ele[12][2] != ele[14][2];
    ele[12][2] != ele[14][3];
    ele[12][2] != ele[14][4];
    ele[12][2] != ele[14][5];
    ele[12][2] != ele[15][0];
    ele[12][2] != ele[15][1];
    ele[12][2] != ele[15][2];
    ele[12][2] != ele[15][3];
    ele[12][2] != ele[15][4];
    ele[12][2] != ele[15][5];
    ele[12][2] != ele[16][0];
    ele[12][2] != ele[16][1];
    ele[12][2] != ele[16][2];
    ele[12][2] != ele[16][3];
    ele[12][2] != ele[16][4];
    ele[12][2] != ele[16][5];
    ele[12][2] != ele[17][0];
    ele[12][2] != ele[17][1];
    ele[12][2] != ele[17][2];
    ele[12][2] != ele[17][3];
    ele[12][2] != ele[17][4];
    ele[12][2] != ele[17][5];
    ele[12][2] != ele[18][2];
    ele[12][2] != ele[19][2];
    ele[12][2] != ele[20][2];
    ele[12][2] != ele[21][2];
    ele[12][2] != ele[22][2];
    ele[12][2] != ele[23][2];
    ele[12][2] != ele[24][2];
    ele[12][2] != ele[25][2];
    ele[12][2] != ele[26][2];
    ele[12][2] != ele[27][2];
    ele[12][2] != ele[28][2];
    ele[12][2] != ele[29][2];
    ele[12][2] != ele[30][2];
    ele[12][2] != ele[31][2];
    ele[12][2] != ele[32][2];
    ele[12][2] != ele[33][2];
    ele[12][2] != ele[34][2];
    ele[12][2] != ele[35][2];
    ele[12][20] != ele[12][21];
    ele[12][20] != ele[12][22];
    ele[12][20] != ele[12][23];
    ele[12][20] != ele[12][24];
    ele[12][20] != ele[12][25];
    ele[12][20] != ele[12][26];
    ele[12][20] != ele[12][27];
    ele[12][20] != ele[12][28];
    ele[12][20] != ele[12][29];
    ele[12][20] != ele[12][30];
    ele[12][20] != ele[12][31];
    ele[12][20] != ele[12][32];
    ele[12][20] != ele[12][33];
    ele[12][20] != ele[12][34];
    ele[12][20] != ele[12][35];
    ele[12][20] != ele[13][18];
    ele[12][20] != ele[13][19];
    ele[12][20] != ele[13][20];
    ele[12][20] != ele[13][21];
    ele[12][20] != ele[13][22];
    ele[12][20] != ele[13][23];
    ele[12][20] != ele[14][18];
    ele[12][20] != ele[14][19];
    ele[12][20] != ele[14][20];
    ele[12][20] != ele[14][21];
    ele[12][20] != ele[14][22];
    ele[12][20] != ele[14][23];
    ele[12][20] != ele[15][18];
    ele[12][20] != ele[15][19];
    ele[12][20] != ele[15][20];
    ele[12][20] != ele[15][21];
    ele[12][20] != ele[15][22];
    ele[12][20] != ele[15][23];
    ele[12][20] != ele[16][18];
    ele[12][20] != ele[16][19];
    ele[12][20] != ele[16][20];
    ele[12][20] != ele[16][21];
    ele[12][20] != ele[16][22];
    ele[12][20] != ele[16][23];
    ele[12][20] != ele[17][18];
    ele[12][20] != ele[17][19];
    ele[12][20] != ele[17][20];
    ele[12][20] != ele[17][21];
    ele[12][20] != ele[17][22];
    ele[12][20] != ele[17][23];
    ele[12][20] != ele[18][20];
    ele[12][20] != ele[19][20];
    ele[12][20] != ele[20][20];
    ele[12][20] != ele[21][20];
    ele[12][20] != ele[22][20];
    ele[12][20] != ele[23][20];
    ele[12][20] != ele[24][20];
    ele[12][20] != ele[25][20];
    ele[12][20] != ele[26][20];
    ele[12][20] != ele[27][20];
    ele[12][20] != ele[28][20];
    ele[12][20] != ele[29][20];
    ele[12][20] != ele[30][20];
    ele[12][20] != ele[31][20];
    ele[12][20] != ele[32][20];
    ele[12][20] != ele[33][20];
    ele[12][20] != ele[34][20];
    ele[12][20] != ele[35][20];
    ele[12][21] != ele[12][22];
    ele[12][21] != ele[12][23];
    ele[12][21] != ele[12][24];
    ele[12][21] != ele[12][25];
    ele[12][21] != ele[12][26];
    ele[12][21] != ele[12][27];
    ele[12][21] != ele[12][28];
    ele[12][21] != ele[12][29];
    ele[12][21] != ele[12][30];
    ele[12][21] != ele[12][31];
    ele[12][21] != ele[12][32];
    ele[12][21] != ele[12][33];
    ele[12][21] != ele[12][34];
    ele[12][21] != ele[12][35];
    ele[12][21] != ele[13][18];
    ele[12][21] != ele[13][19];
    ele[12][21] != ele[13][20];
    ele[12][21] != ele[13][21];
    ele[12][21] != ele[13][22];
    ele[12][21] != ele[13][23];
    ele[12][21] != ele[14][18];
    ele[12][21] != ele[14][19];
    ele[12][21] != ele[14][20];
    ele[12][21] != ele[14][21];
    ele[12][21] != ele[14][22];
    ele[12][21] != ele[14][23];
    ele[12][21] != ele[15][18];
    ele[12][21] != ele[15][19];
    ele[12][21] != ele[15][20];
    ele[12][21] != ele[15][21];
    ele[12][21] != ele[15][22];
    ele[12][21] != ele[15][23];
    ele[12][21] != ele[16][18];
    ele[12][21] != ele[16][19];
    ele[12][21] != ele[16][20];
    ele[12][21] != ele[16][21];
    ele[12][21] != ele[16][22];
    ele[12][21] != ele[16][23];
    ele[12][21] != ele[17][18];
    ele[12][21] != ele[17][19];
    ele[12][21] != ele[17][20];
    ele[12][21] != ele[17][21];
    ele[12][21] != ele[17][22];
    ele[12][21] != ele[17][23];
    ele[12][21] != ele[18][21];
    ele[12][21] != ele[19][21];
    ele[12][21] != ele[20][21];
    ele[12][21] != ele[21][21];
    ele[12][21] != ele[22][21];
    ele[12][21] != ele[23][21];
    ele[12][21] != ele[24][21];
    ele[12][21] != ele[25][21];
    ele[12][21] != ele[26][21];
    ele[12][21] != ele[27][21];
    ele[12][21] != ele[28][21];
    ele[12][21] != ele[29][21];
    ele[12][21] != ele[30][21];
    ele[12][21] != ele[31][21];
    ele[12][21] != ele[32][21];
    ele[12][21] != ele[33][21];
    ele[12][21] != ele[34][21];
    ele[12][21] != ele[35][21];
    ele[12][22] != ele[12][23];
    ele[12][22] != ele[12][24];
    ele[12][22] != ele[12][25];
    ele[12][22] != ele[12][26];
    ele[12][22] != ele[12][27];
    ele[12][22] != ele[12][28];
    ele[12][22] != ele[12][29];
    ele[12][22] != ele[12][30];
    ele[12][22] != ele[12][31];
    ele[12][22] != ele[12][32];
    ele[12][22] != ele[12][33];
    ele[12][22] != ele[12][34];
    ele[12][22] != ele[12][35];
    ele[12][22] != ele[13][18];
    ele[12][22] != ele[13][19];
    ele[12][22] != ele[13][20];
    ele[12][22] != ele[13][21];
    ele[12][22] != ele[13][22];
    ele[12][22] != ele[13][23];
    ele[12][22] != ele[14][18];
    ele[12][22] != ele[14][19];
    ele[12][22] != ele[14][20];
    ele[12][22] != ele[14][21];
    ele[12][22] != ele[14][22];
    ele[12][22] != ele[14][23];
    ele[12][22] != ele[15][18];
    ele[12][22] != ele[15][19];
    ele[12][22] != ele[15][20];
    ele[12][22] != ele[15][21];
    ele[12][22] != ele[15][22];
    ele[12][22] != ele[15][23];
    ele[12][22] != ele[16][18];
    ele[12][22] != ele[16][19];
    ele[12][22] != ele[16][20];
    ele[12][22] != ele[16][21];
    ele[12][22] != ele[16][22];
    ele[12][22] != ele[16][23];
    ele[12][22] != ele[17][18];
    ele[12][22] != ele[17][19];
    ele[12][22] != ele[17][20];
    ele[12][22] != ele[17][21];
    ele[12][22] != ele[17][22];
    ele[12][22] != ele[17][23];
    ele[12][22] != ele[18][22];
    ele[12][22] != ele[19][22];
    ele[12][22] != ele[20][22];
    ele[12][22] != ele[21][22];
    ele[12][22] != ele[22][22];
    ele[12][22] != ele[23][22];
    ele[12][22] != ele[24][22];
    ele[12][22] != ele[25][22];
    ele[12][22] != ele[26][22];
    ele[12][22] != ele[27][22];
    ele[12][22] != ele[28][22];
    ele[12][22] != ele[29][22];
    ele[12][22] != ele[30][22];
    ele[12][22] != ele[31][22];
    ele[12][22] != ele[32][22];
    ele[12][22] != ele[33][22];
    ele[12][22] != ele[34][22];
    ele[12][22] != ele[35][22];
    ele[12][23] != ele[12][24];
    ele[12][23] != ele[12][25];
    ele[12][23] != ele[12][26];
    ele[12][23] != ele[12][27];
    ele[12][23] != ele[12][28];
    ele[12][23] != ele[12][29];
    ele[12][23] != ele[12][30];
    ele[12][23] != ele[12][31];
    ele[12][23] != ele[12][32];
    ele[12][23] != ele[12][33];
    ele[12][23] != ele[12][34];
    ele[12][23] != ele[12][35];
    ele[12][23] != ele[13][18];
    ele[12][23] != ele[13][19];
    ele[12][23] != ele[13][20];
    ele[12][23] != ele[13][21];
    ele[12][23] != ele[13][22];
    ele[12][23] != ele[13][23];
    ele[12][23] != ele[14][18];
    ele[12][23] != ele[14][19];
    ele[12][23] != ele[14][20];
    ele[12][23] != ele[14][21];
    ele[12][23] != ele[14][22];
    ele[12][23] != ele[14][23];
    ele[12][23] != ele[15][18];
    ele[12][23] != ele[15][19];
    ele[12][23] != ele[15][20];
    ele[12][23] != ele[15][21];
    ele[12][23] != ele[15][22];
    ele[12][23] != ele[15][23];
    ele[12][23] != ele[16][18];
    ele[12][23] != ele[16][19];
    ele[12][23] != ele[16][20];
    ele[12][23] != ele[16][21];
    ele[12][23] != ele[16][22];
    ele[12][23] != ele[16][23];
    ele[12][23] != ele[17][18];
    ele[12][23] != ele[17][19];
    ele[12][23] != ele[17][20];
    ele[12][23] != ele[17][21];
    ele[12][23] != ele[17][22];
    ele[12][23] != ele[17][23];
    ele[12][23] != ele[18][23];
    ele[12][23] != ele[19][23];
    ele[12][23] != ele[20][23];
    ele[12][23] != ele[21][23];
    ele[12][23] != ele[22][23];
    ele[12][23] != ele[23][23];
    ele[12][23] != ele[24][23];
    ele[12][23] != ele[25][23];
    ele[12][23] != ele[26][23];
    ele[12][23] != ele[27][23];
    ele[12][23] != ele[28][23];
    ele[12][23] != ele[29][23];
    ele[12][23] != ele[30][23];
    ele[12][23] != ele[31][23];
    ele[12][23] != ele[32][23];
    ele[12][23] != ele[33][23];
    ele[12][23] != ele[34][23];
    ele[12][23] != ele[35][23];
    ele[12][24] != ele[12][25];
    ele[12][24] != ele[12][26];
    ele[12][24] != ele[12][27];
    ele[12][24] != ele[12][28];
    ele[12][24] != ele[12][29];
    ele[12][24] != ele[12][30];
    ele[12][24] != ele[12][31];
    ele[12][24] != ele[12][32];
    ele[12][24] != ele[12][33];
    ele[12][24] != ele[12][34];
    ele[12][24] != ele[12][35];
    ele[12][24] != ele[13][24];
    ele[12][24] != ele[13][25];
    ele[12][24] != ele[13][26];
    ele[12][24] != ele[13][27];
    ele[12][24] != ele[13][28];
    ele[12][24] != ele[13][29];
    ele[12][24] != ele[14][24];
    ele[12][24] != ele[14][25];
    ele[12][24] != ele[14][26];
    ele[12][24] != ele[14][27];
    ele[12][24] != ele[14][28];
    ele[12][24] != ele[14][29];
    ele[12][24] != ele[15][24];
    ele[12][24] != ele[15][25];
    ele[12][24] != ele[15][26];
    ele[12][24] != ele[15][27];
    ele[12][24] != ele[15][28];
    ele[12][24] != ele[15][29];
    ele[12][24] != ele[16][24];
    ele[12][24] != ele[16][25];
    ele[12][24] != ele[16][26];
    ele[12][24] != ele[16][27];
    ele[12][24] != ele[16][28];
    ele[12][24] != ele[16][29];
    ele[12][24] != ele[17][24];
    ele[12][24] != ele[17][25];
    ele[12][24] != ele[17][26];
    ele[12][24] != ele[17][27];
    ele[12][24] != ele[17][28];
    ele[12][24] != ele[17][29];
    ele[12][24] != ele[18][24];
    ele[12][24] != ele[19][24];
    ele[12][24] != ele[20][24];
    ele[12][24] != ele[21][24];
    ele[12][24] != ele[22][24];
    ele[12][24] != ele[23][24];
    ele[12][24] != ele[24][24];
    ele[12][24] != ele[25][24];
    ele[12][24] != ele[26][24];
    ele[12][24] != ele[27][24];
    ele[12][24] != ele[28][24];
    ele[12][24] != ele[29][24];
    ele[12][24] != ele[30][24];
    ele[12][24] != ele[31][24];
    ele[12][24] != ele[32][24];
    ele[12][24] != ele[33][24];
    ele[12][24] != ele[34][24];
    ele[12][24] != ele[35][24];
    ele[12][25] != ele[12][26];
    ele[12][25] != ele[12][27];
    ele[12][25] != ele[12][28];
    ele[12][25] != ele[12][29];
    ele[12][25] != ele[12][30];
    ele[12][25] != ele[12][31];
    ele[12][25] != ele[12][32];
    ele[12][25] != ele[12][33];
    ele[12][25] != ele[12][34];
    ele[12][25] != ele[12][35];
    ele[12][25] != ele[13][24];
    ele[12][25] != ele[13][25];
    ele[12][25] != ele[13][26];
    ele[12][25] != ele[13][27];
    ele[12][25] != ele[13][28];
    ele[12][25] != ele[13][29];
    ele[12][25] != ele[14][24];
    ele[12][25] != ele[14][25];
    ele[12][25] != ele[14][26];
    ele[12][25] != ele[14][27];
    ele[12][25] != ele[14][28];
    ele[12][25] != ele[14][29];
    ele[12][25] != ele[15][24];
    ele[12][25] != ele[15][25];
    ele[12][25] != ele[15][26];
    ele[12][25] != ele[15][27];
    ele[12][25] != ele[15][28];
    ele[12][25] != ele[15][29];
    ele[12][25] != ele[16][24];
    ele[12][25] != ele[16][25];
    ele[12][25] != ele[16][26];
    ele[12][25] != ele[16][27];
    ele[12][25] != ele[16][28];
    ele[12][25] != ele[16][29];
    ele[12][25] != ele[17][24];
    ele[12][25] != ele[17][25];
    ele[12][25] != ele[17][26];
    ele[12][25] != ele[17][27];
    ele[12][25] != ele[17][28];
    ele[12][25] != ele[17][29];
    ele[12][25] != ele[18][25];
    ele[12][25] != ele[19][25];
    ele[12][25] != ele[20][25];
    ele[12][25] != ele[21][25];
    ele[12][25] != ele[22][25];
    ele[12][25] != ele[23][25];
    ele[12][25] != ele[24][25];
    ele[12][25] != ele[25][25];
    ele[12][25] != ele[26][25];
    ele[12][25] != ele[27][25];
    ele[12][25] != ele[28][25];
    ele[12][25] != ele[29][25];
    ele[12][25] != ele[30][25];
    ele[12][25] != ele[31][25];
    ele[12][25] != ele[32][25];
    ele[12][25] != ele[33][25];
    ele[12][25] != ele[34][25];
    ele[12][25] != ele[35][25];
    ele[12][26] != ele[12][27];
    ele[12][26] != ele[12][28];
    ele[12][26] != ele[12][29];
    ele[12][26] != ele[12][30];
    ele[12][26] != ele[12][31];
    ele[12][26] != ele[12][32];
    ele[12][26] != ele[12][33];
    ele[12][26] != ele[12][34];
    ele[12][26] != ele[12][35];
    ele[12][26] != ele[13][24];
    ele[12][26] != ele[13][25];
    ele[12][26] != ele[13][26];
    ele[12][26] != ele[13][27];
    ele[12][26] != ele[13][28];
    ele[12][26] != ele[13][29];
    ele[12][26] != ele[14][24];
    ele[12][26] != ele[14][25];
    ele[12][26] != ele[14][26];
    ele[12][26] != ele[14][27];
    ele[12][26] != ele[14][28];
    ele[12][26] != ele[14][29];
    ele[12][26] != ele[15][24];
    ele[12][26] != ele[15][25];
    ele[12][26] != ele[15][26];
    ele[12][26] != ele[15][27];
    ele[12][26] != ele[15][28];
    ele[12][26] != ele[15][29];
    ele[12][26] != ele[16][24];
    ele[12][26] != ele[16][25];
    ele[12][26] != ele[16][26];
    ele[12][26] != ele[16][27];
    ele[12][26] != ele[16][28];
    ele[12][26] != ele[16][29];
    ele[12][26] != ele[17][24];
    ele[12][26] != ele[17][25];
    ele[12][26] != ele[17][26];
    ele[12][26] != ele[17][27];
    ele[12][26] != ele[17][28];
    ele[12][26] != ele[17][29];
    ele[12][26] != ele[18][26];
    ele[12][26] != ele[19][26];
    ele[12][26] != ele[20][26];
    ele[12][26] != ele[21][26];
    ele[12][26] != ele[22][26];
    ele[12][26] != ele[23][26];
    ele[12][26] != ele[24][26];
    ele[12][26] != ele[25][26];
    ele[12][26] != ele[26][26];
    ele[12][26] != ele[27][26];
    ele[12][26] != ele[28][26];
    ele[12][26] != ele[29][26];
    ele[12][26] != ele[30][26];
    ele[12][26] != ele[31][26];
    ele[12][26] != ele[32][26];
    ele[12][26] != ele[33][26];
    ele[12][26] != ele[34][26];
    ele[12][26] != ele[35][26];
    ele[12][27] != ele[12][28];
    ele[12][27] != ele[12][29];
    ele[12][27] != ele[12][30];
    ele[12][27] != ele[12][31];
    ele[12][27] != ele[12][32];
    ele[12][27] != ele[12][33];
    ele[12][27] != ele[12][34];
    ele[12][27] != ele[12][35];
    ele[12][27] != ele[13][24];
    ele[12][27] != ele[13][25];
    ele[12][27] != ele[13][26];
    ele[12][27] != ele[13][27];
    ele[12][27] != ele[13][28];
    ele[12][27] != ele[13][29];
    ele[12][27] != ele[14][24];
    ele[12][27] != ele[14][25];
    ele[12][27] != ele[14][26];
    ele[12][27] != ele[14][27];
    ele[12][27] != ele[14][28];
    ele[12][27] != ele[14][29];
    ele[12][27] != ele[15][24];
    ele[12][27] != ele[15][25];
    ele[12][27] != ele[15][26];
    ele[12][27] != ele[15][27];
    ele[12][27] != ele[15][28];
    ele[12][27] != ele[15][29];
    ele[12][27] != ele[16][24];
    ele[12][27] != ele[16][25];
    ele[12][27] != ele[16][26];
    ele[12][27] != ele[16][27];
    ele[12][27] != ele[16][28];
    ele[12][27] != ele[16][29];
    ele[12][27] != ele[17][24];
    ele[12][27] != ele[17][25];
    ele[12][27] != ele[17][26];
    ele[12][27] != ele[17][27];
    ele[12][27] != ele[17][28];
    ele[12][27] != ele[17][29];
    ele[12][27] != ele[18][27];
    ele[12][27] != ele[19][27];
    ele[12][27] != ele[20][27];
    ele[12][27] != ele[21][27];
    ele[12][27] != ele[22][27];
    ele[12][27] != ele[23][27];
    ele[12][27] != ele[24][27];
    ele[12][27] != ele[25][27];
    ele[12][27] != ele[26][27];
    ele[12][27] != ele[27][27];
    ele[12][27] != ele[28][27];
    ele[12][27] != ele[29][27];
    ele[12][27] != ele[30][27];
    ele[12][27] != ele[31][27];
    ele[12][27] != ele[32][27];
    ele[12][27] != ele[33][27];
    ele[12][27] != ele[34][27];
    ele[12][27] != ele[35][27];
    ele[12][28] != ele[12][29];
    ele[12][28] != ele[12][30];
    ele[12][28] != ele[12][31];
    ele[12][28] != ele[12][32];
    ele[12][28] != ele[12][33];
    ele[12][28] != ele[12][34];
    ele[12][28] != ele[12][35];
    ele[12][28] != ele[13][24];
    ele[12][28] != ele[13][25];
    ele[12][28] != ele[13][26];
    ele[12][28] != ele[13][27];
    ele[12][28] != ele[13][28];
    ele[12][28] != ele[13][29];
    ele[12][28] != ele[14][24];
    ele[12][28] != ele[14][25];
    ele[12][28] != ele[14][26];
    ele[12][28] != ele[14][27];
    ele[12][28] != ele[14][28];
    ele[12][28] != ele[14][29];
    ele[12][28] != ele[15][24];
    ele[12][28] != ele[15][25];
    ele[12][28] != ele[15][26];
    ele[12][28] != ele[15][27];
    ele[12][28] != ele[15][28];
    ele[12][28] != ele[15][29];
    ele[12][28] != ele[16][24];
    ele[12][28] != ele[16][25];
    ele[12][28] != ele[16][26];
    ele[12][28] != ele[16][27];
    ele[12][28] != ele[16][28];
    ele[12][28] != ele[16][29];
    ele[12][28] != ele[17][24];
    ele[12][28] != ele[17][25];
    ele[12][28] != ele[17][26];
    ele[12][28] != ele[17][27];
    ele[12][28] != ele[17][28];
    ele[12][28] != ele[17][29];
    ele[12][28] != ele[18][28];
    ele[12][28] != ele[19][28];
    ele[12][28] != ele[20][28];
    ele[12][28] != ele[21][28];
    ele[12][28] != ele[22][28];
    ele[12][28] != ele[23][28];
    ele[12][28] != ele[24][28];
    ele[12][28] != ele[25][28];
    ele[12][28] != ele[26][28];
    ele[12][28] != ele[27][28];
    ele[12][28] != ele[28][28];
    ele[12][28] != ele[29][28];
    ele[12][28] != ele[30][28];
    ele[12][28] != ele[31][28];
    ele[12][28] != ele[32][28];
    ele[12][28] != ele[33][28];
    ele[12][28] != ele[34][28];
    ele[12][28] != ele[35][28];
    ele[12][29] != ele[12][30];
    ele[12][29] != ele[12][31];
    ele[12][29] != ele[12][32];
    ele[12][29] != ele[12][33];
    ele[12][29] != ele[12][34];
    ele[12][29] != ele[12][35];
    ele[12][29] != ele[13][24];
    ele[12][29] != ele[13][25];
    ele[12][29] != ele[13][26];
    ele[12][29] != ele[13][27];
    ele[12][29] != ele[13][28];
    ele[12][29] != ele[13][29];
    ele[12][29] != ele[14][24];
    ele[12][29] != ele[14][25];
    ele[12][29] != ele[14][26];
    ele[12][29] != ele[14][27];
    ele[12][29] != ele[14][28];
    ele[12][29] != ele[14][29];
    ele[12][29] != ele[15][24];
    ele[12][29] != ele[15][25];
    ele[12][29] != ele[15][26];
    ele[12][29] != ele[15][27];
    ele[12][29] != ele[15][28];
    ele[12][29] != ele[15][29];
    ele[12][29] != ele[16][24];
    ele[12][29] != ele[16][25];
    ele[12][29] != ele[16][26];
    ele[12][29] != ele[16][27];
    ele[12][29] != ele[16][28];
    ele[12][29] != ele[16][29];
    ele[12][29] != ele[17][24];
    ele[12][29] != ele[17][25];
    ele[12][29] != ele[17][26];
    ele[12][29] != ele[17][27];
    ele[12][29] != ele[17][28];
    ele[12][29] != ele[17][29];
    ele[12][29] != ele[18][29];
    ele[12][29] != ele[19][29];
    ele[12][29] != ele[20][29];
    ele[12][29] != ele[21][29];
    ele[12][29] != ele[22][29];
    ele[12][29] != ele[23][29];
    ele[12][29] != ele[24][29];
    ele[12][29] != ele[25][29];
    ele[12][29] != ele[26][29];
    ele[12][29] != ele[27][29];
    ele[12][29] != ele[28][29];
    ele[12][29] != ele[29][29];
    ele[12][29] != ele[30][29];
    ele[12][29] != ele[31][29];
    ele[12][29] != ele[32][29];
    ele[12][29] != ele[33][29];
    ele[12][29] != ele[34][29];
    ele[12][29] != ele[35][29];
    ele[12][3] != ele[12][10];
    ele[12][3] != ele[12][11];
    ele[12][3] != ele[12][12];
    ele[12][3] != ele[12][13];
    ele[12][3] != ele[12][14];
    ele[12][3] != ele[12][15];
    ele[12][3] != ele[12][16];
    ele[12][3] != ele[12][17];
    ele[12][3] != ele[12][18];
    ele[12][3] != ele[12][19];
    ele[12][3] != ele[12][20];
    ele[12][3] != ele[12][21];
    ele[12][3] != ele[12][22];
    ele[12][3] != ele[12][23];
    ele[12][3] != ele[12][24];
    ele[12][3] != ele[12][25];
    ele[12][3] != ele[12][26];
    ele[12][3] != ele[12][27];
    ele[12][3] != ele[12][28];
    ele[12][3] != ele[12][29];
    ele[12][3] != ele[12][30];
    ele[12][3] != ele[12][31];
    ele[12][3] != ele[12][32];
    ele[12][3] != ele[12][33];
    ele[12][3] != ele[12][34];
    ele[12][3] != ele[12][35];
    ele[12][3] != ele[12][4];
    ele[12][3] != ele[12][5];
    ele[12][3] != ele[12][6];
    ele[12][3] != ele[12][7];
    ele[12][3] != ele[12][8];
    ele[12][3] != ele[12][9];
    ele[12][3] != ele[13][0];
    ele[12][3] != ele[13][1];
    ele[12][3] != ele[13][2];
    ele[12][3] != ele[13][3];
    ele[12][3] != ele[13][4];
    ele[12][3] != ele[13][5];
    ele[12][3] != ele[14][0];
    ele[12][3] != ele[14][1];
    ele[12][3] != ele[14][2];
    ele[12][3] != ele[14][3];
    ele[12][3] != ele[14][4];
    ele[12][3] != ele[14][5];
    ele[12][3] != ele[15][0];
    ele[12][3] != ele[15][1];
    ele[12][3] != ele[15][2];
    ele[12][3] != ele[15][3];
    ele[12][3] != ele[15][4];
    ele[12][3] != ele[15][5];
    ele[12][3] != ele[16][0];
    ele[12][3] != ele[16][1];
    ele[12][3] != ele[16][2];
    ele[12][3] != ele[16][3];
    ele[12][3] != ele[16][4];
    ele[12][3] != ele[16][5];
    ele[12][3] != ele[17][0];
    ele[12][3] != ele[17][1];
    ele[12][3] != ele[17][2];
    ele[12][3] != ele[17][3];
    ele[12][3] != ele[17][4];
    ele[12][3] != ele[17][5];
    ele[12][3] != ele[18][3];
    ele[12][3] != ele[19][3];
    ele[12][3] != ele[20][3];
    ele[12][3] != ele[21][3];
    ele[12][3] != ele[22][3];
    ele[12][3] != ele[23][3];
    ele[12][3] != ele[24][3];
    ele[12][3] != ele[25][3];
    ele[12][3] != ele[26][3];
    ele[12][3] != ele[27][3];
    ele[12][3] != ele[28][3];
    ele[12][3] != ele[29][3];
    ele[12][3] != ele[30][3];
    ele[12][3] != ele[31][3];
    ele[12][3] != ele[32][3];
    ele[12][3] != ele[33][3];
    ele[12][3] != ele[34][3];
    ele[12][3] != ele[35][3];
    ele[12][30] != ele[12][31];
    ele[12][30] != ele[12][32];
    ele[12][30] != ele[12][33];
    ele[12][30] != ele[12][34];
    ele[12][30] != ele[12][35];
    ele[12][30] != ele[13][30];
    ele[12][30] != ele[13][31];
    ele[12][30] != ele[13][32];
    ele[12][30] != ele[13][33];
    ele[12][30] != ele[13][34];
    ele[12][30] != ele[13][35];
    ele[12][30] != ele[14][30];
    ele[12][30] != ele[14][31];
    ele[12][30] != ele[14][32];
    ele[12][30] != ele[14][33];
    ele[12][30] != ele[14][34];
    ele[12][30] != ele[14][35];
    ele[12][30] != ele[15][30];
    ele[12][30] != ele[15][31];
    ele[12][30] != ele[15][32];
    ele[12][30] != ele[15][33];
    ele[12][30] != ele[15][34];
    ele[12][30] != ele[15][35];
    ele[12][30] != ele[16][30];
    ele[12][30] != ele[16][31];
    ele[12][30] != ele[16][32];
    ele[12][30] != ele[16][33];
    ele[12][30] != ele[16][34];
    ele[12][30] != ele[16][35];
    ele[12][30] != ele[17][30];
    ele[12][30] != ele[17][31];
    ele[12][30] != ele[17][32];
    ele[12][30] != ele[17][33];
    ele[12][30] != ele[17][34];
    ele[12][30] != ele[17][35];
    ele[12][30] != ele[18][30];
    ele[12][30] != ele[19][30];
    ele[12][30] != ele[20][30];
    ele[12][30] != ele[21][30];
    ele[12][30] != ele[22][30];
    ele[12][30] != ele[23][30];
    ele[12][30] != ele[24][30];
    ele[12][30] != ele[25][30];
    ele[12][30] != ele[26][30];
    ele[12][30] != ele[27][30];
    ele[12][30] != ele[28][30];
    ele[12][30] != ele[29][30];
    ele[12][30] != ele[30][30];
    ele[12][30] != ele[31][30];
    ele[12][30] != ele[32][30];
    ele[12][30] != ele[33][30];
    ele[12][30] != ele[34][30];
    ele[12][30] != ele[35][30];
    ele[12][31] != ele[12][32];
    ele[12][31] != ele[12][33];
    ele[12][31] != ele[12][34];
    ele[12][31] != ele[12][35];
    ele[12][31] != ele[13][30];
    ele[12][31] != ele[13][31];
    ele[12][31] != ele[13][32];
    ele[12][31] != ele[13][33];
    ele[12][31] != ele[13][34];
    ele[12][31] != ele[13][35];
    ele[12][31] != ele[14][30];
    ele[12][31] != ele[14][31];
    ele[12][31] != ele[14][32];
    ele[12][31] != ele[14][33];
    ele[12][31] != ele[14][34];
    ele[12][31] != ele[14][35];
    ele[12][31] != ele[15][30];
    ele[12][31] != ele[15][31];
    ele[12][31] != ele[15][32];
    ele[12][31] != ele[15][33];
    ele[12][31] != ele[15][34];
    ele[12][31] != ele[15][35];
    ele[12][31] != ele[16][30];
    ele[12][31] != ele[16][31];
    ele[12][31] != ele[16][32];
    ele[12][31] != ele[16][33];
    ele[12][31] != ele[16][34];
    ele[12][31] != ele[16][35];
    ele[12][31] != ele[17][30];
    ele[12][31] != ele[17][31];
    ele[12][31] != ele[17][32];
    ele[12][31] != ele[17][33];
    ele[12][31] != ele[17][34];
    ele[12][31] != ele[17][35];
    ele[12][31] != ele[18][31];
    ele[12][31] != ele[19][31];
    ele[12][31] != ele[20][31];
    ele[12][31] != ele[21][31];
    ele[12][31] != ele[22][31];
    ele[12][31] != ele[23][31];
    ele[12][31] != ele[24][31];
    ele[12][31] != ele[25][31];
    ele[12][31] != ele[26][31];
    ele[12][31] != ele[27][31];
    ele[12][31] != ele[28][31];
    ele[12][31] != ele[29][31];
    ele[12][31] != ele[30][31];
    ele[12][31] != ele[31][31];
    ele[12][31] != ele[32][31];
    ele[12][31] != ele[33][31];
    ele[12][31] != ele[34][31];
    ele[12][31] != ele[35][31];
    ele[12][32] != ele[12][33];
    ele[12][32] != ele[12][34];
    ele[12][32] != ele[12][35];
    ele[12][32] != ele[13][30];
    ele[12][32] != ele[13][31];
    ele[12][32] != ele[13][32];
    ele[12][32] != ele[13][33];
    ele[12][32] != ele[13][34];
    ele[12][32] != ele[13][35];
    ele[12][32] != ele[14][30];
    ele[12][32] != ele[14][31];
    ele[12][32] != ele[14][32];
    ele[12][32] != ele[14][33];
    ele[12][32] != ele[14][34];
    ele[12][32] != ele[14][35];
    ele[12][32] != ele[15][30];
    ele[12][32] != ele[15][31];
    ele[12][32] != ele[15][32];
    ele[12][32] != ele[15][33];
    ele[12][32] != ele[15][34];
    ele[12][32] != ele[15][35];
    ele[12][32] != ele[16][30];
    ele[12][32] != ele[16][31];
    ele[12][32] != ele[16][32];
    ele[12][32] != ele[16][33];
    ele[12][32] != ele[16][34];
    ele[12][32] != ele[16][35];
    ele[12][32] != ele[17][30];
    ele[12][32] != ele[17][31];
    ele[12][32] != ele[17][32];
    ele[12][32] != ele[17][33];
    ele[12][32] != ele[17][34];
    ele[12][32] != ele[17][35];
    ele[12][32] != ele[18][32];
    ele[12][32] != ele[19][32];
    ele[12][32] != ele[20][32];
    ele[12][32] != ele[21][32];
    ele[12][32] != ele[22][32];
    ele[12][32] != ele[23][32];
    ele[12][32] != ele[24][32];
    ele[12][32] != ele[25][32];
    ele[12][32] != ele[26][32];
    ele[12][32] != ele[27][32];
    ele[12][32] != ele[28][32];
    ele[12][32] != ele[29][32];
    ele[12][32] != ele[30][32];
    ele[12][32] != ele[31][32];
    ele[12][32] != ele[32][32];
    ele[12][32] != ele[33][32];
    ele[12][32] != ele[34][32];
    ele[12][32] != ele[35][32];
    ele[12][33] != ele[12][34];
    ele[12][33] != ele[12][35];
    ele[12][33] != ele[13][30];
    ele[12][33] != ele[13][31];
    ele[12][33] != ele[13][32];
    ele[12][33] != ele[13][33];
    ele[12][33] != ele[13][34];
    ele[12][33] != ele[13][35];
    ele[12][33] != ele[14][30];
    ele[12][33] != ele[14][31];
    ele[12][33] != ele[14][32];
    ele[12][33] != ele[14][33];
    ele[12][33] != ele[14][34];
    ele[12][33] != ele[14][35];
    ele[12][33] != ele[15][30];
    ele[12][33] != ele[15][31];
    ele[12][33] != ele[15][32];
    ele[12][33] != ele[15][33];
    ele[12][33] != ele[15][34];
    ele[12][33] != ele[15][35];
    ele[12][33] != ele[16][30];
    ele[12][33] != ele[16][31];
    ele[12][33] != ele[16][32];
    ele[12][33] != ele[16][33];
    ele[12][33] != ele[16][34];
    ele[12][33] != ele[16][35];
    ele[12][33] != ele[17][30];
    ele[12][33] != ele[17][31];
    ele[12][33] != ele[17][32];
    ele[12][33] != ele[17][33];
    ele[12][33] != ele[17][34];
    ele[12][33] != ele[17][35];
    ele[12][33] != ele[18][33];
    ele[12][33] != ele[19][33];
    ele[12][33] != ele[20][33];
    ele[12][33] != ele[21][33];
    ele[12][33] != ele[22][33];
    ele[12][33] != ele[23][33];
    ele[12][33] != ele[24][33];
    ele[12][33] != ele[25][33];
    ele[12][33] != ele[26][33];
    ele[12][33] != ele[27][33];
    ele[12][33] != ele[28][33];
    ele[12][33] != ele[29][33];
    ele[12][33] != ele[30][33];
    ele[12][33] != ele[31][33];
    ele[12][33] != ele[32][33];
    ele[12][33] != ele[33][33];
    ele[12][33] != ele[34][33];
    ele[12][33] != ele[35][33];
    ele[12][34] != ele[12][35];
    ele[12][34] != ele[13][30];
    ele[12][34] != ele[13][31];
    ele[12][34] != ele[13][32];
    ele[12][34] != ele[13][33];
    ele[12][34] != ele[13][34];
    ele[12][34] != ele[13][35];
    ele[12][34] != ele[14][30];
    ele[12][34] != ele[14][31];
    ele[12][34] != ele[14][32];
    ele[12][34] != ele[14][33];
    ele[12][34] != ele[14][34];
    ele[12][34] != ele[14][35];
    ele[12][34] != ele[15][30];
    ele[12][34] != ele[15][31];
    ele[12][34] != ele[15][32];
    ele[12][34] != ele[15][33];
    ele[12][34] != ele[15][34];
    ele[12][34] != ele[15][35];
    ele[12][34] != ele[16][30];
    ele[12][34] != ele[16][31];
    ele[12][34] != ele[16][32];
    ele[12][34] != ele[16][33];
    ele[12][34] != ele[16][34];
    ele[12][34] != ele[16][35];
    ele[12][34] != ele[17][30];
    ele[12][34] != ele[17][31];
    ele[12][34] != ele[17][32];
    ele[12][34] != ele[17][33];
    ele[12][34] != ele[17][34];
    ele[12][34] != ele[17][35];
    ele[12][34] != ele[18][34];
    ele[12][34] != ele[19][34];
    ele[12][34] != ele[20][34];
    ele[12][34] != ele[21][34];
    ele[12][34] != ele[22][34];
    ele[12][34] != ele[23][34];
    ele[12][34] != ele[24][34];
    ele[12][34] != ele[25][34];
    ele[12][34] != ele[26][34];
    ele[12][34] != ele[27][34];
    ele[12][34] != ele[28][34];
    ele[12][34] != ele[29][34];
    ele[12][34] != ele[30][34];
    ele[12][34] != ele[31][34];
    ele[12][34] != ele[32][34];
    ele[12][34] != ele[33][34];
    ele[12][34] != ele[34][34];
    ele[12][34] != ele[35][34];
    ele[12][35] != ele[13][30];
    ele[12][35] != ele[13][31];
    ele[12][35] != ele[13][32];
    ele[12][35] != ele[13][33];
    ele[12][35] != ele[13][34];
    ele[12][35] != ele[13][35];
    ele[12][35] != ele[14][30];
    ele[12][35] != ele[14][31];
    ele[12][35] != ele[14][32];
    ele[12][35] != ele[14][33];
    ele[12][35] != ele[14][34];
    ele[12][35] != ele[14][35];
    ele[12][35] != ele[15][30];
    ele[12][35] != ele[15][31];
    ele[12][35] != ele[15][32];
    ele[12][35] != ele[15][33];
    ele[12][35] != ele[15][34];
    ele[12][35] != ele[15][35];
    ele[12][35] != ele[16][30];
    ele[12][35] != ele[16][31];
    ele[12][35] != ele[16][32];
    ele[12][35] != ele[16][33];
    ele[12][35] != ele[16][34];
    ele[12][35] != ele[16][35];
    ele[12][35] != ele[17][30];
    ele[12][35] != ele[17][31];
    ele[12][35] != ele[17][32];
    ele[12][35] != ele[17][33];
    ele[12][35] != ele[17][34];
    ele[12][35] != ele[17][35];
    ele[12][35] != ele[18][35];
    ele[12][35] != ele[19][35];
    ele[12][35] != ele[20][35];
    ele[12][35] != ele[21][35];
    ele[12][35] != ele[22][35];
    ele[12][35] != ele[23][35];
    ele[12][35] != ele[24][35];
    ele[12][35] != ele[25][35];
    ele[12][35] != ele[26][35];
    ele[12][35] != ele[27][35];
    ele[12][35] != ele[28][35];
    ele[12][35] != ele[29][35];
    ele[12][35] != ele[30][35];
    ele[12][35] != ele[31][35];
    ele[12][35] != ele[32][35];
    ele[12][35] != ele[33][35];
    ele[12][35] != ele[34][35];
    ele[12][35] != ele[35][35];
    ele[12][4] != ele[12][10];
    ele[12][4] != ele[12][11];
    ele[12][4] != ele[12][12];
    ele[12][4] != ele[12][13];
    ele[12][4] != ele[12][14];
    ele[12][4] != ele[12][15];
    ele[12][4] != ele[12][16];
    ele[12][4] != ele[12][17];
    ele[12][4] != ele[12][18];
    ele[12][4] != ele[12][19];
    ele[12][4] != ele[12][20];
    ele[12][4] != ele[12][21];
    ele[12][4] != ele[12][22];
    ele[12][4] != ele[12][23];
    ele[12][4] != ele[12][24];
    ele[12][4] != ele[12][25];
    ele[12][4] != ele[12][26];
    ele[12][4] != ele[12][27];
    ele[12][4] != ele[12][28];
    ele[12][4] != ele[12][29];
    ele[12][4] != ele[12][30];
    ele[12][4] != ele[12][31];
    ele[12][4] != ele[12][32];
    ele[12][4] != ele[12][33];
    ele[12][4] != ele[12][34];
    ele[12][4] != ele[12][35];
    ele[12][4] != ele[12][5];
    ele[12][4] != ele[12][6];
    ele[12][4] != ele[12][7];
    ele[12][4] != ele[12][8];
    ele[12][4] != ele[12][9];
    ele[12][4] != ele[13][0];
    ele[12][4] != ele[13][1];
    ele[12][4] != ele[13][2];
    ele[12][4] != ele[13][3];
    ele[12][4] != ele[13][4];
    ele[12][4] != ele[13][5];
    ele[12][4] != ele[14][0];
    ele[12][4] != ele[14][1];
    ele[12][4] != ele[14][2];
    ele[12][4] != ele[14][3];
    ele[12][4] != ele[14][4];
    ele[12][4] != ele[14][5];
    ele[12][4] != ele[15][0];
    ele[12][4] != ele[15][1];
    ele[12][4] != ele[15][2];
    ele[12][4] != ele[15][3];
    ele[12][4] != ele[15][4];
    ele[12][4] != ele[15][5];
    ele[12][4] != ele[16][0];
    ele[12][4] != ele[16][1];
    ele[12][4] != ele[16][2];
    ele[12][4] != ele[16][3];
    ele[12][4] != ele[16][4];
    ele[12][4] != ele[16][5];
    ele[12][4] != ele[17][0];
    ele[12][4] != ele[17][1];
    ele[12][4] != ele[17][2];
    ele[12][4] != ele[17][3];
    ele[12][4] != ele[17][4];
    ele[12][4] != ele[17][5];
    ele[12][4] != ele[18][4];
    ele[12][4] != ele[19][4];
    ele[12][4] != ele[20][4];
    ele[12][4] != ele[21][4];
    ele[12][4] != ele[22][4];
    ele[12][4] != ele[23][4];
    ele[12][4] != ele[24][4];
    ele[12][4] != ele[25][4];
    ele[12][4] != ele[26][4];
    ele[12][4] != ele[27][4];
    ele[12][4] != ele[28][4];
    ele[12][4] != ele[29][4];
    ele[12][4] != ele[30][4];
    ele[12][4] != ele[31][4];
    ele[12][4] != ele[32][4];
    ele[12][4] != ele[33][4];
    ele[12][4] != ele[34][4];
    ele[12][4] != ele[35][4];
    ele[12][5] != ele[12][10];
    ele[12][5] != ele[12][11];
    ele[12][5] != ele[12][12];
    ele[12][5] != ele[12][13];
    ele[12][5] != ele[12][14];
    ele[12][5] != ele[12][15];
    ele[12][5] != ele[12][16];
    ele[12][5] != ele[12][17];
    ele[12][5] != ele[12][18];
    ele[12][5] != ele[12][19];
    ele[12][5] != ele[12][20];
    ele[12][5] != ele[12][21];
    ele[12][5] != ele[12][22];
    ele[12][5] != ele[12][23];
    ele[12][5] != ele[12][24];
    ele[12][5] != ele[12][25];
    ele[12][5] != ele[12][26];
    ele[12][5] != ele[12][27];
    ele[12][5] != ele[12][28];
    ele[12][5] != ele[12][29];
    ele[12][5] != ele[12][30];
    ele[12][5] != ele[12][31];
    ele[12][5] != ele[12][32];
    ele[12][5] != ele[12][33];
    ele[12][5] != ele[12][34];
    ele[12][5] != ele[12][35];
    ele[12][5] != ele[12][6];
    ele[12][5] != ele[12][7];
    ele[12][5] != ele[12][8];
    ele[12][5] != ele[12][9];
    ele[12][5] != ele[13][0];
    ele[12][5] != ele[13][1];
    ele[12][5] != ele[13][2];
    ele[12][5] != ele[13][3];
    ele[12][5] != ele[13][4];
    ele[12][5] != ele[13][5];
    ele[12][5] != ele[14][0];
    ele[12][5] != ele[14][1];
    ele[12][5] != ele[14][2];
    ele[12][5] != ele[14][3];
    ele[12][5] != ele[14][4];
    ele[12][5] != ele[14][5];
    ele[12][5] != ele[15][0];
    ele[12][5] != ele[15][1];
    ele[12][5] != ele[15][2];
    ele[12][5] != ele[15][3];
    ele[12][5] != ele[15][4];
    ele[12][5] != ele[15][5];
    ele[12][5] != ele[16][0];
    ele[12][5] != ele[16][1];
    ele[12][5] != ele[16][2];
    ele[12][5] != ele[16][3];
    ele[12][5] != ele[16][4];
    ele[12][5] != ele[16][5];
    ele[12][5] != ele[17][0];
    ele[12][5] != ele[17][1];
    ele[12][5] != ele[17][2];
    ele[12][5] != ele[17][3];
    ele[12][5] != ele[17][4];
    ele[12][5] != ele[17][5];
    ele[12][5] != ele[18][5];
    ele[12][5] != ele[19][5];
    ele[12][5] != ele[20][5];
    ele[12][5] != ele[21][5];
    ele[12][5] != ele[22][5];
    ele[12][5] != ele[23][5];
    ele[12][5] != ele[24][5];
    ele[12][5] != ele[25][5];
    ele[12][5] != ele[26][5];
    ele[12][5] != ele[27][5];
    ele[12][5] != ele[28][5];
    ele[12][5] != ele[29][5];
    ele[12][5] != ele[30][5];
    ele[12][5] != ele[31][5];
    ele[12][5] != ele[32][5];
    ele[12][5] != ele[33][5];
    ele[12][5] != ele[34][5];
    ele[12][5] != ele[35][5];
    ele[12][6] != ele[12][10];
    ele[12][6] != ele[12][11];
    ele[12][6] != ele[12][12];
    ele[12][6] != ele[12][13];
    ele[12][6] != ele[12][14];
    ele[12][6] != ele[12][15];
    ele[12][6] != ele[12][16];
    ele[12][6] != ele[12][17];
    ele[12][6] != ele[12][18];
    ele[12][6] != ele[12][19];
    ele[12][6] != ele[12][20];
    ele[12][6] != ele[12][21];
    ele[12][6] != ele[12][22];
    ele[12][6] != ele[12][23];
    ele[12][6] != ele[12][24];
    ele[12][6] != ele[12][25];
    ele[12][6] != ele[12][26];
    ele[12][6] != ele[12][27];
    ele[12][6] != ele[12][28];
    ele[12][6] != ele[12][29];
    ele[12][6] != ele[12][30];
    ele[12][6] != ele[12][31];
    ele[12][6] != ele[12][32];
    ele[12][6] != ele[12][33];
    ele[12][6] != ele[12][34];
    ele[12][6] != ele[12][35];
    ele[12][6] != ele[12][7];
    ele[12][6] != ele[12][8];
    ele[12][6] != ele[12][9];
    ele[12][6] != ele[13][10];
    ele[12][6] != ele[13][11];
    ele[12][6] != ele[13][6];
    ele[12][6] != ele[13][7];
    ele[12][6] != ele[13][8];
    ele[12][6] != ele[13][9];
    ele[12][6] != ele[14][10];
    ele[12][6] != ele[14][11];
    ele[12][6] != ele[14][6];
    ele[12][6] != ele[14][7];
    ele[12][6] != ele[14][8];
    ele[12][6] != ele[14][9];
    ele[12][6] != ele[15][10];
    ele[12][6] != ele[15][11];
    ele[12][6] != ele[15][6];
    ele[12][6] != ele[15][7];
    ele[12][6] != ele[15][8];
    ele[12][6] != ele[15][9];
    ele[12][6] != ele[16][10];
    ele[12][6] != ele[16][11];
    ele[12][6] != ele[16][6];
    ele[12][6] != ele[16][7];
    ele[12][6] != ele[16][8];
    ele[12][6] != ele[16][9];
    ele[12][6] != ele[17][10];
    ele[12][6] != ele[17][11];
    ele[12][6] != ele[17][6];
    ele[12][6] != ele[17][7];
    ele[12][6] != ele[17][8];
    ele[12][6] != ele[17][9];
    ele[12][6] != ele[18][6];
    ele[12][6] != ele[19][6];
    ele[12][6] != ele[20][6];
    ele[12][6] != ele[21][6];
    ele[12][6] != ele[22][6];
    ele[12][6] != ele[23][6];
    ele[12][6] != ele[24][6];
    ele[12][6] != ele[25][6];
    ele[12][6] != ele[26][6];
    ele[12][6] != ele[27][6];
    ele[12][6] != ele[28][6];
    ele[12][6] != ele[29][6];
    ele[12][6] != ele[30][6];
    ele[12][6] != ele[31][6];
    ele[12][6] != ele[32][6];
    ele[12][6] != ele[33][6];
    ele[12][6] != ele[34][6];
    ele[12][6] != ele[35][6];
    ele[12][7] != ele[12][10];
    ele[12][7] != ele[12][11];
    ele[12][7] != ele[12][12];
    ele[12][7] != ele[12][13];
    ele[12][7] != ele[12][14];
    ele[12][7] != ele[12][15];
    ele[12][7] != ele[12][16];
    ele[12][7] != ele[12][17];
    ele[12][7] != ele[12][18];
    ele[12][7] != ele[12][19];
    ele[12][7] != ele[12][20];
    ele[12][7] != ele[12][21];
    ele[12][7] != ele[12][22];
    ele[12][7] != ele[12][23];
    ele[12][7] != ele[12][24];
    ele[12][7] != ele[12][25];
    ele[12][7] != ele[12][26];
    ele[12][7] != ele[12][27];
    ele[12][7] != ele[12][28];
    ele[12][7] != ele[12][29];
    ele[12][7] != ele[12][30];
    ele[12][7] != ele[12][31];
    ele[12][7] != ele[12][32];
    ele[12][7] != ele[12][33];
    ele[12][7] != ele[12][34];
    ele[12][7] != ele[12][35];
    ele[12][7] != ele[12][8];
    ele[12][7] != ele[12][9];
    ele[12][7] != ele[13][10];
    ele[12][7] != ele[13][11];
    ele[12][7] != ele[13][6];
    ele[12][7] != ele[13][7];
    ele[12][7] != ele[13][8];
    ele[12][7] != ele[13][9];
    ele[12][7] != ele[14][10];
    ele[12][7] != ele[14][11];
    ele[12][7] != ele[14][6];
    ele[12][7] != ele[14][7];
    ele[12][7] != ele[14][8];
    ele[12][7] != ele[14][9];
    ele[12][7] != ele[15][10];
    ele[12][7] != ele[15][11];
    ele[12][7] != ele[15][6];
    ele[12][7] != ele[15][7];
    ele[12][7] != ele[15][8];
    ele[12][7] != ele[15][9];
    ele[12][7] != ele[16][10];
    ele[12][7] != ele[16][11];
    ele[12][7] != ele[16][6];
    ele[12][7] != ele[16][7];
    ele[12][7] != ele[16][8];
    ele[12][7] != ele[16][9];
    ele[12][7] != ele[17][10];
    ele[12][7] != ele[17][11];
    ele[12][7] != ele[17][6];
    ele[12][7] != ele[17][7];
    ele[12][7] != ele[17][8];
    ele[12][7] != ele[17][9];
    ele[12][7] != ele[18][7];
    ele[12][7] != ele[19][7];
    ele[12][7] != ele[20][7];
    ele[12][7] != ele[21][7];
    ele[12][7] != ele[22][7];
    ele[12][7] != ele[23][7];
    ele[12][7] != ele[24][7];
    ele[12][7] != ele[25][7];
    ele[12][7] != ele[26][7];
    ele[12][7] != ele[27][7];
    ele[12][7] != ele[28][7];
    ele[12][7] != ele[29][7];
    ele[12][7] != ele[30][7];
    ele[12][7] != ele[31][7];
    ele[12][7] != ele[32][7];
    ele[12][7] != ele[33][7];
    ele[12][7] != ele[34][7];
    ele[12][7] != ele[35][7];
    ele[12][8] != ele[12][10];
    ele[12][8] != ele[12][11];
    ele[12][8] != ele[12][12];
    ele[12][8] != ele[12][13];
    ele[12][8] != ele[12][14];
    ele[12][8] != ele[12][15];
    ele[12][8] != ele[12][16];
    ele[12][8] != ele[12][17];
    ele[12][8] != ele[12][18];
    ele[12][8] != ele[12][19];
    ele[12][8] != ele[12][20];
    ele[12][8] != ele[12][21];
    ele[12][8] != ele[12][22];
    ele[12][8] != ele[12][23];
    ele[12][8] != ele[12][24];
    ele[12][8] != ele[12][25];
    ele[12][8] != ele[12][26];
    ele[12][8] != ele[12][27];
    ele[12][8] != ele[12][28];
    ele[12][8] != ele[12][29];
    ele[12][8] != ele[12][30];
    ele[12][8] != ele[12][31];
    ele[12][8] != ele[12][32];
    ele[12][8] != ele[12][33];
    ele[12][8] != ele[12][34];
    ele[12][8] != ele[12][35];
    ele[12][8] != ele[12][9];
    ele[12][8] != ele[13][10];
    ele[12][8] != ele[13][11];
    ele[12][8] != ele[13][6];
    ele[12][8] != ele[13][7];
    ele[12][8] != ele[13][8];
    ele[12][8] != ele[13][9];
    ele[12][8] != ele[14][10];
    ele[12][8] != ele[14][11];
    ele[12][8] != ele[14][6];
    ele[12][8] != ele[14][7];
    ele[12][8] != ele[14][8];
    ele[12][8] != ele[14][9];
    ele[12][8] != ele[15][10];
    ele[12][8] != ele[15][11];
    ele[12][8] != ele[15][6];
    ele[12][8] != ele[15][7];
    ele[12][8] != ele[15][8];
    ele[12][8] != ele[15][9];
    ele[12][8] != ele[16][10];
    ele[12][8] != ele[16][11];
    ele[12][8] != ele[16][6];
    ele[12][8] != ele[16][7];
    ele[12][8] != ele[16][8];
    ele[12][8] != ele[16][9];
    ele[12][8] != ele[17][10];
    ele[12][8] != ele[17][11];
    ele[12][8] != ele[17][6];
    ele[12][8] != ele[17][7];
    ele[12][8] != ele[17][8];
    ele[12][8] != ele[17][9];
    ele[12][8] != ele[18][8];
    ele[12][8] != ele[19][8];
    ele[12][8] != ele[20][8];
    ele[12][8] != ele[21][8];
    ele[12][8] != ele[22][8];
    ele[12][8] != ele[23][8];
    ele[12][8] != ele[24][8];
    ele[12][8] != ele[25][8];
    ele[12][8] != ele[26][8];
    ele[12][8] != ele[27][8];
    ele[12][8] != ele[28][8];
    ele[12][8] != ele[29][8];
    ele[12][8] != ele[30][8];
    ele[12][8] != ele[31][8];
    ele[12][8] != ele[32][8];
    ele[12][8] != ele[33][8];
    ele[12][8] != ele[34][8];
    ele[12][8] != ele[35][8];
    ele[12][9] != ele[12][10];
    ele[12][9] != ele[12][11];
    ele[12][9] != ele[12][12];
    ele[12][9] != ele[12][13];
    ele[12][9] != ele[12][14];
    ele[12][9] != ele[12][15];
    ele[12][9] != ele[12][16];
    ele[12][9] != ele[12][17];
    ele[12][9] != ele[12][18];
    ele[12][9] != ele[12][19];
    ele[12][9] != ele[12][20];
    ele[12][9] != ele[12][21];
    ele[12][9] != ele[12][22];
    ele[12][9] != ele[12][23];
    ele[12][9] != ele[12][24];
    ele[12][9] != ele[12][25];
    ele[12][9] != ele[12][26];
    ele[12][9] != ele[12][27];
    ele[12][9] != ele[12][28];
    ele[12][9] != ele[12][29];
    ele[12][9] != ele[12][30];
    ele[12][9] != ele[12][31];
    ele[12][9] != ele[12][32];
    ele[12][9] != ele[12][33];
    ele[12][9] != ele[12][34];
    ele[12][9] != ele[12][35];
    ele[12][9] != ele[13][10];
    ele[12][9] != ele[13][11];
    ele[12][9] != ele[13][6];
    ele[12][9] != ele[13][7];
    ele[12][9] != ele[13][8];
    ele[12][9] != ele[13][9];
    ele[12][9] != ele[14][10];
    ele[12][9] != ele[14][11];
    ele[12][9] != ele[14][6];
    ele[12][9] != ele[14][7];
    ele[12][9] != ele[14][8];
    ele[12][9] != ele[14][9];
    ele[12][9] != ele[15][10];
    ele[12][9] != ele[15][11];
    ele[12][9] != ele[15][6];
    ele[12][9] != ele[15][7];
    ele[12][9] != ele[15][8];
    ele[12][9] != ele[15][9];
    ele[12][9] != ele[16][10];
    ele[12][9] != ele[16][11];
    ele[12][9] != ele[16][6];
    ele[12][9] != ele[16][7];
    ele[12][9] != ele[16][8];
    ele[12][9] != ele[16][9];
    ele[12][9] != ele[17][10];
    ele[12][9] != ele[17][11];
    ele[12][9] != ele[17][6];
    ele[12][9] != ele[17][7];
    ele[12][9] != ele[17][8];
    ele[12][9] != ele[17][9];
    ele[12][9] != ele[18][9];
    ele[12][9] != ele[19][9];
    ele[12][9] != ele[20][9];
    ele[12][9] != ele[21][9];
    ele[12][9] != ele[22][9];
    ele[12][9] != ele[23][9];
    ele[12][9] != ele[24][9];
    ele[12][9] != ele[25][9];
    ele[12][9] != ele[26][9];
    ele[12][9] != ele[27][9];
    ele[12][9] != ele[28][9];
    ele[12][9] != ele[29][9];
    ele[12][9] != ele[30][9];
    ele[12][9] != ele[31][9];
    ele[12][9] != ele[32][9];
    ele[12][9] != ele[33][9];
    ele[12][9] != ele[34][9];
    ele[12][9] != ele[35][9];
    ele[13][0] != ele[13][1];
    ele[13][0] != ele[13][10];
    ele[13][0] != ele[13][11];
    ele[13][0] != ele[13][12];
    ele[13][0] != ele[13][13];
    ele[13][0] != ele[13][14];
    ele[13][0] != ele[13][15];
    ele[13][0] != ele[13][16];
    ele[13][0] != ele[13][17];
    ele[13][0] != ele[13][18];
    ele[13][0] != ele[13][19];
    ele[13][0] != ele[13][2];
    ele[13][0] != ele[13][20];
    ele[13][0] != ele[13][21];
    ele[13][0] != ele[13][22];
    ele[13][0] != ele[13][23];
    ele[13][0] != ele[13][24];
    ele[13][0] != ele[13][25];
    ele[13][0] != ele[13][26];
    ele[13][0] != ele[13][27];
    ele[13][0] != ele[13][28];
    ele[13][0] != ele[13][29];
    ele[13][0] != ele[13][3];
    ele[13][0] != ele[13][30];
    ele[13][0] != ele[13][31];
    ele[13][0] != ele[13][32];
    ele[13][0] != ele[13][33];
    ele[13][0] != ele[13][34];
    ele[13][0] != ele[13][35];
    ele[13][0] != ele[13][4];
    ele[13][0] != ele[13][5];
    ele[13][0] != ele[13][6];
    ele[13][0] != ele[13][7];
    ele[13][0] != ele[13][8];
    ele[13][0] != ele[13][9];
    ele[13][0] != ele[14][0];
    ele[13][0] != ele[14][1];
    ele[13][0] != ele[14][2];
    ele[13][0] != ele[14][3];
    ele[13][0] != ele[14][4];
    ele[13][0] != ele[14][5];
    ele[13][0] != ele[15][0];
    ele[13][0] != ele[15][1];
    ele[13][0] != ele[15][2];
    ele[13][0] != ele[15][3];
    ele[13][0] != ele[15][4];
    ele[13][0] != ele[15][5];
    ele[13][0] != ele[16][0];
    ele[13][0] != ele[16][1];
    ele[13][0] != ele[16][2];
    ele[13][0] != ele[16][3];
    ele[13][0] != ele[16][4];
    ele[13][0] != ele[16][5];
    ele[13][0] != ele[17][0];
    ele[13][0] != ele[17][1];
    ele[13][0] != ele[17][2];
    ele[13][0] != ele[17][3];
    ele[13][0] != ele[17][4];
    ele[13][0] != ele[17][5];
    ele[13][0] != ele[18][0];
    ele[13][0] != ele[19][0];
    ele[13][0] != ele[20][0];
    ele[13][0] != ele[21][0];
    ele[13][0] != ele[22][0];
    ele[13][0] != ele[23][0];
    ele[13][0] != ele[24][0];
    ele[13][0] != ele[25][0];
    ele[13][0] != ele[26][0];
    ele[13][0] != ele[27][0];
    ele[13][0] != ele[28][0];
    ele[13][0] != ele[29][0];
    ele[13][0] != ele[30][0];
    ele[13][0] != ele[31][0];
    ele[13][0] != ele[32][0];
    ele[13][0] != ele[33][0];
    ele[13][0] != ele[34][0];
    ele[13][0] != ele[35][0];
    ele[13][1] != ele[13][10];
    ele[13][1] != ele[13][11];
    ele[13][1] != ele[13][12];
    ele[13][1] != ele[13][13];
    ele[13][1] != ele[13][14];
    ele[13][1] != ele[13][15];
    ele[13][1] != ele[13][16];
    ele[13][1] != ele[13][17];
    ele[13][1] != ele[13][18];
    ele[13][1] != ele[13][19];
    ele[13][1] != ele[13][2];
    ele[13][1] != ele[13][20];
    ele[13][1] != ele[13][21];
    ele[13][1] != ele[13][22];
    ele[13][1] != ele[13][23];
    ele[13][1] != ele[13][24];
    ele[13][1] != ele[13][25];
    ele[13][1] != ele[13][26];
    ele[13][1] != ele[13][27];
    ele[13][1] != ele[13][28];
    ele[13][1] != ele[13][29];
    ele[13][1] != ele[13][3];
    ele[13][1] != ele[13][30];
    ele[13][1] != ele[13][31];
    ele[13][1] != ele[13][32];
    ele[13][1] != ele[13][33];
    ele[13][1] != ele[13][34];
    ele[13][1] != ele[13][35];
    ele[13][1] != ele[13][4];
    ele[13][1] != ele[13][5];
    ele[13][1] != ele[13][6];
    ele[13][1] != ele[13][7];
    ele[13][1] != ele[13][8];
    ele[13][1] != ele[13][9];
    ele[13][1] != ele[14][0];
    ele[13][1] != ele[14][1];
    ele[13][1] != ele[14][2];
    ele[13][1] != ele[14][3];
    ele[13][1] != ele[14][4];
    ele[13][1] != ele[14][5];
    ele[13][1] != ele[15][0];
    ele[13][1] != ele[15][1];
    ele[13][1] != ele[15][2];
    ele[13][1] != ele[15][3];
    ele[13][1] != ele[15][4];
    ele[13][1] != ele[15][5];
    ele[13][1] != ele[16][0];
    ele[13][1] != ele[16][1];
    ele[13][1] != ele[16][2];
    ele[13][1] != ele[16][3];
    ele[13][1] != ele[16][4];
    ele[13][1] != ele[16][5];
    ele[13][1] != ele[17][0];
    ele[13][1] != ele[17][1];
    ele[13][1] != ele[17][2];
    ele[13][1] != ele[17][3];
    ele[13][1] != ele[17][4];
    ele[13][1] != ele[17][5];
    ele[13][1] != ele[18][1];
    ele[13][1] != ele[19][1];
    ele[13][1] != ele[20][1];
    ele[13][1] != ele[21][1];
    ele[13][1] != ele[22][1];
    ele[13][1] != ele[23][1];
    ele[13][1] != ele[24][1];
    ele[13][1] != ele[25][1];
    ele[13][1] != ele[26][1];
    ele[13][1] != ele[27][1];
    ele[13][1] != ele[28][1];
    ele[13][1] != ele[29][1];
    ele[13][1] != ele[30][1];
    ele[13][1] != ele[31][1];
    ele[13][1] != ele[32][1];
    ele[13][1] != ele[33][1];
    ele[13][1] != ele[34][1];
    ele[13][1] != ele[35][1];
    ele[13][10] != ele[13][11];
    ele[13][10] != ele[13][12];
    ele[13][10] != ele[13][13];
    ele[13][10] != ele[13][14];
    ele[13][10] != ele[13][15];
    ele[13][10] != ele[13][16];
    ele[13][10] != ele[13][17];
    ele[13][10] != ele[13][18];
    ele[13][10] != ele[13][19];
    ele[13][10] != ele[13][20];
    ele[13][10] != ele[13][21];
    ele[13][10] != ele[13][22];
    ele[13][10] != ele[13][23];
    ele[13][10] != ele[13][24];
    ele[13][10] != ele[13][25];
    ele[13][10] != ele[13][26];
    ele[13][10] != ele[13][27];
    ele[13][10] != ele[13][28];
    ele[13][10] != ele[13][29];
    ele[13][10] != ele[13][30];
    ele[13][10] != ele[13][31];
    ele[13][10] != ele[13][32];
    ele[13][10] != ele[13][33];
    ele[13][10] != ele[13][34];
    ele[13][10] != ele[13][35];
    ele[13][10] != ele[14][10];
    ele[13][10] != ele[14][11];
    ele[13][10] != ele[14][6];
    ele[13][10] != ele[14][7];
    ele[13][10] != ele[14][8];
    ele[13][10] != ele[14][9];
    ele[13][10] != ele[15][10];
    ele[13][10] != ele[15][11];
    ele[13][10] != ele[15][6];
    ele[13][10] != ele[15][7];
    ele[13][10] != ele[15][8];
    ele[13][10] != ele[15][9];
    ele[13][10] != ele[16][10];
    ele[13][10] != ele[16][11];
    ele[13][10] != ele[16][6];
    ele[13][10] != ele[16][7];
    ele[13][10] != ele[16][8];
    ele[13][10] != ele[16][9];
    ele[13][10] != ele[17][10];
    ele[13][10] != ele[17][11];
    ele[13][10] != ele[17][6];
    ele[13][10] != ele[17][7];
    ele[13][10] != ele[17][8];
    ele[13][10] != ele[17][9];
    ele[13][10] != ele[18][10];
    ele[13][10] != ele[19][10];
    ele[13][10] != ele[20][10];
    ele[13][10] != ele[21][10];
    ele[13][10] != ele[22][10];
    ele[13][10] != ele[23][10];
    ele[13][10] != ele[24][10];
    ele[13][10] != ele[25][10];
    ele[13][10] != ele[26][10];
    ele[13][10] != ele[27][10];
    ele[13][10] != ele[28][10];
    ele[13][10] != ele[29][10];
    ele[13][10] != ele[30][10];
    ele[13][10] != ele[31][10];
    ele[13][10] != ele[32][10];
    ele[13][10] != ele[33][10];
    ele[13][10] != ele[34][10];
    ele[13][10] != ele[35][10];
    ele[13][11] != ele[13][12];
    ele[13][11] != ele[13][13];
    ele[13][11] != ele[13][14];
    ele[13][11] != ele[13][15];
    ele[13][11] != ele[13][16];
    ele[13][11] != ele[13][17];
    ele[13][11] != ele[13][18];
    ele[13][11] != ele[13][19];
    ele[13][11] != ele[13][20];
    ele[13][11] != ele[13][21];
    ele[13][11] != ele[13][22];
    ele[13][11] != ele[13][23];
    ele[13][11] != ele[13][24];
    ele[13][11] != ele[13][25];
    ele[13][11] != ele[13][26];
    ele[13][11] != ele[13][27];
    ele[13][11] != ele[13][28];
    ele[13][11] != ele[13][29];
    ele[13][11] != ele[13][30];
    ele[13][11] != ele[13][31];
    ele[13][11] != ele[13][32];
    ele[13][11] != ele[13][33];
    ele[13][11] != ele[13][34];
    ele[13][11] != ele[13][35];
    ele[13][11] != ele[14][10];
    ele[13][11] != ele[14][11];
    ele[13][11] != ele[14][6];
    ele[13][11] != ele[14][7];
    ele[13][11] != ele[14][8];
    ele[13][11] != ele[14][9];
    ele[13][11] != ele[15][10];
    ele[13][11] != ele[15][11];
    ele[13][11] != ele[15][6];
    ele[13][11] != ele[15][7];
    ele[13][11] != ele[15][8];
    ele[13][11] != ele[15][9];
    ele[13][11] != ele[16][10];
    ele[13][11] != ele[16][11];
    ele[13][11] != ele[16][6];
    ele[13][11] != ele[16][7];
    ele[13][11] != ele[16][8];
    ele[13][11] != ele[16][9];
    ele[13][11] != ele[17][10];
    ele[13][11] != ele[17][11];
    ele[13][11] != ele[17][6];
    ele[13][11] != ele[17][7];
    ele[13][11] != ele[17][8];
    ele[13][11] != ele[17][9];
    ele[13][11] != ele[18][11];
    ele[13][11] != ele[19][11];
    ele[13][11] != ele[20][11];
    ele[13][11] != ele[21][11];
    ele[13][11] != ele[22][11];
    ele[13][11] != ele[23][11];
    ele[13][11] != ele[24][11];
    ele[13][11] != ele[25][11];
    ele[13][11] != ele[26][11];
    ele[13][11] != ele[27][11];
    ele[13][11] != ele[28][11];
    ele[13][11] != ele[29][11];
    ele[13][11] != ele[30][11];
    ele[13][11] != ele[31][11];
    ele[13][11] != ele[32][11];
    ele[13][11] != ele[33][11];
    ele[13][11] != ele[34][11];
    ele[13][11] != ele[35][11];
    ele[13][12] != ele[13][13];
    ele[13][12] != ele[13][14];
    ele[13][12] != ele[13][15];
    ele[13][12] != ele[13][16];
    ele[13][12] != ele[13][17];
    ele[13][12] != ele[13][18];
    ele[13][12] != ele[13][19];
    ele[13][12] != ele[13][20];
    ele[13][12] != ele[13][21];
    ele[13][12] != ele[13][22];
    ele[13][12] != ele[13][23];
    ele[13][12] != ele[13][24];
    ele[13][12] != ele[13][25];
    ele[13][12] != ele[13][26];
    ele[13][12] != ele[13][27];
    ele[13][12] != ele[13][28];
    ele[13][12] != ele[13][29];
    ele[13][12] != ele[13][30];
    ele[13][12] != ele[13][31];
    ele[13][12] != ele[13][32];
    ele[13][12] != ele[13][33];
    ele[13][12] != ele[13][34];
    ele[13][12] != ele[13][35];
    ele[13][12] != ele[14][12];
    ele[13][12] != ele[14][13];
    ele[13][12] != ele[14][14];
    ele[13][12] != ele[14][15];
    ele[13][12] != ele[14][16];
    ele[13][12] != ele[14][17];
    ele[13][12] != ele[15][12];
    ele[13][12] != ele[15][13];
    ele[13][12] != ele[15][14];
    ele[13][12] != ele[15][15];
    ele[13][12] != ele[15][16];
    ele[13][12] != ele[15][17];
    ele[13][12] != ele[16][12];
    ele[13][12] != ele[16][13];
    ele[13][12] != ele[16][14];
    ele[13][12] != ele[16][15];
    ele[13][12] != ele[16][16];
    ele[13][12] != ele[16][17];
    ele[13][12] != ele[17][12];
    ele[13][12] != ele[17][13];
    ele[13][12] != ele[17][14];
    ele[13][12] != ele[17][15];
    ele[13][12] != ele[17][16];
    ele[13][12] != ele[17][17];
    ele[13][12] != ele[18][12];
    ele[13][12] != ele[19][12];
    ele[13][12] != ele[20][12];
    ele[13][12] != ele[21][12];
    ele[13][12] != ele[22][12];
    ele[13][12] != ele[23][12];
    ele[13][12] != ele[24][12];
    ele[13][12] != ele[25][12];
    ele[13][12] != ele[26][12];
    ele[13][12] != ele[27][12];
    ele[13][12] != ele[28][12];
    ele[13][12] != ele[29][12];
    ele[13][12] != ele[30][12];
    ele[13][12] != ele[31][12];
    ele[13][12] != ele[32][12];
    ele[13][12] != ele[33][12];
    ele[13][12] != ele[34][12];
    ele[13][12] != ele[35][12];
    ele[13][13] != ele[13][14];
    ele[13][13] != ele[13][15];
    ele[13][13] != ele[13][16];
    ele[13][13] != ele[13][17];
    ele[13][13] != ele[13][18];
    ele[13][13] != ele[13][19];
    ele[13][13] != ele[13][20];
    ele[13][13] != ele[13][21];
    ele[13][13] != ele[13][22];
    ele[13][13] != ele[13][23];
    ele[13][13] != ele[13][24];
    ele[13][13] != ele[13][25];
    ele[13][13] != ele[13][26];
    ele[13][13] != ele[13][27];
    ele[13][13] != ele[13][28];
    ele[13][13] != ele[13][29];
    ele[13][13] != ele[13][30];
    ele[13][13] != ele[13][31];
    ele[13][13] != ele[13][32];
    ele[13][13] != ele[13][33];
    ele[13][13] != ele[13][34];
    ele[13][13] != ele[13][35];
    ele[13][13] != ele[14][12];
    ele[13][13] != ele[14][13];
    ele[13][13] != ele[14][14];
    ele[13][13] != ele[14][15];
    ele[13][13] != ele[14][16];
    ele[13][13] != ele[14][17];
    ele[13][13] != ele[15][12];
    ele[13][13] != ele[15][13];
    ele[13][13] != ele[15][14];
    ele[13][13] != ele[15][15];
    ele[13][13] != ele[15][16];
    ele[13][13] != ele[15][17];
    ele[13][13] != ele[16][12];
    ele[13][13] != ele[16][13];
    ele[13][13] != ele[16][14];
    ele[13][13] != ele[16][15];
    ele[13][13] != ele[16][16];
    ele[13][13] != ele[16][17];
    ele[13][13] != ele[17][12];
    ele[13][13] != ele[17][13];
    ele[13][13] != ele[17][14];
    ele[13][13] != ele[17][15];
    ele[13][13] != ele[17][16];
    ele[13][13] != ele[17][17];
    ele[13][13] != ele[18][13];
    ele[13][13] != ele[19][13];
    ele[13][13] != ele[20][13];
    ele[13][13] != ele[21][13];
    ele[13][13] != ele[22][13];
    ele[13][13] != ele[23][13];
    ele[13][13] != ele[24][13];
    ele[13][13] != ele[25][13];
    ele[13][13] != ele[26][13];
    ele[13][13] != ele[27][13];
    ele[13][13] != ele[28][13];
    ele[13][13] != ele[29][13];
    ele[13][13] != ele[30][13];
    ele[13][13] != ele[31][13];
    ele[13][13] != ele[32][13];
    ele[13][13] != ele[33][13];
    ele[13][13] != ele[34][13];
    ele[13][13] != ele[35][13];
    ele[13][14] != ele[13][15];
    ele[13][14] != ele[13][16];
    ele[13][14] != ele[13][17];
    ele[13][14] != ele[13][18];
    ele[13][14] != ele[13][19];
    ele[13][14] != ele[13][20];
    ele[13][14] != ele[13][21];
    ele[13][14] != ele[13][22];
    ele[13][14] != ele[13][23];
    ele[13][14] != ele[13][24];
    ele[13][14] != ele[13][25];
    ele[13][14] != ele[13][26];
    ele[13][14] != ele[13][27];
    ele[13][14] != ele[13][28];
    ele[13][14] != ele[13][29];
    ele[13][14] != ele[13][30];
    ele[13][14] != ele[13][31];
    ele[13][14] != ele[13][32];
    ele[13][14] != ele[13][33];
    ele[13][14] != ele[13][34];
    ele[13][14] != ele[13][35];
    ele[13][14] != ele[14][12];
    ele[13][14] != ele[14][13];
    ele[13][14] != ele[14][14];
    ele[13][14] != ele[14][15];
    ele[13][14] != ele[14][16];
    ele[13][14] != ele[14][17];
    ele[13][14] != ele[15][12];
    ele[13][14] != ele[15][13];
    ele[13][14] != ele[15][14];
    ele[13][14] != ele[15][15];
    ele[13][14] != ele[15][16];
    ele[13][14] != ele[15][17];
    ele[13][14] != ele[16][12];
    ele[13][14] != ele[16][13];
    ele[13][14] != ele[16][14];
    ele[13][14] != ele[16][15];
    ele[13][14] != ele[16][16];
    ele[13][14] != ele[16][17];
    ele[13][14] != ele[17][12];
    ele[13][14] != ele[17][13];
    ele[13][14] != ele[17][14];
    ele[13][14] != ele[17][15];
    ele[13][14] != ele[17][16];
    ele[13][14] != ele[17][17];
    ele[13][14] != ele[18][14];
    ele[13][14] != ele[19][14];
    ele[13][14] != ele[20][14];
    ele[13][14] != ele[21][14];
    ele[13][14] != ele[22][14];
    ele[13][14] != ele[23][14];
    ele[13][14] != ele[24][14];
    ele[13][14] != ele[25][14];
    ele[13][14] != ele[26][14];
    ele[13][14] != ele[27][14];
    ele[13][14] != ele[28][14];
    ele[13][14] != ele[29][14];
    ele[13][14] != ele[30][14];
    ele[13][14] != ele[31][14];
    ele[13][14] != ele[32][14];
    ele[13][14] != ele[33][14];
    ele[13][14] != ele[34][14];
    ele[13][14] != ele[35][14];
    ele[13][15] != ele[13][16];
    ele[13][15] != ele[13][17];
    ele[13][15] != ele[13][18];
    ele[13][15] != ele[13][19];
    ele[13][15] != ele[13][20];
    ele[13][15] != ele[13][21];
    ele[13][15] != ele[13][22];
    ele[13][15] != ele[13][23];
    ele[13][15] != ele[13][24];
    ele[13][15] != ele[13][25];
    ele[13][15] != ele[13][26];
    ele[13][15] != ele[13][27];
    ele[13][15] != ele[13][28];
    ele[13][15] != ele[13][29];
    ele[13][15] != ele[13][30];
    ele[13][15] != ele[13][31];
    ele[13][15] != ele[13][32];
    ele[13][15] != ele[13][33];
    ele[13][15] != ele[13][34];
    ele[13][15] != ele[13][35];
    ele[13][15] != ele[14][12];
    ele[13][15] != ele[14][13];
    ele[13][15] != ele[14][14];
    ele[13][15] != ele[14][15];
    ele[13][15] != ele[14][16];
    ele[13][15] != ele[14][17];
    ele[13][15] != ele[15][12];
    ele[13][15] != ele[15][13];
    ele[13][15] != ele[15][14];
    ele[13][15] != ele[15][15];
    ele[13][15] != ele[15][16];
    ele[13][15] != ele[15][17];
    ele[13][15] != ele[16][12];
    ele[13][15] != ele[16][13];
    ele[13][15] != ele[16][14];
    ele[13][15] != ele[16][15];
    ele[13][15] != ele[16][16];
    ele[13][15] != ele[16][17];
    ele[13][15] != ele[17][12];
    ele[13][15] != ele[17][13];
    ele[13][15] != ele[17][14];
    ele[13][15] != ele[17][15];
    ele[13][15] != ele[17][16];
    ele[13][15] != ele[17][17];
    ele[13][15] != ele[18][15];
    ele[13][15] != ele[19][15];
    ele[13][15] != ele[20][15];
    ele[13][15] != ele[21][15];
    ele[13][15] != ele[22][15];
    ele[13][15] != ele[23][15];
    ele[13][15] != ele[24][15];
    ele[13][15] != ele[25][15];
    ele[13][15] != ele[26][15];
    ele[13][15] != ele[27][15];
    ele[13][15] != ele[28][15];
    ele[13][15] != ele[29][15];
    ele[13][15] != ele[30][15];
    ele[13][15] != ele[31][15];
    ele[13][15] != ele[32][15];
    ele[13][15] != ele[33][15];
    ele[13][15] != ele[34][15];
    ele[13][15] != ele[35][15];
    ele[13][16] != ele[13][17];
    ele[13][16] != ele[13][18];
    ele[13][16] != ele[13][19];
    ele[13][16] != ele[13][20];
    ele[13][16] != ele[13][21];
    ele[13][16] != ele[13][22];
    ele[13][16] != ele[13][23];
    ele[13][16] != ele[13][24];
    ele[13][16] != ele[13][25];
    ele[13][16] != ele[13][26];
    ele[13][16] != ele[13][27];
    ele[13][16] != ele[13][28];
    ele[13][16] != ele[13][29];
    ele[13][16] != ele[13][30];
    ele[13][16] != ele[13][31];
    ele[13][16] != ele[13][32];
    ele[13][16] != ele[13][33];
    ele[13][16] != ele[13][34];
    ele[13][16] != ele[13][35];
    ele[13][16] != ele[14][12];
    ele[13][16] != ele[14][13];
    ele[13][16] != ele[14][14];
    ele[13][16] != ele[14][15];
    ele[13][16] != ele[14][16];
    ele[13][16] != ele[14][17];
    ele[13][16] != ele[15][12];
    ele[13][16] != ele[15][13];
    ele[13][16] != ele[15][14];
    ele[13][16] != ele[15][15];
    ele[13][16] != ele[15][16];
    ele[13][16] != ele[15][17];
    ele[13][16] != ele[16][12];
    ele[13][16] != ele[16][13];
    ele[13][16] != ele[16][14];
    ele[13][16] != ele[16][15];
    ele[13][16] != ele[16][16];
    ele[13][16] != ele[16][17];
    ele[13][16] != ele[17][12];
    ele[13][16] != ele[17][13];
    ele[13][16] != ele[17][14];
    ele[13][16] != ele[17][15];
    ele[13][16] != ele[17][16];
    ele[13][16] != ele[17][17];
    ele[13][16] != ele[18][16];
    ele[13][16] != ele[19][16];
    ele[13][16] != ele[20][16];
    ele[13][16] != ele[21][16];
    ele[13][16] != ele[22][16];
    ele[13][16] != ele[23][16];
    ele[13][16] != ele[24][16];
    ele[13][16] != ele[25][16];
    ele[13][16] != ele[26][16];
    ele[13][16] != ele[27][16];
    ele[13][16] != ele[28][16];
    ele[13][16] != ele[29][16];
    ele[13][16] != ele[30][16];
    ele[13][16] != ele[31][16];
    ele[13][16] != ele[32][16];
    ele[13][16] != ele[33][16];
    ele[13][16] != ele[34][16];
    ele[13][16] != ele[35][16];
    ele[13][17] != ele[13][18];
    ele[13][17] != ele[13][19];
    ele[13][17] != ele[13][20];
    ele[13][17] != ele[13][21];
    ele[13][17] != ele[13][22];
    ele[13][17] != ele[13][23];
    ele[13][17] != ele[13][24];
    ele[13][17] != ele[13][25];
    ele[13][17] != ele[13][26];
    ele[13][17] != ele[13][27];
    ele[13][17] != ele[13][28];
    ele[13][17] != ele[13][29];
    ele[13][17] != ele[13][30];
    ele[13][17] != ele[13][31];
    ele[13][17] != ele[13][32];
    ele[13][17] != ele[13][33];
    ele[13][17] != ele[13][34];
    ele[13][17] != ele[13][35];
    ele[13][17] != ele[14][12];
    ele[13][17] != ele[14][13];
    ele[13][17] != ele[14][14];
    ele[13][17] != ele[14][15];
    ele[13][17] != ele[14][16];
    ele[13][17] != ele[14][17];
    ele[13][17] != ele[15][12];
    ele[13][17] != ele[15][13];
    ele[13][17] != ele[15][14];
    ele[13][17] != ele[15][15];
    ele[13][17] != ele[15][16];
    ele[13][17] != ele[15][17];
    ele[13][17] != ele[16][12];
    ele[13][17] != ele[16][13];
    ele[13][17] != ele[16][14];
    ele[13][17] != ele[16][15];
    ele[13][17] != ele[16][16];
    ele[13][17] != ele[16][17];
    ele[13][17] != ele[17][12];
    ele[13][17] != ele[17][13];
    ele[13][17] != ele[17][14];
    ele[13][17] != ele[17][15];
    ele[13][17] != ele[17][16];
    ele[13][17] != ele[17][17];
    ele[13][17] != ele[18][17];
    ele[13][17] != ele[19][17];
    ele[13][17] != ele[20][17];
    ele[13][17] != ele[21][17];
    ele[13][17] != ele[22][17];
    ele[13][17] != ele[23][17];
    ele[13][17] != ele[24][17];
    ele[13][17] != ele[25][17];
    ele[13][17] != ele[26][17];
    ele[13][17] != ele[27][17];
    ele[13][17] != ele[28][17];
    ele[13][17] != ele[29][17];
    ele[13][17] != ele[30][17];
    ele[13][17] != ele[31][17];
    ele[13][17] != ele[32][17];
    ele[13][17] != ele[33][17];
    ele[13][17] != ele[34][17];
    ele[13][17] != ele[35][17];
    ele[13][18] != ele[13][19];
    ele[13][18] != ele[13][20];
    ele[13][18] != ele[13][21];
    ele[13][18] != ele[13][22];
    ele[13][18] != ele[13][23];
    ele[13][18] != ele[13][24];
    ele[13][18] != ele[13][25];
    ele[13][18] != ele[13][26];
    ele[13][18] != ele[13][27];
    ele[13][18] != ele[13][28];
    ele[13][18] != ele[13][29];
    ele[13][18] != ele[13][30];
    ele[13][18] != ele[13][31];
    ele[13][18] != ele[13][32];
    ele[13][18] != ele[13][33];
    ele[13][18] != ele[13][34];
    ele[13][18] != ele[13][35];
    ele[13][18] != ele[14][18];
    ele[13][18] != ele[14][19];
    ele[13][18] != ele[14][20];
    ele[13][18] != ele[14][21];
    ele[13][18] != ele[14][22];
    ele[13][18] != ele[14][23];
    ele[13][18] != ele[15][18];
    ele[13][18] != ele[15][19];
    ele[13][18] != ele[15][20];
    ele[13][18] != ele[15][21];
    ele[13][18] != ele[15][22];
    ele[13][18] != ele[15][23];
    ele[13][18] != ele[16][18];
    ele[13][18] != ele[16][19];
    ele[13][18] != ele[16][20];
    ele[13][18] != ele[16][21];
    ele[13][18] != ele[16][22];
    ele[13][18] != ele[16][23];
    ele[13][18] != ele[17][18];
    ele[13][18] != ele[17][19];
    ele[13][18] != ele[17][20];
    ele[13][18] != ele[17][21];
    ele[13][18] != ele[17][22];
    ele[13][18] != ele[17][23];
    ele[13][18] != ele[18][18];
    ele[13][18] != ele[19][18];
    ele[13][18] != ele[20][18];
    ele[13][18] != ele[21][18];
    ele[13][18] != ele[22][18];
    ele[13][18] != ele[23][18];
    ele[13][18] != ele[24][18];
    ele[13][18] != ele[25][18];
    ele[13][18] != ele[26][18];
    ele[13][18] != ele[27][18];
    ele[13][18] != ele[28][18];
    ele[13][18] != ele[29][18];
    ele[13][18] != ele[30][18];
    ele[13][18] != ele[31][18];
    ele[13][18] != ele[32][18];
    ele[13][18] != ele[33][18];
    ele[13][18] != ele[34][18];
    ele[13][18] != ele[35][18];
    ele[13][19] != ele[13][20];
    ele[13][19] != ele[13][21];
    ele[13][19] != ele[13][22];
    ele[13][19] != ele[13][23];
    ele[13][19] != ele[13][24];
    ele[13][19] != ele[13][25];
    ele[13][19] != ele[13][26];
    ele[13][19] != ele[13][27];
    ele[13][19] != ele[13][28];
    ele[13][19] != ele[13][29];
    ele[13][19] != ele[13][30];
    ele[13][19] != ele[13][31];
    ele[13][19] != ele[13][32];
    ele[13][19] != ele[13][33];
    ele[13][19] != ele[13][34];
    ele[13][19] != ele[13][35];
    ele[13][19] != ele[14][18];
    ele[13][19] != ele[14][19];
    ele[13][19] != ele[14][20];
    ele[13][19] != ele[14][21];
    ele[13][19] != ele[14][22];
    ele[13][19] != ele[14][23];
    ele[13][19] != ele[15][18];
    ele[13][19] != ele[15][19];
    ele[13][19] != ele[15][20];
    ele[13][19] != ele[15][21];
    ele[13][19] != ele[15][22];
    ele[13][19] != ele[15][23];
    ele[13][19] != ele[16][18];
    ele[13][19] != ele[16][19];
    ele[13][19] != ele[16][20];
    ele[13][19] != ele[16][21];
    ele[13][19] != ele[16][22];
    ele[13][19] != ele[16][23];
    ele[13][19] != ele[17][18];
    ele[13][19] != ele[17][19];
    ele[13][19] != ele[17][20];
    ele[13][19] != ele[17][21];
    ele[13][19] != ele[17][22];
    ele[13][19] != ele[17][23];
    ele[13][19] != ele[18][19];
    ele[13][19] != ele[19][19];
    ele[13][19] != ele[20][19];
    ele[13][19] != ele[21][19];
    ele[13][19] != ele[22][19];
    ele[13][19] != ele[23][19];
    ele[13][19] != ele[24][19];
    ele[13][19] != ele[25][19];
    ele[13][19] != ele[26][19];
    ele[13][19] != ele[27][19];
    ele[13][19] != ele[28][19];
    ele[13][19] != ele[29][19];
    ele[13][19] != ele[30][19];
    ele[13][19] != ele[31][19];
    ele[13][19] != ele[32][19];
    ele[13][19] != ele[33][19];
    ele[13][19] != ele[34][19];
    ele[13][19] != ele[35][19];
    ele[13][2] != ele[13][10];
    ele[13][2] != ele[13][11];
    ele[13][2] != ele[13][12];
    ele[13][2] != ele[13][13];
    ele[13][2] != ele[13][14];
    ele[13][2] != ele[13][15];
    ele[13][2] != ele[13][16];
    ele[13][2] != ele[13][17];
    ele[13][2] != ele[13][18];
    ele[13][2] != ele[13][19];
    ele[13][2] != ele[13][20];
    ele[13][2] != ele[13][21];
    ele[13][2] != ele[13][22];
    ele[13][2] != ele[13][23];
    ele[13][2] != ele[13][24];
    ele[13][2] != ele[13][25];
    ele[13][2] != ele[13][26];
    ele[13][2] != ele[13][27];
    ele[13][2] != ele[13][28];
    ele[13][2] != ele[13][29];
    ele[13][2] != ele[13][3];
    ele[13][2] != ele[13][30];
    ele[13][2] != ele[13][31];
    ele[13][2] != ele[13][32];
    ele[13][2] != ele[13][33];
    ele[13][2] != ele[13][34];
    ele[13][2] != ele[13][35];
    ele[13][2] != ele[13][4];
    ele[13][2] != ele[13][5];
    ele[13][2] != ele[13][6];
    ele[13][2] != ele[13][7];
    ele[13][2] != ele[13][8];
    ele[13][2] != ele[13][9];
    ele[13][2] != ele[14][0];
    ele[13][2] != ele[14][1];
    ele[13][2] != ele[14][2];
    ele[13][2] != ele[14][3];
    ele[13][2] != ele[14][4];
    ele[13][2] != ele[14][5];
    ele[13][2] != ele[15][0];
    ele[13][2] != ele[15][1];
    ele[13][2] != ele[15][2];
    ele[13][2] != ele[15][3];
    ele[13][2] != ele[15][4];
    ele[13][2] != ele[15][5];
    ele[13][2] != ele[16][0];
    ele[13][2] != ele[16][1];
    ele[13][2] != ele[16][2];
    ele[13][2] != ele[16][3];
    ele[13][2] != ele[16][4];
    ele[13][2] != ele[16][5];
    ele[13][2] != ele[17][0];
    ele[13][2] != ele[17][1];
    ele[13][2] != ele[17][2];
    ele[13][2] != ele[17][3];
    ele[13][2] != ele[17][4];
    ele[13][2] != ele[17][5];
    ele[13][2] != ele[18][2];
    ele[13][2] != ele[19][2];
    ele[13][2] != ele[20][2];
    ele[13][2] != ele[21][2];
    ele[13][2] != ele[22][2];
    ele[13][2] != ele[23][2];
    ele[13][2] != ele[24][2];
    ele[13][2] != ele[25][2];
    ele[13][2] != ele[26][2];
    ele[13][2] != ele[27][2];
    ele[13][2] != ele[28][2];
    ele[13][2] != ele[29][2];
    ele[13][2] != ele[30][2];
    ele[13][2] != ele[31][2];
    ele[13][2] != ele[32][2];
    ele[13][2] != ele[33][2];
    ele[13][2] != ele[34][2];
    ele[13][2] != ele[35][2];
    ele[13][20] != ele[13][21];
    ele[13][20] != ele[13][22];
    ele[13][20] != ele[13][23];
    ele[13][20] != ele[13][24];
    ele[13][20] != ele[13][25];
    ele[13][20] != ele[13][26];
    ele[13][20] != ele[13][27];
    ele[13][20] != ele[13][28];
    ele[13][20] != ele[13][29];
    ele[13][20] != ele[13][30];
    ele[13][20] != ele[13][31];
    ele[13][20] != ele[13][32];
    ele[13][20] != ele[13][33];
    ele[13][20] != ele[13][34];
    ele[13][20] != ele[13][35];
    ele[13][20] != ele[14][18];
    ele[13][20] != ele[14][19];
    ele[13][20] != ele[14][20];
    ele[13][20] != ele[14][21];
    ele[13][20] != ele[14][22];
    ele[13][20] != ele[14][23];
    ele[13][20] != ele[15][18];
    ele[13][20] != ele[15][19];
    ele[13][20] != ele[15][20];
    ele[13][20] != ele[15][21];
    ele[13][20] != ele[15][22];
    ele[13][20] != ele[15][23];
    ele[13][20] != ele[16][18];
    ele[13][20] != ele[16][19];
    ele[13][20] != ele[16][20];
    ele[13][20] != ele[16][21];
    ele[13][20] != ele[16][22];
    ele[13][20] != ele[16][23];
    ele[13][20] != ele[17][18];
    ele[13][20] != ele[17][19];
    ele[13][20] != ele[17][20];
    ele[13][20] != ele[17][21];
    ele[13][20] != ele[17][22];
    ele[13][20] != ele[17][23];
    ele[13][20] != ele[18][20];
    ele[13][20] != ele[19][20];
    ele[13][20] != ele[20][20];
    ele[13][20] != ele[21][20];
    ele[13][20] != ele[22][20];
    ele[13][20] != ele[23][20];
    ele[13][20] != ele[24][20];
    ele[13][20] != ele[25][20];
    ele[13][20] != ele[26][20];
    ele[13][20] != ele[27][20];
    ele[13][20] != ele[28][20];
    ele[13][20] != ele[29][20];
    ele[13][20] != ele[30][20];
    ele[13][20] != ele[31][20];
    ele[13][20] != ele[32][20];
    ele[13][20] != ele[33][20];
    ele[13][20] != ele[34][20];
    ele[13][20] != ele[35][20];
    ele[13][21] != ele[13][22];
    ele[13][21] != ele[13][23];
    ele[13][21] != ele[13][24];
    ele[13][21] != ele[13][25];
    ele[13][21] != ele[13][26];
    ele[13][21] != ele[13][27];
    ele[13][21] != ele[13][28];
    ele[13][21] != ele[13][29];
    ele[13][21] != ele[13][30];
    ele[13][21] != ele[13][31];
    ele[13][21] != ele[13][32];
    ele[13][21] != ele[13][33];
    ele[13][21] != ele[13][34];
    ele[13][21] != ele[13][35];
    ele[13][21] != ele[14][18];
    ele[13][21] != ele[14][19];
    ele[13][21] != ele[14][20];
    ele[13][21] != ele[14][21];
    ele[13][21] != ele[14][22];
    ele[13][21] != ele[14][23];
    ele[13][21] != ele[15][18];
    ele[13][21] != ele[15][19];
    ele[13][21] != ele[15][20];
    ele[13][21] != ele[15][21];
    ele[13][21] != ele[15][22];
    ele[13][21] != ele[15][23];
    ele[13][21] != ele[16][18];
    ele[13][21] != ele[16][19];
    ele[13][21] != ele[16][20];
    ele[13][21] != ele[16][21];
    ele[13][21] != ele[16][22];
    ele[13][21] != ele[16][23];
    ele[13][21] != ele[17][18];
    ele[13][21] != ele[17][19];
    ele[13][21] != ele[17][20];
    ele[13][21] != ele[17][21];
    ele[13][21] != ele[17][22];
    ele[13][21] != ele[17][23];
    ele[13][21] != ele[18][21];
    ele[13][21] != ele[19][21];
    ele[13][21] != ele[20][21];
    ele[13][21] != ele[21][21];
    ele[13][21] != ele[22][21];
    ele[13][21] != ele[23][21];
    ele[13][21] != ele[24][21];
    ele[13][21] != ele[25][21];
    ele[13][21] != ele[26][21];
    ele[13][21] != ele[27][21];
    ele[13][21] != ele[28][21];
    ele[13][21] != ele[29][21];
    ele[13][21] != ele[30][21];
    ele[13][21] != ele[31][21];
    ele[13][21] != ele[32][21];
    ele[13][21] != ele[33][21];
    ele[13][21] != ele[34][21];
    ele[13][21] != ele[35][21];
    ele[13][22] != ele[13][23];
    ele[13][22] != ele[13][24];
    ele[13][22] != ele[13][25];
    ele[13][22] != ele[13][26];
    ele[13][22] != ele[13][27];
    ele[13][22] != ele[13][28];
    ele[13][22] != ele[13][29];
    ele[13][22] != ele[13][30];
    ele[13][22] != ele[13][31];
    ele[13][22] != ele[13][32];
    ele[13][22] != ele[13][33];
    ele[13][22] != ele[13][34];
    ele[13][22] != ele[13][35];
    ele[13][22] != ele[14][18];
    ele[13][22] != ele[14][19];
    ele[13][22] != ele[14][20];
    ele[13][22] != ele[14][21];
    ele[13][22] != ele[14][22];
    ele[13][22] != ele[14][23];
    ele[13][22] != ele[15][18];
    ele[13][22] != ele[15][19];
    ele[13][22] != ele[15][20];
    ele[13][22] != ele[15][21];
    ele[13][22] != ele[15][22];
    ele[13][22] != ele[15][23];
    ele[13][22] != ele[16][18];
    ele[13][22] != ele[16][19];
    ele[13][22] != ele[16][20];
    ele[13][22] != ele[16][21];
    ele[13][22] != ele[16][22];
    ele[13][22] != ele[16][23];
    ele[13][22] != ele[17][18];
    ele[13][22] != ele[17][19];
    ele[13][22] != ele[17][20];
    ele[13][22] != ele[17][21];
    ele[13][22] != ele[17][22];
    ele[13][22] != ele[17][23];
    ele[13][22] != ele[18][22];
    ele[13][22] != ele[19][22];
    ele[13][22] != ele[20][22];
    ele[13][22] != ele[21][22];
    ele[13][22] != ele[22][22];
    ele[13][22] != ele[23][22];
    ele[13][22] != ele[24][22];
    ele[13][22] != ele[25][22];
    ele[13][22] != ele[26][22];
    ele[13][22] != ele[27][22];
    ele[13][22] != ele[28][22];
    ele[13][22] != ele[29][22];
    ele[13][22] != ele[30][22];
    ele[13][22] != ele[31][22];
    ele[13][22] != ele[32][22];
    ele[13][22] != ele[33][22];
    ele[13][22] != ele[34][22];
    ele[13][22] != ele[35][22];
    ele[13][23] != ele[13][24];
    ele[13][23] != ele[13][25];
    ele[13][23] != ele[13][26];
    ele[13][23] != ele[13][27];
    ele[13][23] != ele[13][28];
    ele[13][23] != ele[13][29];
    ele[13][23] != ele[13][30];
    ele[13][23] != ele[13][31];
    ele[13][23] != ele[13][32];
    ele[13][23] != ele[13][33];
    ele[13][23] != ele[13][34];
    ele[13][23] != ele[13][35];
    ele[13][23] != ele[14][18];
    ele[13][23] != ele[14][19];
    ele[13][23] != ele[14][20];
    ele[13][23] != ele[14][21];
    ele[13][23] != ele[14][22];
    ele[13][23] != ele[14][23];
    ele[13][23] != ele[15][18];
    ele[13][23] != ele[15][19];
    ele[13][23] != ele[15][20];
    ele[13][23] != ele[15][21];
    ele[13][23] != ele[15][22];
    ele[13][23] != ele[15][23];
    ele[13][23] != ele[16][18];
    ele[13][23] != ele[16][19];
    ele[13][23] != ele[16][20];
    ele[13][23] != ele[16][21];
    ele[13][23] != ele[16][22];
    ele[13][23] != ele[16][23];
    ele[13][23] != ele[17][18];
    ele[13][23] != ele[17][19];
    ele[13][23] != ele[17][20];
    ele[13][23] != ele[17][21];
    ele[13][23] != ele[17][22];
    ele[13][23] != ele[17][23];
    ele[13][23] != ele[18][23];
    ele[13][23] != ele[19][23];
    ele[13][23] != ele[20][23];
    ele[13][23] != ele[21][23];
    ele[13][23] != ele[22][23];
    ele[13][23] != ele[23][23];
    ele[13][23] != ele[24][23];
    ele[13][23] != ele[25][23];
    ele[13][23] != ele[26][23];
    ele[13][23] != ele[27][23];
    ele[13][23] != ele[28][23];
    ele[13][23] != ele[29][23];
    ele[13][23] != ele[30][23];
    ele[13][23] != ele[31][23];
    ele[13][23] != ele[32][23];
    ele[13][23] != ele[33][23];
    ele[13][23] != ele[34][23];
    ele[13][23] != ele[35][23];
    ele[13][24] != ele[13][25];
    ele[13][24] != ele[13][26];
    ele[13][24] != ele[13][27];
    ele[13][24] != ele[13][28];
    ele[13][24] != ele[13][29];
    ele[13][24] != ele[13][30];
    ele[13][24] != ele[13][31];
    ele[13][24] != ele[13][32];
    ele[13][24] != ele[13][33];
    ele[13][24] != ele[13][34];
    ele[13][24] != ele[13][35];
    ele[13][24] != ele[14][24];
    ele[13][24] != ele[14][25];
    ele[13][24] != ele[14][26];
    ele[13][24] != ele[14][27];
    ele[13][24] != ele[14][28];
    ele[13][24] != ele[14][29];
    ele[13][24] != ele[15][24];
    ele[13][24] != ele[15][25];
    ele[13][24] != ele[15][26];
    ele[13][24] != ele[15][27];
    ele[13][24] != ele[15][28];
    ele[13][24] != ele[15][29];
    ele[13][24] != ele[16][24];
    ele[13][24] != ele[16][25];
    ele[13][24] != ele[16][26];
    ele[13][24] != ele[16][27];
    ele[13][24] != ele[16][28];
    ele[13][24] != ele[16][29];
    ele[13][24] != ele[17][24];
    ele[13][24] != ele[17][25];
    ele[13][24] != ele[17][26];
    ele[13][24] != ele[17][27];
    ele[13][24] != ele[17][28];
    ele[13][24] != ele[17][29];
    ele[13][24] != ele[18][24];
    ele[13][24] != ele[19][24];
    ele[13][24] != ele[20][24];
    ele[13][24] != ele[21][24];
    ele[13][24] != ele[22][24];
    ele[13][24] != ele[23][24];
    ele[13][24] != ele[24][24];
    ele[13][24] != ele[25][24];
    ele[13][24] != ele[26][24];
    ele[13][24] != ele[27][24];
    ele[13][24] != ele[28][24];
    ele[13][24] != ele[29][24];
    ele[13][24] != ele[30][24];
    ele[13][24] != ele[31][24];
    ele[13][24] != ele[32][24];
    ele[13][24] != ele[33][24];
    ele[13][24] != ele[34][24];
    ele[13][24] != ele[35][24];
    ele[13][25] != ele[13][26];
    ele[13][25] != ele[13][27];
    ele[13][25] != ele[13][28];
    ele[13][25] != ele[13][29];
    ele[13][25] != ele[13][30];
    ele[13][25] != ele[13][31];
    ele[13][25] != ele[13][32];
    ele[13][25] != ele[13][33];
    ele[13][25] != ele[13][34];
    ele[13][25] != ele[13][35];
    ele[13][25] != ele[14][24];
    ele[13][25] != ele[14][25];
    ele[13][25] != ele[14][26];
    ele[13][25] != ele[14][27];
    ele[13][25] != ele[14][28];
    ele[13][25] != ele[14][29];
    ele[13][25] != ele[15][24];
    ele[13][25] != ele[15][25];
    ele[13][25] != ele[15][26];
    ele[13][25] != ele[15][27];
    ele[13][25] != ele[15][28];
    ele[13][25] != ele[15][29];
    ele[13][25] != ele[16][24];
    ele[13][25] != ele[16][25];
    ele[13][25] != ele[16][26];
    ele[13][25] != ele[16][27];
    ele[13][25] != ele[16][28];
    ele[13][25] != ele[16][29];
    ele[13][25] != ele[17][24];
    ele[13][25] != ele[17][25];
    ele[13][25] != ele[17][26];
    ele[13][25] != ele[17][27];
    ele[13][25] != ele[17][28];
    ele[13][25] != ele[17][29];
    ele[13][25] != ele[18][25];
    ele[13][25] != ele[19][25];
    ele[13][25] != ele[20][25];
    ele[13][25] != ele[21][25];
    ele[13][25] != ele[22][25];
    ele[13][25] != ele[23][25];
    ele[13][25] != ele[24][25];
    ele[13][25] != ele[25][25];
    ele[13][25] != ele[26][25];
    ele[13][25] != ele[27][25];
    ele[13][25] != ele[28][25];
    ele[13][25] != ele[29][25];
    ele[13][25] != ele[30][25];
    ele[13][25] != ele[31][25];
    ele[13][25] != ele[32][25];
    ele[13][25] != ele[33][25];
    ele[13][25] != ele[34][25];
    ele[13][25] != ele[35][25];
    ele[13][26] != ele[13][27];
    ele[13][26] != ele[13][28];
    ele[13][26] != ele[13][29];
    ele[13][26] != ele[13][30];
    ele[13][26] != ele[13][31];
    ele[13][26] != ele[13][32];
    ele[13][26] != ele[13][33];
    ele[13][26] != ele[13][34];
    ele[13][26] != ele[13][35];
    ele[13][26] != ele[14][24];
    ele[13][26] != ele[14][25];
    ele[13][26] != ele[14][26];
    ele[13][26] != ele[14][27];
    ele[13][26] != ele[14][28];
    ele[13][26] != ele[14][29];
    ele[13][26] != ele[15][24];
    ele[13][26] != ele[15][25];
    ele[13][26] != ele[15][26];
    ele[13][26] != ele[15][27];
    ele[13][26] != ele[15][28];
    ele[13][26] != ele[15][29];
    ele[13][26] != ele[16][24];
    ele[13][26] != ele[16][25];
    ele[13][26] != ele[16][26];
    ele[13][26] != ele[16][27];
    ele[13][26] != ele[16][28];
    ele[13][26] != ele[16][29];
    ele[13][26] != ele[17][24];
    ele[13][26] != ele[17][25];
    ele[13][26] != ele[17][26];
    ele[13][26] != ele[17][27];
    ele[13][26] != ele[17][28];
    ele[13][26] != ele[17][29];
    ele[13][26] != ele[18][26];
    ele[13][26] != ele[19][26];
    ele[13][26] != ele[20][26];
    ele[13][26] != ele[21][26];
    ele[13][26] != ele[22][26];
    ele[13][26] != ele[23][26];
    ele[13][26] != ele[24][26];
    ele[13][26] != ele[25][26];
    ele[13][26] != ele[26][26];
    ele[13][26] != ele[27][26];
    ele[13][26] != ele[28][26];
    ele[13][26] != ele[29][26];
    ele[13][26] != ele[30][26];
    ele[13][26] != ele[31][26];
    ele[13][26] != ele[32][26];
    ele[13][26] != ele[33][26];
    ele[13][26] != ele[34][26];
    ele[13][26] != ele[35][26];
    ele[13][27] != ele[13][28];
    ele[13][27] != ele[13][29];
    ele[13][27] != ele[13][30];
    ele[13][27] != ele[13][31];
    ele[13][27] != ele[13][32];
    ele[13][27] != ele[13][33];
    ele[13][27] != ele[13][34];
    ele[13][27] != ele[13][35];
    ele[13][27] != ele[14][24];
    ele[13][27] != ele[14][25];
    ele[13][27] != ele[14][26];
    ele[13][27] != ele[14][27];
    ele[13][27] != ele[14][28];
    ele[13][27] != ele[14][29];
    ele[13][27] != ele[15][24];
    ele[13][27] != ele[15][25];
    ele[13][27] != ele[15][26];
    ele[13][27] != ele[15][27];
    ele[13][27] != ele[15][28];
    ele[13][27] != ele[15][29];
    ele[13][27] != ele[16][24];
    ele[13][27] != ele[16][25];
    ele[13][27] != ele[16][26];
    ele[13][27] != ele[16][27];
    ele[13][27] != ele[16][28];
    ele[13][27] != ele[16][29];
    ele[13][27] != ele[17][24];
    ele[13][27] != ele[17][25];
    ele[13][27] != ele[17][26];
    ele[13][27] != ele[17][27];
    ele[13][27] != ele[17][28];
    ele[13][27] != ele[17][29];
    ele[13][27] != ele[18][27];
    ele[13][27] != ele[19][27];
    ele[13][27] != ele[20][27];
    ele[13][27] != ele[21][27];
    ele[13][27] != ele[22][27];
    ele[13][27] != ele[23][27];
    ele[13][27] != ele[24][27];
    ele[13][27] != ele[25][27];
    ele[13][27] != ele[26][27];
    ele[13][27] != ele[27][27];
    ele[13][27] != ele[28][27];
    ele[13][27] != ele[29][27];
    ele[13][27] != ele[30][27];
    ele[13][27] != ele[31][27];
    ele[13][27] != ele[32][27];
    ele[13][27] != ele[33][27];
    ele[13][27] != ele[34][27];
    ele[13][27] != ele[35][27];
    ele[13][28] != ele[13][29];
    ele[13][28] != ele[13][30];
    ele[13][28] != ele[13][31];
    ele[13][28] != ele[13][32];
    ele[13][28] != ele[13][33];
    ele[13][28] != ele[13][34];
    ele[13][28] != ele[13][35];
    ele[13][28] != ele[14][24];
    ele[13][28] != ele[14][25];
    ele[13][28] != ele[14][26];
    ele[13][28] != ele[14][27];
    ele[13][28] != ele[14][28];
    ele[13][28] != ele[14][29];
    ele[13][28] != ele[15][24];
    ele[13][28] != ele[15][25];
    ele[13][28] != ele[15][26];
    ele[13][28] != ele[15][27];
    ele[13][28] != ele[15][28];
    ele[13][28] != ele[15][29];
    ele[13][28] != ele[16][24];
    ele[13][28] != ele[16][25];
    ele[13][28] != ele[16][26];
    ele[13][28] != ele[16][27];
    ele[13][28] != ele[16][28];
    ele[13][28] != ele[16][29];
    ele[13][28] != ele[17][24];
    ele[13][28] != ele[17][25];
    ele[13][28] != ele[17][26];
    ele[13][28] != ele[17][27];
    ele[13][28] != ele[17][28];
    ele[13][28] != ele[17][29];
    ele[13][28] != ele[18][28];
    ele[13][28] != ele[19][28];
    ele[13][28] != ele[20][28];
    ele[13][28] != ele[21][28];
    ele[13][28] != ele[22][28];
    ele[13][28] != ele[23][28];
    ele[13][28] != ele[24][28];
    ele[13][28] != ele[25][28];
    ele[13][28] != ele[26][28];
    ele[13][28] != ele[27][28];
    ele[13][28] != ele[28][28];
    ele[13][28] != ele[29][28];
    ele[13][28] != ele[30][28];
    ele[13][28] != ele[31][28];
    ele[13][28] != ele[32][28];
    ele[13][28] != ele[33][28];
    ele[13][28] != ele[34][28];
    ele[13][28] != ele[35][28];
    ele[13][29] != ele[13][30];
    ele[13][29] != ele[13][31];
    ele[13][29] != ele[13][32];
    ele[13][29] != ele[13][33];
    ele[13][29] != ele[13][34];
    ele[13][29] != ele[13][35];
    ele[13][29] != ele[14][24];
    ele[13][29] != ele[14][25];
    ele[13][29] != ele[14][26];
    ele[13][29] != ele[14][27];
    ele[13][29] != ele[14][28];
    ele[13][29] != ele[14][29];
    ele[13][29] != ele[15][24];
    ele[13][29] != ele[15][25];
    ele[13][29] != ele[15][26];
    ele[13][29] != ele[15][27];
    ele[13][29] != ele[15][28];
    ele[13][29] != ele[15][29];
    ele[13][29] != ele[16][24];
    ele[13][29] != ele[16][25];
    ele[13][29] != ele[16][26];
    ele[13][29] != ele[16][27];
    ele[13][29] != ele[16][28];
    ele[13][29] != ele[16][29];
    ele[13][29] != ele[17][24];
    ele[13][29] != ele[17][25];
    ele[13][29] != ele[17][26];
    ele[13][29] != ele[17][27];
    ele[13][29] != ele[17][28];
    ele[13][29] != ele[17][29];
    ele[13][29] != ele[18][29];
    ele[13][29] != ele[19][29];
    ele[13][29] != ele[20][29];
    ele[13][29] != ele[21][29];
    ele[13][29] != ele[22][29];
    ele[13][29] != ele[23][29];
    ele[13][29] != ele[24][29];
    ele[13][29] != ele[25][29];
    ele[13][29] != ele[26][29];
    ele[13][29] != ele[27][29];
    ele[13][29] != ele[28][29];
    ele[13][29] != ele[29][29];
    ele[13][29] != ele[30][29];
    ele[13][29] != ele[31][29];
    ele[13][29] != ele[32][29];
    ele[13][29] != ele[33][29];
    ele[13][29] != ele[34][29];
    ele[13][29] != ele[35][29];
    ele[13][3] != ele[13][10];
    ele[13][3] != ele[13][11];
    ele[13][3] != ele[13][12];
    ele[13][3] != ele[13][13];
    ele[13][3] != ele[13][14];
    ele[13][3] != ele[13][15];
    ele[13][3] != ele[13][16];
    ele[13][3] != ele[13][17];
    ele[13][3] != ele[13][18];
    ele[13][3] != ele[13][19];
    ele[13][3] != ele[13][20];
    ele[13][3] != ele[13][21];
    ele[13][3] != ele[13][22];
    ele[13][3] != ele[13][23];
    ele[13][3] != ele[13][24];
    ele[13][3] != ele[13][25];
    ele[13][3] != ele[13][26];
    ele[13][3] != ele[13][27];
    ele[13][3] != ele[13][28];
    ele[13][3] != ele[13][29];
    ele[13][3] != ele[13][30];
    ele[13][3] != ele[13][31];
    ele[13][3] != ele[13][32];
    ele[13][3] != ele[13][33];
    ele[13][3] != ele[13][34];
    ele[13][3] != ele[13][35];
    ele[13][3] != ele[13][4];
    ele[13][3] != ele[13][5];
    ele[13][3] != ele[13][6];
    ele[13][3] != ele[13][7];
    ele[13][3] != ele[13][8];
    ele[13][3] != ele[13][9];
    ele[13][3] != ele[14][0];
    ele[13][3] != ele[14][1];
    ele[13][3] != ele[14][2];
    ele[13][3] != ele[14][3];
    ele[13][3] != ele[14][4];
    ele[13][3] != ele[14][5];
    ele[13][3] != ele[15][0];
    ele[13][3] != ele[15][1];
    ele[13][3] != ele[15][2];
    ele[13][3] != ele[15][3];
    ele[13][3] != ele[15][4];
    ele[13][3] != ele[15][5];
    ele[13][3] != ele[16][0];
    ele[13][3] != ele[16][1];
    ele[13][3] != ele[16][2];
    ele[13][3] != ele[16][3];
    ele[13][3] != ele[16][4];
    ele[13][3] != ele[16][5];
    ele[13][3] != ele[17][0];
    ele[13][3] != ele[17][1];
    ele[13][3] != ele[17][2];
    ele[13][3] != ele[17][3];
    ele[13][3] != ele[17][4];
    ele[13][3] != ele[17][5];
    ele[13][3] != ele[18][3];
    ele[13][3] != ele[19][3];
    ele[13][3] != ele[20][3];
    ele[13][3] != ele[21][3];
    ele[13][3] != ele[22][3];
    ele[13][3] != ele[23][3];
    ele[13][3] != ele[24][3];
    ele[13][3] != ele[25][3];
    ele[13][3] != ele[26][3];
    ele[13][3] != ele[27][3];
    ele[13][3] != ele[28][3];
    ele[13][3] != ele[29][3];
    ele[13][3] != ele[30][3];
    ele[13][3] != ele[31][3];
    ele[13][3] != ele[32][3];
    ele[13][3] != ele[33][3];
    ele[13][3] != ele[34][3];
    ele[13][3] != ele[35][3];
    ele[13][30] != ele[13][31];
    ele[13][30] != ele[13][32];
    ele[13][30] != ele[13][33];
    ele[13][30] != ele[13][34];
    ele[13][30] != ele[13][35];
    ele[13][30] != ele[14][30];
    ele[13][30] != ele[14][31];
    ele[13][30] != ele[14][32];
    ele[13][30] != ele[14][33];
    ele[13][30] != ele[14][34];
    ele[13][30] != ele[14][35];
    ele[13][30] != ele[15][30];
    ele[13][30] != ele[15][31];
    ele[13][30] != ele[15][32];
    ele[13][30] != ele[15][33];
    ele[13][30] != ele[15][34];
    ele[13][30] != ele[15][35];
    ele[13][30] != ele[16][30];
    ele[13][30] != ele[16][31];
    ele[13][30] != ele[16][32];
    ele[13][30] != ele[16][33];
    ele[13][30] != ele[16][34];
    ele[13][30] != ele[16][35];
    ele[13][30] != ele[17][30];
    ele[13][30] != ele[17][31];
    ele[13][30] != ele[17][32];
    ele[13][30] != ele[17][33];
    ele[13][30] != ele[17][34];
    ele[13][30] != ele[17][35];
    ele[13][30] != ele[18][30];
    ele[13][30] != ele[19][30];
    ele[13][30] != ele[20][30];
    ele[13][30] != ele[21][30];
    ele[13][30] != ele[22][30];
    ele[13][30] != ele[23][30];
    ele[13][30] != ele[24][30];
    ele[13][30] != ele[25][30];
    ele[13][30] != ele[26][30];
    ele[13][30] != ele[27][30];
    ele[13][30] != ele[28][30];
    ele[13][30] != ele[29][30];
    ele[13][30] != ele[30][30];
    ele[13][30] != ele[31][30];
    ele[13][30] != ele[32][30];
    ele[13][30] != ele[33][30];
    ele[13][30] != ele[34][30];
    ele[13][30] != ele[35][30];
    ele[13][31] != ele[13][32];
    ele[13][31] != ele[13][33];
    ele[13][31] != ele[13][34];
    ele[13][31] != ele[13][35];
    ele[13][31] != ele[14][30];
    ele[13][31] != ele[14][31];
    ele[13][31] != ele[14][32];
    ele[13][31] != ele[14][33];
    ele[13][31] != ele[14][34];
    ele[13][31] != ele[14][35];
    ele[13][31] != ele[15][30];
    ele[13][31] != ele[15][31];
    ele[13][31] != ele[15][32];
    ele[13][31] != ele[15][33];
    ele[13][31] != ele[15][34];
    ele[13][31] != ele[15][35];
    ele[13][31] != ele[16][30];
    ele[13][31] != ele[16][31];
    ele[13][31] != ele[16][32];
    ele[13][31] != ele[16][33];
    ele[13][31] != ele[16][34];
    ele[13][31] != ele[16][35];
    ele[13][31] != ele[17][30];
    ele[13][31] != ele[17][31];
    ele[13][31] != ele[17][32];
    ele[13][31] != ele[17][33];
    ele[13][31] != ele[17][34];
    ele[13][31] != ele[17][35];
    ele[13][31] != ele[18][31];
    ele[13][31] != ele[19][31];
    ele[13][31] != ele[20][31];
    ele[13][31] != ele[21][31];
    ele[13][31] != ele[22][31];
    ele[13][31] != ele[23][31];
    ele[13][31] != ele[24][31];
    ele[13][31] != ele[25][31];
    ele[13][31] != ele[26][31];
    ele[13][31] != ele[27][31];
    ele[13][31] != ele[28][31];
    ele[13][31] != ele[29][31];
    ele[13][31] != ele[30][31];
    ele[13][31] != ele[31][31];
    ele[13][31] != ele[32][31];
    ele[13][31] != ele[33][31];
    ele[13][31] != ele[34][31];
    ele[13][31] != ele[35][31];
    ele[13][32] != ele[13][33];
    ele[13][32] != ele[13][34];
    ele[13][32] != ele[13][35];
    ele[13][32] != ele[14][30];
    ele[13][32] != ele[14][31];
    ele[13][32] != ele[14][32];
    ele[13][32] != ele[14][33];
    ele[13][32] != ele[14][34];
    ele[13][32] != ele[14][35];
    ele[13][32] != ele[15][30];
    ele[13][32] != ele[15][31];
    ele[13][32] != ele[15][32];
    ele[13][32] != ele[15][33];
    ele[13][32] != ele[15][34];
    ele[13][32] != ele[15][35];
    ele[13][32] != ele[16][30];
    ele[13][32] != ele[16][31];
    ele[13][32] != ele[16][32];
    ele[13][32] != ele[16][33];
    ele[13][32] != ele[16][34];
    ele[13][32] != ele[16][35];
    ele[13][32] != ele[17][30];
    ele[13][32] != ele[17][31];
    ele[13][32] != ele[17][32];
    ele[13][32] != ele[17][33];
    ele[13][32] != ele[17][34];
    ele[13][32] != ele[17][35];
    ele[13][32] != ele[18][32];
    ele[13][32] != ele[19][32];
    ele[13][32] != ele[20][32];
    ele[13][32] != ele[21][32];
    ele[13][32] != ele[22][32];
    ele[13][32] != ele[23][32];
    ele[13][32] != ele[24][32];
    ele[13][32] != ele[25][32];
    ele[13][32] != ele[26][32];
    ele[13][32] != ele[27][32];
    ele[13][32] != ele[28][32];
    ele[13][32] != ele[29][32];
    ele[13][32] != ele[30][32];
    ele[13][32] != ele[31][32];
    ele[13][32] != ele[32][32];
    ele[13][32] != ele[33][32];
    ele[13][32] != ele[34][32];
    ele[13][32] != ele[35][32];
    ele[13][33] != ele[13][34];
    ele[13][33] != ele[13][35];
    ele[13][33] != ele[14][30];
    ele[13][33] != ele[14][31];
    ele[13][33] != ele[14][32];
    ele[13][33] != ele[14][33];
    ele[13][33] != ele[14][34];
    ele[13][33] != ele[14][35];
    ele[13][33] != ele[15][30];
    ele[13][33] != ele[15][31];
    ele[13][33] != ele[15][32];
    ele[13][33] != ele[15][33];
    ele[13][33] != ele[15][34];
    ele[13][33] != ele[15][35];
    ele[13][33] != ele[16][30];
    ele[13][33] != ele[16][31];
    ele[13][33] != ele[16][32];
    ele[13][33] != ele[16][33];
    ele[13][33] != ele[16][34];
    ele[13][33] != ele[16][35];
    ele[13][33] != ele[17][30];
    ele[13][33] != ele[17][31];
    ele[13][33] != ele[17][32];
    ele[13][33] != ele[17][33];
    ele[13][33] != ele[17][34];
    ele[13][33] != ele[17][35];
    ele[13][33] != ele[18][33];
    ele[13][33] != ele[19][33];
    ele[13][33] != ele[20][33];
    ele[13][33] != ele[21][33];
    ele[13][33] != ele[22][33];
    ele[13][33] != ele[23][33];
    ele[13][33] != ele[24][33];
    ele[13][33] != ele[25][33];
    ele[13][33] != ele[26][33];
    ele[13][33] != ele[27][33];
    ele[13][33] != ele[28][33];
    ele[13][33] != ele[29][33];
    ele[13][33] != ele[30][33];
    ele[13][33] != ele[31][33];
    ele[13][33] != ele[32][33];
    ele[13][33] != ele[33][33];
    ele[13][33] != ele[34][33];
    ele[13][33] != ele[35][33];
    ele[13][34] != ele[13][35];
    ele[13][34] != ele[14][30];
    ele[13][34] != ele[14][31];
    ele[13][34] != ele[14][32];
    ele[13][34] != ele[14][33];
    ele[13][34] != ele[14][34];
    ele[13][34] != ele[14][35];
    ele[13][34] != ele[15][30];
    ele[13][34] != ele[15][31];
    ele[13][34] != ele[15][32];
    ele[13][34] != ele[15][33];
    ele[13][34] != ele[15][34];
    ele[13][34] != ele[15][35];
    ele[13][34] != ele[16][30];
    ele[13][34] != ele[16][31];
    ele[13][34] != ele[16][32];
    ele[13][34] != ele[16][33];
    ele[13][34] != ele[16][34];
    ele[13][34] != ele[16][35];
    ele[13][34] != ele[17][30];
    ele[13][34] != ele[17][31];
    ele[13][34] != ele[17][32];
    ele[13][34] != ele[17][33];
    ele[13][34] != ele[17][34];
    ele[13][34] != ele[17][35];
    ele[13][34] != ele[18][34];
    ele[13][34] != ele[19][34];
    ele[13][34] != ele[20][34];
    ele[13][34] != ele[21][34];
    ele[13][34] != ele[22][34];
    ele[13][34] != ele[23][34];
    ele[13][34] != ele[24][34];
    ele[13][34] != ele[25][34];
    ele[13][34] != ele[26][34];
    ele[13][34] != ele[27][34];
    ele[13][34] != ele[28][34];
    ele[13][34] != ele[29][34];
    ele[13][34] != ele[30][34];
    ele[13][34] != ele[31][34];
    ele[13][34] != ele[32][34];
    ele[13][34] != ele[33][34];
    ele[13][34] != ele[34][34];
    ele[13][34] != ele[35][34];
    ele[13][35] != ele[14][30];
    ele[13][35] != ele[14][31];
    ele[13][35] != ele[14][32];
    ele[13][35] != ele[14][33];
    ele[13][35] != ele[14][34];
    ele[13][35] != ele[14][35];
    ele[13][35] != ele[15][30];
    ele[13][35] != ele[15][31];
    ele[13][35] != ele[15][32];
    ele[13][35] != ele[15][33];
    ele[13][35] != ele[15][34];
    ele[13][35] != ele[15][35];
    ele[13][35] != ele[16][30];
    ele[13][35] != ele[16][31];
    ele[13][35] != ele[16][32];
    ele[13][35] != ele[16][33];
    ele[13][35] != ele[16][34];
    ele[13][35] != ele[16][35];
    ele[13][35] != ele[17][30];
    ele[13][35] != ele[17][31];
    ele[13][35] != ele[17][32];
    ele[13][35] != ele[17][33];
    ele[13][35] != ele[17][34];
    ele[13][35] != ele[17][35];
    ele[13][35] != ele[18][35];
    ele[13][35] != ele[19][35];
    ele[13][35] != ele[20][35];
    ele[13][35] != ele[21][35];
    ele[13][35] != ele[22][35];
    ele[13][35] != ele[23][35];
    ele[13][35] != ele[24][35];
    ele[13][35] != ele[25][35];
    ele[13][35] != ele[26][35];
    ele[13][35] != ele[27][35];
    ele[13][35] != ele[28][35];
    ele[13][35] != ele[29][35];
    ele[13][35] != ele[30][35];
    ele[13][35] != ele[31][35];
    ele[13][35] != ele[32][35];
    ele[13][35] != ele[33][35];
    ele[13][35] != ele[34][35];
    ele[13][35] != ele[35][35];
    ele[13][4] != ele[13][10];
    ele[13][4] != ele[13][11];
    ele[13][4] != ele[13][12];
    ele[13][4] != ele[13][13];
    ele[13][4] != ele[13][14];
    ele[13][4] != ele[13][15];
    ele[13][4] != ele[13][16];
    ele[13][4] != ele[13][17];
    ele[13][4] != ele[13][18];
    ele[13][4] != ele[13][19];
    ele[13][4] != ele[13][20];
    ele[13][4] != ele[13][21];
    ele[13][4] != ele[13][22];
    ele[13][4] != ele[13][23];
    ele[13][4] != ele[13][24];
    ele[13][4] != ele[13][25];
    ele[13][4] != ele[13][26];
    ele[13][4] != ele[13][27];
    ele[13][4] != ele[13][28];
    ele[13][4] != ele[13][29];
    ele[13][4] != ele[13][30];
    ele[13][4] != ele[13][31];
    ele[13][4] != ele[13][32];
    ele[13][4] != ele[13][33];
    ele[13][4] != ele[13][34];
    ele[13][4] != ele[13][35];
    ele[13][4] != ele[13][5];
    ele[13][4] != ele[13][6];
    ele[13][4] != ele[13][7];
    ele[13][4] != ele[13][8];
    ele[13][4] != ele[13][9];
    ele[13][4] != ele[14][0];
    ele[13][4] != ele[14][1];
    ele[13][4] != ele[14][2];
    ele[13][4] != ele[14][3];
    ele[13][4] != ele[14][4];
    ele[13][4] != ele[14][5];
    ele[13][4] != ele[15][0];
    ele[13][4] != ele[15][1];
    ele[13][4] != ele[15][2];
    ele[13][4] != ele[15][3];
    ele[13][4] != ele[15][4];
    ele[13][4] != ele[15][5];
    ele[13][4] != ele[16][0];
    ele[13][4] != ele[16][1];
    ele[13][4] != ele[16][2];
    ele[13][4] != ele[16][3];
    ele[13][4] != ele[16][4];
    ele[13][4] != ele[16][5];
    ele[13][4] != ele[17][0];
    ele[13][4] != ele[17][1];
    ele[13][4] != ele[17][2];
    ele[13][4] != ele[17][3];
    ele[13][4] != ele[17][4];
    ele[13][4] != ele[17][5];
    ele[13][4] != ele[18][4];
    ele[13][4] != ele[19][4];
    ele[13][4] != ele[20][4];
    ele[13][4] != ele[21][4];
    ele[13][4] != ele[22][4];
    ele[13][4] != ele[23][4];
    ele[13][4] != ele[24][4];
    ele[13][4] != ele[25][4];
    ele[13][4] != ele[26][4];
    ele[13][4] != ele[27][4];
    ele[13][4] != ele[28][4];
    ele[13][4] != ele[29][4];
    ele[13][4] != ele[30][4];
    ele[13][4] != ele[31][4];
    ele[13][4] != ele[32][4];
    ele[13][4] != ele[33][4];
    ele[13][4] != ele[34][4];
    ele[13][4] != ele[35][4];
    ele[13][5] != ele[13][10];
    ele[13][5] != ele[13][11];
    ele[13][5] != ele[13][12];
    ele[13][5] != ele[13][13];
    ele[13][5] != ele[13][14];
    ele[13][5] != ele[13][15];
    ele[13][5] != ele[13][16];
    ele[13][5] != ele[13][17];
    ele[13][5] != ele[13][18];
    ele[13][5] != ele[13][19];
    ele[13][5] != ele[13][20];
    ele[13][5] != ele[13][21];
    ele[13][5] != ele[13][22];
    ele[13][5] != ele[13][23];
    ele[13][5] != ele[13][24];
    ele[13][5] != ele[13][25];
    ele[13][5] != ele[13][26];
    ele[13][5] != ele[13][27];
    ele[13][5] != ele[13][28];
    ele[13][5] != ele[13][29];
    ele[13][5] != ele[13][30];
    ele[13][5] != ele[13][31];
    ele[13][5] != ele[13][32];
    ele[13][5] != ele[13][33];
    ele[13][5] != ele[13][34];
    ele[13][5] != ele[13][35];
    ele[13][5] != ele[13][6];
    ele[13][5] != ele[13][7];
    ele[13][5] != ele[13][8];
    ele[13][5] != ele[13][9];
    ele[13][5] != ele[14][0];
    ele[13][5] != ele[14][1];
    ele[13][5] != ele[14][2];
    ele[13][5] != ele[14][3];
    ele[13][5] != ele[14][4];
    ele[13][5] != ele[14][5];
    ele[13][5] != ele[15][0];
    ele[13][5] != ele[15][1];
    ele[13][5] != ele[15][2];
    ele[13][5] != ele[15][3];
    ele[13][5] != ele[15][4];
    ele[13][5] != ele[15][5];
    ele[13][5] != ele[16][0];
    ele[13][5] != ele[16][1];
    ele[13][5] != ele[16][2];
    ele[13][5] != ele[16][3];
    ele[13][5] != ele[16][4];
    ele[13][5] != ele[16][5];
    ele[13][5] != ele[17][0];
    ele[13][5] != ele[17][1];
    ele[13][5] != ele[17][2];
    ele[13][5] != ele[17][3];
    ele[13][5] != ele[17][4];
    ele[13][5] != ele[17][5];
    ele[13][5] != ele[18][5];
    ele[13][5] != ele[19][5];
    ele[13][5] != ele[20][5];
    ele[13][5] != ele[21][5];
    ele[13][5] != ele[22][5];
    ele[13][5] != ele[23][5];
    ele[13][5] != ele[24][5];
    ele[13][5] != ele[25][5];
    ele[13][5] != ele[26][5];
    ele[13][5] != ele[27][5];
    ele[13][5] != ele[28][5];
    ele[13][5] != ele[29][5];
    ele[13][5] != ele[30][5];
    ele[13][5] != ele[31][5];
    ele[13][5] != ele[32][5];
    ele[13][5] != ele[33][5];
    ele[13][5] != ele[34][5];
    ele[13][5] != ele[35][5];
    ele[13][6] != ele[13][10];
    ele[13][6] != ele[13][11];
    ele[13][6] != ele[13][12];
    ele[13][6] != ele[13][13];
    ele[13][6] != ele[13][14];
    ele[13][6] != ele[13][15];
    ele[13][6] != ele[13][16];
    ele[13][6] != ele[13][17];
    ele[13][6] != ele[13][18];
    ele[13][6] != ele[13][19];
    ele[13][6] != ele[13][20];
    ele[13][6] != ele[13][21];
    ele[13][6] != ele[13][22];
    ele[13][6] != ele[13][23];
    ele[13][6] != ele[13][24];
    ele[13][6] != ele[13][25];
    ele[13][6] != ele[13][26];
    ele[13][6] != ele[13][27];
    ele[13][6] != ele[13][28];
    ele[13][6] != ele[13][29];
    ele[13][6] != ele[13][30];
    ele[13][6] != ele[13][31];
    ele[13][6] != ele[13][32];
    ele[13][6] != ele[13][33];
    ele[13][6] != ele[13][34];
    ele[13][6] != ele[13][35];
    ele[13][6] != ele[13][7];
    ele[13][6] != ele[13][8];
    ele[13][6] != ele[13][9];
    ele[13][6] != ele[14][10];
    ele[13][6] != ele[14][11];
    ele[13][6] != ele[14][6];
    ele[13][6] != ele[14][7];
    ele[13][6] != ele[14][8];
    ele[13][6] != ele[14][9];
    ele[13][6] != ele[15][10];
    ele[13][6] != ele[15][11];
    ele[13][6] != ele[15][6];
    ele[13][6] != ele[15][7];
    ele[13][6] != ele[15][8];
    ele[13][6] != ele[15][9];
    ele[13][6] != ele[16][10];
    ele[13][6] != ele[16][11];
    ele[13][6] != ele[16][6];
    ele[13][6] != ele[16][7];
    ele[13][6] != ele[16][8];
    ele[13][6] != ele[16][9];
    ele[13][6] != ele[17][10];
    ele[13][6] != ele[17][11];
    ele[13][6] != ele[17][6];
    ele[13][6] != ele[17][7];
    ele[13][6] != ele[17][8];
    ele[13][6] != ele[17][9];
    ele[13][6] != ele[18][6];
    ele[13][6] != ele[19][6];
    ele[13][6] != ele[20][6];
    ele[13][6] != ele[21][6];
    ele[13][6] != ele[22][6];
    ele[13][6] != ele[23][6];
    ele[13][6] != ele[24][6];
    ele[13][6] != ele[25][6];
    ele[13][6] != ele[26][6];
    ele[13][6] != ele[27][6];
    ele[13][6] != ele[28][6];
    ele[13][6] != ele[29][6];
    ele[13][6] != ele[30][6];
    ele[13][6] != ele[31][6];
    ele[13][6] != ele[32][6];
    ele[13][6] != ele[33][6];
    ele[13][6] != ele[34][6];
    ele[13][6] != ele[35][6];
    ele[13][7] != ele[13][10];
    ele[13][7] != ele[13][11];
    ele[13][7] != ele[13][12];
    ele[13][7] != ele[13][13];
    ele[13][7] != ele[13][14];
    ele[13][7] != ele[13][15];
    ele[13][7] != ele[13][16];
    ele[13][7] != ele[13][17];
    ele[13][7] != ele[13][18];
    ele[13][7] != ele[13][19];
    ele[13][7] != ele[13][20];
    ele[13][7] != ele[13][21];
    ele[13][7] != ele[13][22];
    ele[13][7] != ele[13][23];
    ele[13][7] != ele[13][24];
    ele[13][7] != ele[13][25];
    ele[13][7] != ele[13][26];
    ele[13][7] != ele[13][27];
    ele[13][7] != ele[13][28];
    ele[13][7] != ele[13][29];
    ele[13][7] != ele[13][30];
    ele[13][7] != ele[13][31];
    ele[13][7] != ele[13][32];
    ele[13][7] != ele[13][33];
    ele[13][7] != ele[13][34];
    ele[13][7] != ele[13][35];
    ele[13][7] != ele[13][8];
    ele[13][7] != ele[13][9];
    ele[13][7] != ele[14][10];
    ele[13][7] != ele[14][11];
    ele[13][7] != ele[14][6];
    ele[13][7] != ele[14][7];
    ele[13][7] != ele[14][8];
    ele[13][7] != ele[14][9];
    ele[13][7] != ele[15][10];
    ele[13][7] != ele[15][11];
    ele[13][7] != ele[15][6];
    ele[13][7] != ele[15][7];
    ele[13][7] != ele[15][8];
    ele[13][7] != ele[15][9];
    ele[13][7] != ele[16][10];
    ele[13][7] != ele[16][11];
    ele[13][7] != ele[16][6];
    ele[13][7] != ele[16][7];
    ele[13][7] != ele[16][8];
    ele[13][7] != ele[16][9];
    ele[13][7] != ele[17][10];
    ele[13][7] != ele[17][11];
    ele[13][7] != ele[17][6];
    ele[13][7] != ele[17][7];
    ele[13][7] != ele[17][8];
    ele[13][7] != ele[17][9];
    ele[13][7] != ele[18][7];
    ele[13][7] != ele[19][7];
    ele[13][7] != ele[20][7];
    ele[13][7] != ele[21][7];
    ele[13][7] != ele[22][7];
    ele[13][7] != ele[23][7];
    ele[13][7] != ele[24][7];
    ele[13][7] != ele[25][7];
    ele[13][7] != ele[26][7];
    ele[13][7] != ele[27][7];
    ele[13][7] != ele[28][7];
    ele[13][7] != ele[29][7];
    ele[13][7] != ele[30][7];
    ele[13][7] != ele[31][7];
    ele[13][7] != ele[32][7];
    ele[13][7] != ele[33][7];
    ele[13][7] != ele[34][7];
    ele[13][7] != ele[35][7];
    ele[13][8] != ele[13][10];
    ele[13][8] != ele[13][11];
    ele[13][8] != ele[13][12];
    ele[13][8] != ele[13][13];
    ele[13][8] != ele[13][14];
    ele[13][8] != ele[13][15];
    ele[13][8] != ele[13][16];
    ele[13][8] != ele[13][17];
    ele[13][8] != ele[13][18];
    ele[13][8] != ele[13][19];
    ele[13][8] != ele[13][20];
    ele[13][8] != ele[13][21];
    ele[13][8] != ele[13][22];
    ele[13][8] != ele[13][23];
    ele[13][8] != ele[13][24];
    ele[13][8] != ele[13][25];
    ele[13][8] != ele[13][26];
    ele[13][8] != ele[13][27];
    ele[13][8] != ele[13][28];
    ele[13][8] != ele[13][29];
    ele[13][8] != ele[13][30];
    ele[13][8] != ele[13][31];
    ele[13][8] != ele[13][32];
    ele[13][8] != ele[13][33];
    ele[13][8] != ele[13][34];
    ele[13][8] != ele[13][35];
    ele[13][8] != ele[13][9];
    ele[13][8] != ele[14][10];
    ele[13][8] != ele[14][11];
    ele[13][8] != ele[14][6];
    ele[13][8] != ele[14][7];
    ele[13][8] != ele[14][8];
    ele[13][8] != ele[14][9];
    ele[13][8] != ele[15][10];
    ele[13][8] != ele[15][11];
    ele[13][8] != ele[15][6];
    ele[13][8] != ele[15][7];
    ele[13][8] != ele[15][8];
    ele[13][8] != ele[15][9];
    ele[13][8] != ele[16][10];
    ele[13][8] != ele[16][11];
    ele[13][8] != ele[16][6];
    ele[13][8] != ele[16][7];
    ele[13][8] != ele[16][8];
    ele[13][8] != ele[16][9];
    ele[13][8] != ele[17][10];
    ele[13][8] != ele[17][11];
    ele[13][8] != ele[17][6];
    ele[13][8] != ele[17][7];
    ele[13][8] != ele[17][8];
    ele[13][8] != ele[17][9];
    ele[13][8] != ele[18][8];
    ele[13][8] != ele[19][8];
    ele[13][8] != ele[20][8];
    ele[13][8] != ele[21][8];
    ele[13][8] != ele[22][8];
    ele[13][8] != ele[23][8];
    ele[13][8] != ele[24][8];
    ele[13][8] != ele[25][8];
    ele[13][8] != ele[26][8];
    ele[13][8] != ele[27][8];
    ele[13][8] != ele[28][8];
    ele[13][8] != ele[29][8];
    ele[13][8] != ele[30][8];
    ele[13][8] != ele[31][8];
    ele[13][8] != ele[32][8];
    ele[13][8] != ele[33][8];
    ele[13][8] != ele[34][8];
    ele[13][8] != ele[35][8];
    ele[13][9] != ele[13][10];
    ele[13][9] != ele[13][11];
    ele[13][9] != ele[13][12];
    ele[13][9] != ele[13][13];
    ele[13][9] != ele[13][14];
    ele[13][9] != ele[13][15];
    ele[13][9] != ele[13][16];
    ele[13][9] != ele[13][17];
    ele[13][9] != ele[13][18];
    ele[13][9] != ele[13][19];
    ele[13][9] != ele[13][20];
    ele[13][9] != ele[13][21];
    ele[13][9] != ele[13][22];
    ele[13][9] != ele[13][23];
    ele[13][9] != ele[13][24];
    ele[13][9] != ele[13][25];
    ele[13][9] != ele[13][26];
    ele[13][9] != ele[13][27];
    ele[13][9] != ele[13][28];
    ele[13][9] != ele[13][29];
    ele[13][9] != ele[13][30];
    ele[13][9] != ele[13][31];
    ele[13][9] != ele[13][32];
    ele[13][9] != ele[13][33];
    ele[13][9] != ele[13][34];
    ele[13][9] != ele[13][35];
    ele[13][9] != ele[14][10];
    ele[13][9] != ele[14][11];
    ele[13][9] != ele[14][6];
    ele[13][9] != ele[14][7];
    ele[13][9] != ele[14][8];
    ele[13][9] != ele[14][9];
    ele[13][9] != ele[15][10];
    ele[13][9] != ele[15][11];
    ele[13][9] != ele[15][6];
    ele[13][9] != ele[15][7];
    ele[13][9] != ele[15][8];
    ele[13][9] != ele[15][9];
    ele[13][9] != ele[16][10];
    ele[13][9] != ele[16][11];
    ele[13][9] != ele[16][6];
    ele[13][9] != ele[16][7];
    ele[13][9] != ele[16][8];
    ele[13][9] != ele[16][9];
    ele[13][9] != ele[17][10];
    ele[13][9] != ele[17][11];
    ele[13][9] != ele[17][6];
    ele[13][9] != ele[17][7];
    ele[13][9] != ele[17][8];
    ele[13][9] != ele[17][9];
    ele[13][9] != ele[18][9];
    ele[13][9] != ele[19][9];
    ele[13][9] != ele[20][9];
    ele[13][9] != ele[21][9];
    ele[13][9] != ele[22][9];
    ele[13][9] != ele[23][9];
    ele[13][9] != ele[24][9];
    ele[13][9] != ele[25][9];
    ele[13][9] != ele[26][9];
    ele[13][9] != ele[27][9];
    ele[13][9] != ele[28][9];
    ele[13][9] != ele[29][9];
    ele[13][9] != ele[30][9];
    ele[13][9] != ele[31][9];
    ele[13][9] != ele[32][9];
    ele[13][9] != ele[33][9];
    ele[13][9] != ele[34][9];
    ele[13][9] != ele[35][9];
    ele[14][0] != ele[14][1];
    ele[14][0] != ele[14][10];
    ele[14][0] != ele[14][11];
    ele[14][0] != ele[14][12];
    ele[14][0] != ele[14][13];
    ele[14][0] != ele[14][14];
    ele[14][0] != ele[14][15];
    ele[14][0] != ele[14][16];
    ele[14][0] != ele[14][17];
    ele[14][0] != ele[14][18];
    ele[14][0] != ele[14][19];
    ele[14][0] != ele[14][2];
    ele[14][0] != ele[14][20];
    ele[14][0] != ele[14][21];
    ele[14][0] != ele[14][22];
    ele[14][0] != ele[14][23];
    ele[14][0] != ele[14][24];
    ele[14][0] != ele[14][25];
    ele[14][0] != ele[14][26];
    ele[14][0] != ele[14][27];
    ele[14][0] != ele[14][28];
    ele[14][0] != ele[14][29];
    ele[14][0] != ele[14][3];
    ele[14][0] != ele[14][30];
    ele[14][0] != ele[14][31];
    ele[14][0] != ele[14][32];
    ele[14][0] != ele[14][33];
    ele[14][0] != ele[14][34];
    ele[14][0] != ele[14][35];
    ele[14][0] != ele[14][4];
    ele[14][0] != ele[14][5];
    ele[14][0] != ele[14][6];
    ele[14][0] != ele[14][7];
    ele[14][0] != ele[14][8];
    ele[14][0] != ele[14][9];
    ele[14][0] != ele[15][0];
    ele[14][0] != ele[15][1];
    ele[14][0] != ele[15][2];
    ele[14][0] != ele[15][3];
    ele[14][0] != ele[15][4];
    ele[14][0] != ele[15][5];
    ele[14][0] != ele[16][0];
    ele[14][0] != ele[16][1];
    ele[14][0] != ele[16][2];
    ele[14][0] != ele[16][3];
    ele[14][0] != ele[16][4];
    ele[14][0] != ele[16][5];
    ele[14][0] != ele[17][0];
    ele[14][0] != ele[17][1];
    ele[14][0] != ele[17][2];
    ele[14][0] != ele[17][3];
    ele[14][0] != ele[17][4];
    ele[14][0] != ele[17][5];
    ele[14][0] != ele[18][0];
    ele[14][0] != ele[19][0];
    ele[14][0] != ele[20][0];
    ele[14][0] != ele[21][0];
    ele[14][0] != ele[22][0];
    ele[14][0] != ele[23][0];
    ele[14][0] != ele[24][0];
    ele[14][0] != ele[25][0];
    ele[14][0] != ele[26][0];
    ele[14][0] != ele[27][0];
    ele[14][0] != ele[28][0];
    ele[14][0] != ele[29][0];
    ele[14][0] != ele[30][0];
    ele[14][0] != ele[31][0];
    ele[14][0] != ele[32][0];
    ele[14][0] != ele[33][0];
    ele[14][0] != ele[34][0];
    ele[14][0] != ele[35][0];
    ele[14][1] != ele[14][10];
    ele[14][1] != ele[14][11];
    ele[14][1] != ele[14][12];
    ele[14][1] != ele[14][13];
    ele[14][1] != ele[14][14];
    ele[14][1] != ele[14][15];
    ele[14][1] != ele[14][16];
    ele[14][1] != ele[14][17];
    ele[14][1] != ele[14][18];
    ele[14][1] != ele[14][19];
    ele[14][1] != ele[14][2];
    ele[14][1] != ele[14][20];
    ele[14][1] != ele[14][21];
    ele[14][1] != ele[14][22];
    ele[14][1] != ele[14][23];
    ele[14][1] != ele[14][24];
    ele[14][1] != ele[14][25];
    ele[14][1] != ele[14][26];
    ele[14][1] != ele[14][27];
    ele[14][1] != ele[14][28];
    ele[14][1] != ele[14][29];
    ele[14][1] != ele[14][3];
    ele[14][1] != ele[14][30];
    ele[14][1] != ele[14][31];
    ele[14][1] != ele[14][32];
    ele[14][1] != ele[14][33];
    ele[14][1] != ele[14][34];
    ele[14][1] != ele[14][35];
    ele[14][1] != ele[14][4];
    ele[14][1] != ele[14][5];
    ele[14][1] != ele[14][6];
    ele[14][1] != ele[14][7];
    ele[14][1] != ele[14][8];
    ele[14][1] != ele[14][9];
    ele[14][1] != ele[15][0];
    ele[14][1] != ele[15][1];
    ele[14][1] != ele[15][2];
    ele[14][1] != ele[15][3];
    ele[14][1] != ele[15][4];
    ele[14][1] != ele[15][5];
    ele[14][1] != ele[16][0];
    ele[14][1] != ele[16][1];
    ele[14][1] != ele[16][2];
    ele[14][1] != ele[16][3];
    ele[14][1] != ele[16][4];
    ele[14][1] != ele[16][5];
    ele[14][1] != ele[17][0];
    ele[14][1] != ele[17][1];
    ele[14][1] != ele[17][2];
    ele[14][1] != ele[17][3];
    ele[14][1] != ele[17][4];
    ele[14][1] != ele[17][5];
    ele[14][1] != ele[18][1];
    ele[14][1] != ele[19][1];
    ele[14][1] != ele[20][1];
    ele[14][1] != ele[21][1];
    ele[14][1] != ele[22][1];
    ele[14][1] != ele[23][1];
    ele[14][1] != ele[24][1];
    ele[14][1] != ele[25][1];
    ele[14][1] != ele[26][1];
    ele[14][1] != ele[27][1];
    ele[14][1] != ele[28][1];
    ele[14][1] != ele[29][1];
    ele[14][1] != ele[30][1];
    ele[14][1] != ele[31][1];
    ele[14][1] != ele[32][1];
    ele[14][1] != ele[33][1];
    ele[14][1] != ele[34][1];
    ele[14][1] != ele[35][1];
    ele[14][10] != ele[14][11];
    ele[14][10] != ele[14][12];
    ele[14][10] != ele[14][13];
    ele[14][10] != ele[14][14];
    ele[14][10] != ele[14][15];
    ele[14][10] != ele[14][16];
    ele[14][10] != ele[14][17];
    ele[14][10] != ele[14][18];
    ele[14][10] != ele[14][19];
    ele[14][10] != ele[14][20];
    ele[14][10] != ele[14][21];
    ele[14][10] != ele[14][22];
    ele[14][10] != ele[14][23];
    ele[14][10] != ele[14][24];
    ele[14][10] != ele[14][25];
    ele[14][10] != ele[14][26];
    ele[14][10] != ele[14][27];
    ele[14][10] != ele[14][28];
    ele[14][10] != ele[14][29];
    ele[14][10] != ele[14][30];
    ele[14][10] != ele[14][31];
    ele[14][10] != ele[14][32];
    ele[14][10] != ele[14][33];
    ele[14][10] != ele[14][34];
    ele[14][10] != ele[14][35];
    ele[14][10] != ele[15][10];
    ele[14][10] != ele[15][11];
    ele[14][10] != ele[15][6];
    ele[14][10] != ele[15][7];
    ele[14][10] != ele[15][8];
    ele[14][10] != ele[15][9];
    ele[14][10] != ele[16][10];
    ele[14][10] != ele[16][11];
    ele[14][10] != ele[16][6];
    ele[14][10] != ele[16][7];
    ele[14][10] != ele[16][8];
    ele[14][10] != ele[16][9];
    ele[14][10] != ele[17][10];
    ele[14][10] != ele[17][11];
    ele[14][10] != ele[17][6];
    ele[14][10] != ele[17][7];
    ele[14][10] != ele[17][8];
    ele[14][10] != ele[17][9];
    ele[14][10] != ele[18][10];
    ele[14][10] != ele[19][10];
    ele[14][10] != ele[20][10];
    ele[14][10] != ele[21][10];
    ele[14][10] != ele[22][10];
    ele[14][10] != ele[23][10];
    ele[14][10] != ele[24][10];
    ele[14][10] != ele[25][10];
    ele[14][10] != ele[26][10];
    ele[14][10] != ele[27][10];
    ele[14][10] != ele[28][10];
    ele[14][10] != ele[29][10];
    ele[14][10] != ele[30][10];
    ele[14][10] != ele[31][10];
    ele[14][10] != ele[32][10];
    ele[14][10] != ele[33][10];
    ele[14][10] != ele[34][10];
    ele[14][10] != ele[35][10];
    ele[14][11] != ele[14][12];
    ele[14][11] != ele[14][13];
    ele[14][11] != ele[14][14];
    ele[14][11] != ele[14][15];
    ele[14][11] != ele[14][16];
    ele[14][11] != ele[14][17];
    ele[14][11] != ele[14][18];
    ele[14][11] != ele[14][19];
    ele[14][11] != ele[14][20];
    ele[14][11] != ele[14][21];
    ele[14][11] != ele[14][22];
    ele[14][11] != ele[14][23];
    ele[14][11] != ele[14][24];
    ele[14][11] != ele[14][25];
    ele[14][11] != ele[14][26];
    ele[14][11] != ele[14][27];
    ele[14][11] != ele[14][28];
    ele[14][11] != ele[14][29];
    ele[14][11] != ele[14][30];
    ele[14][11] != ele[14][31];
    ele[14][11] != ele[14][32];
    ele[14][11] != ele[14][33];
    ele[14][11] != ele[14][34];
    ele[14][11] != ele[14][35];
    ele[14][11] != ele[15][10];
    ele[14][11] != ele[15][11];
    ele[14][11] != ele[15][6];
    ele[14][11] != ele[15][7];
    ele[14][11] != ele[15][8];
    ele[14][11] != ele[15][9];
    ele[14][11] != ele[16][10];
    ele[14][11] != ele[16][11];
    ele[14][11] != ele[16][6];
    ele[14][11] != ele[16][7];
    ele[14][11] != ele[16][8];
    ele[14][11] != ele[16][9];
    ele[14][11] != ele[17][10];
    ele[14][11] != ele[17][11];
    ele[14][11] != ele[17][6];
    ele[14][11] != ele[17][7];
    ele[14][11] != ele[17][8];
    ele[14][11] != ele[17][9];
    ele[14][11] != ele[18][11];
    ele[14][11] != ele[19][11];
    ele[14][11] != ele[20][11];
    ele[14][11] != ele[21][11];
    ele[14][11] != ele[22][11];
    ele[14][11] != ele[23][11];
    ele[14][11] != ele[24][11];
    ele[14][11] != ele[25][11];
    ele[14][11] != ele[26][11];
    ele[14][11] != ele[27][11];
    ele[14][11] != ele[28][11];
    ele[14][11] != ele[29][11];
    ele[14][11] != ele[30][11];
    ele[14][11] != ele[31][11];
    ele[14][11] != ele[32][11];
    ele[14][11] != ele[33][11];
    ele[14][11] != ele[34][11];
    ele[14][11] != ele[35][11];
    ele[14][12] != ele[14][13];
    ele[14][12] != ele[14][14];
    ele[14][12] != ele[14][15];
    ele[14][12] != ele[14][16];
    ele[14][12] != ele[14][17];
    ele[14][12] != ele[14][18];
    ele[14][12] != ele[14][19];
    ele[14][12] != ele[14][20];
    ele[14][12] != ele[14][21];
    ele[14][12] != ele[14][22];
    ele[14][12] != ele[14][23];
    ele[14][12] != ele[14][24];
    ele[14][12] != ele[14][25];
    ele[14][12] != ele[14][26];
    ele[14][12] != ele[14][27];
    ele[14][12] != ele[14][28];
    ele[14][12] != ele[14][29];
    ele[14][12] != ele[14][30];
    ele[14][12] != ele[14][31];
    ele[14][12] != ele[14][32];
    ele[14][12] != ele[14][33];
    ele[14][12] != ele[14][34];
    ele[14][12] != ele[14][35];
    ele[14][12] != ele[15][12];
    ele[14][12] != ele[15][13];
    ele[14][12] != ele[15][14];
    ele[14][12] != ele[15][15];
    ele[14][12] != ele[15][16];
    ele[14][12] != ele[15][17];
    ele[14][12] != ele[16][12];
    ele[14][12] != ele[16][13];
    ele[14][12] != ele[16][14];
    ele[14][12] != ele[16][15];
    ele[14][12] != ele[16][16];
    ele[14][12] != ele[16][17];
    ele[14][12] != ele[17][12];
    ele[14][12] != ele[17][13];
    ele[14][12] != ele[17][14];
    ele[14][12] != ele[17][15];
    ele[14][12] != ele[17][16];
    ele[14][12] != ele[17][17];
    ele[14][12] != ele[18][12];
    ele[14][12] != ele[19][12];
    ele[14][12] != ele[20][12];
    ele[14][12] != ele[21][12];
    ele[14][12] != ele[22][12];
    ele[14][12] != ele[23][12];
    ele[14][12] != ele[24][12];
    ele[14][12] != ele[25][12];
    ele[14][12] != ele[26][12];
    ele[14][12] != ele[27][12];
    ele[14][12] != ele[28][12];
    ele[14][12] != ele[29][12];
    ele[14][12] != ele[30][12];
    ele[14][12] != ele[31][12];
    ele[14][12] != ele[32][12];
    ele[14][12] != ele[33][12];
    ele[14][12] != ele[34][12];
    ele[14][12] != ele[35][12];
    ele[14][13] != ele[14][14];
    ele[14][13] != ele[14][15];
    ele[14][13] != ele[14][16];
    ele[14][13] != ele[14][17];
    ele[14][13] != ele[14][18];
    ele[14][13] != ele[14][19];
    ele[14][13] != ele[14][20];
    ele[14][13] != ele[14][21];
    ele[14][13] != ele[14][22];
    ele[14][13] != ele[14][23];
    ele[14][13] != ele[14][24];
    ele[14][13] != ele[14][25];
    ele[14][13] != ele[14][26];
    ele[14][13] != ele[14][27];
    ele[14][13] != ele[14][28];
    ele[14][13] != ele[14][29];
    ele[14][13] != ele[14][30];
    ele[14][13] != ele[14][31];
    ele[14][13] != ele[14][32];
    ele[14][13] != ele[14][33];
    ele[14][13] != ele[14][34];
    ele[14][13] != ele[14][35];
    ele[14][13] != ele[15][12];
    ele[14][13] != ele[15][13];
    ele[14][13] != ele[15][14];
    ele[14][13] != ele[15][15];
    ele[14][13] != ele[15][16];
    ele[14][13] != ele[15][17];
    ele[14][13] != ele[16][12];
    ele[14][13] != ele[16][13];
    ele[14][13] != ele[16][14];
    ele[14][13] != ele[16][15];
    ele[14][13] != ele[16][16];
    ele[14][13] != ele[16][17];
    ele[14][13] != ele[17][12];
    ele[14][13] != ele[17][13];
    ele[14][13] != ele[17][14];
    ele[14][13] != ele[17][15];
    ele[14][13] != ele[17][16];
    ele[14][13] != ele[17][17];
    ele[14][13] != ele[18][13];
    ele[14][13] != ele[19][13];
    ele[14][13] != ele[20][13];
    ele[14][13] != ele[21][13];
    ele[14][13] != ele[22][13];
    ele[14][13] != ele[23][13];
    ele[14][13] != ele[24][13];
    ele[14][13] != ele[25][13];
    ele[14][13] != ele[26][13];
    ele[14][13] != ele[27][13];
    ele[14][13] != ele[28][13];
    ele[14][13] != ele[29][13];
    ele[14][13] != ele[30][13];
    ele[14][13] != ele[31][13];
    ele[14][13] != ele[32][13];
    ele[14][13] != ele[33][13];
    ele[14][13] != ele[34][13];
    ele[14][13] != ele[35][13];
    ele[14][14] != ele[14][15];
    ele[14][14] != ele[14][16];
    ele[14][14] != ele[14][17];
    ele[14][14] != ele[14][18];
    ele[14][14] != ele[14][19];
    ele[14][14] != ele[14][20];
    ele[14][14] != ele[14][21];
    ele[14][14] != ele[14][22];
    ele[14][14] != ele[14][23];
    ele[14][14] != ele[14][24];
    ele[14][14] != ele[14][25];
    ele[14][14] != ele[14][26];
    ele[14][14] != ele[14][27];
    ele[14][14] != ele[14][28];
    ele[14][14] != ele[14][29];
    ele[14][14] != ele[14][30];
    ele[14][14] != ele[14][31];
    ele[14][14] != ele[14][32];
    ele[14][14] != ele[14][33];
    ele[14][14] != ele[14][34];
    ele[14][14] != ele[14][35];
    ele[14][14] != ele[15][12];
    ele[14][14] != ele[15][13];
    ele[14][14] != ele[15][14];
    ele[14][14] != ele[15][15];
    ele[14][14] != ele[15][16];
    ele[14][14] != ele[15][17];
    ele[14][14] != ele[16][12];
    ele[14][14] != ele[16][13];
    ele[14][14] != ele[16][14];
    ele[14][14] != ele[16][15];
    ele[14][14] != ele[16][16];
    ele[14][14] != ele[16][17];
    ele[14][14] != ele[17][12];
    ele[14][14] != ele[17][13];
    ele[14][14] != ele[17][14];
    ele[14][14] != ele[17][15];
    ele[14][14] != ele[17][16];
    ele[14][14] != ele[17][17];
    ele[14][14] != ele[18][14];
    ele[14][14] != ele[19][14];
    ele[14][14] != ele[20][14];
    ele[14][14] != ele[21][14];
    ele[14][14] != ele[22][14];
    ele[14][14] != ele[23][14];
    ele[14][14] != ele[24][14];
    ele[14][14] != ele[25][14];
    ele[14][14] != ele[26][14];
    ele[14][14] != ele[27][14];
    ele[14][14] != ele[28][14];
    ele[14][14] != ele[29][14];
    ele[14][14] != ele[30][14];
    ele[14][14] != ele[31][14];
    ele[14][14] != ele[32][14];
    ele[14][14] != ele[33][14];
    ele[14][14] != ele[34][14];
    ele[14][14] != ele[35][14];
    ele[14][15] != ele[14][16];
    ele[14][15] != ele[14][17];
    ele[14][15] != ele[14][18];
    ele[14][15] != ele[14][19];
    ele[14][15] != ele[14][20];
    ele[14][15] != ele[14][21];
    ele[14][15] != ele[14][22];
    ele[14][15] != ele[14][23];
    ele[14][15] != ele[14][24];
    ele[14][15] != ele[14][25];
    ele[14][15] != ele[14][26];
    ele[14][15] != ele[14][27];
    ele[14][15] != ele[14][28];
    ele[14][15] != ele[14][29];
    ele[14][15] != ele[14][30];
    ele[14][15] != ele[14][31];
    ele[14][15] != ele[14][32];
    ele[14][15] != ele[14][33];
    ele[14][15] != ele[14][34];
    ele[14][15] != ele[14][35];
    ele[14][15] != ele[15][12];
    ele[14][15] != ele[15][13];
    ele[14][15] != ele[15][14];
    ele[14][15] != ele[15][15];
    ele[14][15] != ele[15][16];
    ele[14][15] != ele[15][17];
    ele[14][15] != ele[16][12];
    ele[14][15] != ele[16][13];
    ele[14][15] != ele[16][14];
    ele[14][15] != ele[16][15];
    ele[14][15] != ele[16][16];
    ele[14][15] != ele[16][17];
    ele[14][15] != ele[17][12];
    ele[14][15] != ele[17][13];
    ele[14][15] != ele[17][14];
    ele[14][15] != ele[17][15];
    ele[14][15] != ele[17][16];
    ele[14][15] != ele[17][17];
    ele[14][15] != ele[18][15];
    ele[14][15] != ele[19][15];
    ele[14][15] != ele[20][15];
    ele[14][15] != ele[21][15];
    ele[14][15] != ele[22][15];
    ele[14][15] != ele[23][15];
    ele[14][15] != ele[24][15];
    ele[14][15] != ele[25][15];
    ele[14][15] != ele[26][15];
    ele[14][15] != ele[27][15];
    ele[14][15] != ele[28][15];
    ele[14][15] != ele[29][15];
    ele[14][15] != ele[30][15];
    ele[14][15] != ele[31][15];
    ele[14][15] != ele[32][15];
    ele[14][15] != ele[33][15];
    ele[14][15] != ele[34][15];
    ele[14][15] != ele[35][15];
    ele[14][16] != ele[14][17];
    ele[14][16] != ele[14][18];
    ele[14][16] != ele[14][19];
    ele[14][16] != ele[14][20];
    ele[14][16] != ele[14][21];
    ele[14][16] != ele[14][22];
    ele[14][16] != ele[14][23];
    ele[14][16] != ele[14][24];
    ele[14][16] != ele[14][25];
    ele[14][16] != ele[14][26];
    ele[14][16] != ele[14][27];
    ele[14][16] != ele[14][28];
    ele[14][16] != ele[14][29];
    ele[14][16] != ele[14][30];
    ele[14][16] != ele[14][31];
    ele[14][16] != ele[14][32];
    ele[14][16] != ele[14][33];
    ele[14][16] != ele[14][34];
    ele[14][16] != ele[14][35];
    ele[14][16] != ele[15][12];
    ele[14][16] != ele[15][13];
    ele[14][16] != ele[15][14];
    ele[14][16] != ele[15][15];
    ele[14][16] != ele[15][16];
    ele[14][16] != ele[15][17];
    ele[14][16] != ele[16][12];
    ele[14][16] != ele[16][13];
    ele[14][16] != ele[16][14];
    ele[14][16] != ele[16][15];
    ele[14][16] != ele[16][16];
    ele[14][16] != ele[16][17];
    ele[14][16] != ele[17][12];
    ele[14][16] != ele[17][13];
    ele[14][16] != ele[17][14];
    ele[14][16] != ele[17][15];
    ele[14][16] != ele[17][16];
    ele[14][16] != ele[17][17];
    ele[14][16] != ele[18][16];
    ele[14][16] != ele[19][16];
    ele[14][16] != ele[20][16];
    ele[14][16] != ele[21][16];
    ele[14][16] != ele[22][16];
    ele[14][16] != ele[23][16];
    ele[14][16] != ele[24][16];
    ele[14][16] != ele[25][16];
    ele[14][16] != ele[26][16];
    ele[14][16] != ele[27][16];
    ele[14][16] != ele[28][16];
    ele[14][16] != ele[29][16];
    ele[14][16] != ele[30][16];
    ele[14][16] != ele[31][16];
    ele[14][16] != ele[32][16];
    ele[14][16] != ele[33][16];
    ele[14][16] != ele[34][16];
    ele[14][16] != ele[35][16];
    ele[14][17] != ele[14][18];
    ele[14][17] != ele[14][19];
    ele[14][17] != ele[14][20];
    ele[14][17] != ele[14][21];
    ele[14][17] != ele[14][22];
    ele[14][17] != ele[14][23];
    ele[14][17] != ele[14][24];
    ele[14][17] != ele[14][25];
    ele[14][17] != ele[14][26];
    ele[14][17] != ele[14][27];
    ele[14][17] != ele[14][28];
    ele[14][17] != ele[14][29];
    ele[14][17] != ele[14][30];
    ele[14][17] != ele[14][31];
    ele[14][17] != ele[14][32];
    ele[14][17] != ele[14][33];
    ele[14][17] != ele[14][34];
    ele[14][17] != ele[14][35];
    ele[14][17] != ele[15][12];
    ele[14][17] != ele[15][13];
    ele[14][17] != ele[15][14];
    ele[14][17] != ele[15][15];
    ele[14][17] != ele[15][16];
    ele[14][17] != ele[15][17];
    ele[14][17] != ele[16][12];
    ele[14][17] != ele[16][13];
    ele[14][17] != ele[16][14];
    ele[14][17] != ele[16][15];
    ele[14][17] != ele[16][16];
    ele[14][17] != ele[16][17];
    ele[14][17] != ele[17][12];
    ele[14][17] != ele[17][13];
    ele[14][17] != ele[17][14];
    ele[14][17] != ele[17][15];
    ele[14][17] != ele[17][16];
    ele[14][17] != ele[17][17];
    ele[14][17] != ele[18][17];
    ele[14][17] != ele[19][17];
    ele[14][17] != ele[20][17];
    ele[14][17] != ele[21][17];
    ele[14][17] != ele[22][17];
    ele[14][17] != ele[23][17];
    ele[14][17] != ele[24][17];
    ele[14][17] != ele[25][17];
    ele[14][17] != ele[26][17];
    ele[14][17] != ele[27][17];
    ele[14][17] != ele[28][17];
    ele[14][17] != ele[29][17];
    ele[14][17] != ele[30][17];
    ele[14][17] != ele[31][17];
    ele[14][17] != ele[32][17];
    ele[14][17] != ele[33][17];
    ele[14][17] != ele[34][17];
    ele[14][17] != ele[35][17];
    ele[14][18] != ele[14][19];
    ele[14][18] != ele[14][20];
    ele[14][18] != ele[14][21];
    ele[14][18] != ele[14][22];
    ele[14][18] != ele[14][23];
    ele[14][18] != ele[14][24];
    ele[14][18] != ele[14][25];
    ele[14][18] != ele[14][26];
    ele[14][18] != ele[14][27];
    ele[14][18] != ele[14][28];
    ele[14][18] != ele[14][29];
    ele[14][18] != ele[14][30];
    ele[14][18] != ele[14][31];
    ele[14][18] != ele[14][32];
    ele[14][18] != ele[14][33];
    ele[14][18] != ele[14][34];
    ele[14][18] != ele[14][35];
    ele[14][18] != ele[15][18];
    ele[14][18] != ele[15][19];
    ele[14][18] != ele[15][20];
    ele[14][18] != ele[15][21];
    ele[14][18] != ele[15][22];
    ele[14][18] != ele[15][23];
    ele[14][18] != ele[16][18];
    ele[14][18] != ele[16][19];
    ele[14][18] != ele[16][20];
    ele[14][18] != ele[16][21];
    ele[14][18] != ele[16][22];
    ele[14][18] != ele[16][23];
    ele[14][18] != ele[17][18];
    ele[14][18] != ele[17][19];
    ele[14][18] != ele[17][20];
    ele[14][18] != ele[17][21];
    ele[14][18] != ele[17][22];
    ele[14][18] != ele[17][23];
    ele[14][18] != ele[18][18];
    ele[14][18] != ele[19][18];
    ele[14][18] != ele[20][18];
    ele[14][18] != ele[21][18];
    ele[14][18] != ele[22][18];
    ele[14][18] != ele[23][18];
    ele[14][18] != ele[24][18];
    ele[14][18] != ele[25][18];
    ele[14][18] != ele[26][18];
    ele[14][18] != ele[27][18];
    ele[14][18] != ele[28][18];
    ele[14][18] != ele[29][18];
    ele[14][18] != ele[30][18];
    ele[14][18] != ele[31][18];
    ele[14][18] != ele[32][18];
    ele[14][18] != ele[33][18];
    ele[14][18] != ele[34][18];
    ele[14][18] != ele[35][18];
    ele[14][19] != ele[14][20];
    ele[14][19] != ele[14][21];
    ele[14][19] != ele[14][22];
    ele[14][19] != ele[14][23];
    ele[14][19] != ele[14][24];
    ele[14][19] != ele[14][25];
    ele[14][19] != ele[14][26];
    ele[14][19] != ele[14][27];
    ele[14][19] != ele[14][28];
    ele[14][19] != ele[14][29];
    ele[14][19] != ele[14][30];
    ele[14][19] != ele[14][31];
    ele[14][19] != ele[14][32];
    ele[14][19] != ele[14][33];
    ele[14][19] != ele[14][34];
    ele[14][19] != ele[14][35];
    ele[14][19] != ele[15][18];
    ele[14][19] != ele[15][19];
    ele[14][19] != ele[15][20];
    ele[14][19] != ele[15][21];
    ele[14][19] != ele[15][22];
    ele[14][19] != ele[15][23];
    ele[14][19] != ele[16][18];
    ele[14][19] != ele[16][19];
    ele[14][19] != ele[16][20];
    ele[14][19] != ele[16][21];
    ele[14][19] != ele[16][22];
    ele[14][19] != ele[16][23];
    ele[14][19] != ele[17][18];
    ele[14][19] != ele[17][19];
    ele[14][19] != ele[17][20];
    ele[14][19] != ele[17][21];
    ele[14][19] != ele[17][22];
    ele[14][19] != ele[17][23];
    ele[14][19] != ele[18][19];
    ele[14][19] != ele[19][19];
    ele[14][19] != ele[20][19];
    ele[14][19] != ele[21][19];
    ele[14][19] != ele[22][19];
    ele[14][19] != ele[23][19];
    ele[14][19] != ele[24][19];
    ele[14][19] != ele[25][19];
    ele[14][19] != ele[26][19];
    ele[14][19] != ele[27][19];
    ele[14][19] != ele[28][19];
    ele[14][19] != ele[29][19];
    ele[14][19] != ele[30][19];
    ele[14][19] != ele[31][19];
    ele[14][19] != ele[32][19];
    ele[14][19] != ele[33][19];
    ele[14][19] != ele[34][19];
    ele[14][19] != ele[35][19];
    ele[14][2] != ele[14][10];
    ele[14][2] != ele[14][11];
    ele[14][2] != ele[14][12];
    ele[14][2] != ele[14][13];
    ele[14][2] != ele[14][14];
    ele[14][2] != ele[14][15];
    ele[14][2] != ele[14][16];
    ele[14][2] != ele[14][17];
    ele[14][2] != ele[14][18];
    ele[14][2] != ele[14][19];
    ele[14][2] != ele[14][20];
    ele[14][2] != ele[14][21];
    ele[14][2] != ele[14][22];
    ele[14][2] != ele[14][23];
    ele[14][2] != ele[14][24];
    ele[14][2] != ele[14][25];
    ele[14][2] != ele[14][26];
    ele[14][2] != ele[14][27];
    ele[14][2] != ele[14][28];
    ele[14][2] != ele[14][29];
    ele[14][2] != ele[14][3];
    ele[14][2] != ele[14][30];
    ele[14][2] != ele[14][31];
    ele[14][2] != ele[14][32];
    ele[14][2] != ele[14][33];
    ele[14][2] != ele[14][34];
    ele[14][2] != ele[14][35];
    ele[14][2] != ele[14][4];
    ele[14][2] != ele[14][5];
    ele[14][2] != ele[14][6];
    ele[14][2] != ele[14][7];
    ele[14][2] != ele[14][8];
    ele[14][2] != ele[14][9];
    ele[14][2] != ele[15][0];
    ele[14][2] != ele[15][1];
    ele[14][2] != ele[15][2];
    ele[14][2] != ele[15][3];
    ele[14][2] != ele[15][4];
    ele[14][2] != ele[15][5];
    ele[14][2] != ele[16][0];
    ele[14][2] != ele[16][1];
    ele[14][2] != ele[16][2];
    ele[14][2] != ele[16][3];
    ele[14][2] != ele[16][4];
    ele[14][2] != ele[16][5];
    ele[14][2] != ele[17][0];
    ele[14][2] != ele[17][1];
    ele[14][2] != ele[17][2];
    ele[14][2] != ele[17][3];
    ele[14][2] != ele[17][4];
    ele[14][2] != ele[17][5];
    ele[14][2] != ele[18][2];
    ele[14][2] != ele[19][2];
    ele[14][2] != ele[20][2];
    ele[14][2] != ele[21][2];
    ele[14][2] != ele[22][2];
    ele[14][2] != ele[23][2];
    ele[14][2] != ele[24][2];
    ele[14][2] != ele[25][2];
    ele[14][2] != ele[26][2];
    ele[14][2] != ele[27][2];
    ele[14][2] != ele[28][2];
    ele[14][2] != ele[29][2];
    ele[14][2] != ele[30][2];
    ele[14][2] != ele[31][2];
    ele[14][2] != ele[32][2];
    ele[14][2] != ele[33][2];
    ele[14][2] != ele[34][2];
    ele[14][2] != ele[35][2];
    ele[14][20] != ele[14][21];
    ele[14][20] != ele[14][22];
    ele[14][20] != ele[14][23];
    ele[14][20] != ele[14][24];
    ele[14][20] != ele[14][25];
    ele[14][20] != ele[14][26];
    ele[14][20] != ele[14][27];
    ele[14][20] != ele[14][28];
    ele[14][20] != ele[14][29];
    ele[14][20] != ele[14][30];
    ele[14][20] != ele[14][31];
    ele[14][20] != ele[14][32];
    ele[14][20] != ele[14][33];
    ele[14][20] != ele[14][34];
    ele[14][20] != ele[14][35];
    ele[14][20] != ele[15][18];
    ele[14][20] != ele[15][19];
    ele[14][20] != ele[15][20];
    ele[14][20] != ele[15][21];
    ele[14][20] != ele[15][22];
    ele[14][20] != ele[15][23];
    ele[14][20] != ele[16][18];
    ele[14][20] != ele[16][19];
    ele[14][20] != ele[16][20];
    ele[14][20] != ele[16][21];
    ele[14][20] != ele[16][22];
    ele[14][20] != ele[16][23];
    ele[14][20] != ele[17][18];
    ele[14][20] != ele[17][19];
    ele[14][20] != ele[17][20];
    ele[14][20] != ele[17][21];
    ele[14][20] != ele[17][22];
    ele[14][20] != ele[17][23];
    ele[14][20] != ele[18][20];
    ele[14][20] != ele[19][20];
    ele[14][20] != ele[20][20];
    ele[14][20] != ele[21][20];
    ele[14][20] != ele[22][20];
    ele[14][20] != ele[23][20];
    ele[14][20] != ele[24][20];
    ele[14][20] != ele[25][20];
    ele[14][20] != ele[26][20];
    ele[14][20] != ele[27][20];
    ele[14][20] != ele[28][20];
    ele[14][20] != ele[29][20];
    ele[14][20] != ele[30][20];
    ele[14][20] != ele[31][20];
    ele[14][20] != ele[32][20];
    ele[14][20] != ele[33][20];
    ele[14][20] != ele[34][20];
    ele[14][20] != ele[35][20];
    ele[14][21] != ele[14][22];
    ele[14][21] != ele[14][23];
    ele[14][21] != ele[14][24];
    ele[14][21] != ele[14][25];
    ele[14][21] != ele[14][26];
    ele[14][21] != ele[14][27];
    ele[14][21] != ele[14][28];
    ele[14][21] != ele[14][29];
    ele[14][21] != ele[14][30];
    ele[14][21] != ele[14][31];
    ele[14][21] != ele[14][32];
    ele[14][21] != ele[14][33];
    ele[14][21] != ele[14][34];
    ele[14][21] != ele[14][35];
    ele[14][21] != ele[15][18];
    ele[14][21] != ele[15][19];
    ele[14][21] != ele[15][20];
    ele[14][21] != ele[15][21];
    ele[14][21] != ele[15][22];
    ele[14][21] != ele[15][23];
    ele[14][21] != ele[16][18];
    ele[14][21] != ele[16][19];
    ele[14][21] != ele[16][20];
    ele[14][21] != ele[16][21];
    ele[14][21] != ele[16][22];
    ele[14][21] != ele[16][23];
    ele[14][21] != ele[17][18];
    ele[14][21] != ele[17][19];
    ele[14][21] != ele[17][20];
    ele[14][21] != ele[17][21];
    ele[14][21] != ele[17][22];
    ele[14][21] != ele[17][23];
    ele[14][21] != ele[18][21];
    ele[14][21] != ele[19][21];
    ele[14][21] != ele[20][21];
    ele[14][21] != ele[21][21];
    ele[14][21] != ele[22][21];
    ele[14][21] != ele[23][21];
    ele[14][21] != ele[24][21];
    ele[14][21] != ele[25][21];
    ele[14][21] != ele[26][21];
    ele[14][21] != ele[27][21];
    ele[14][21] != ele[28][21];
    ele[14][21] != ele[29][21];
    ele[14][21] != ele[30][21];
    ele[14][21] != ele[31][21];
    ele[14][21] != ele[32][21];
    ele[14][21] != ele[33][21];
    ele[14][21] != ele[34][21];
    ele[14][21] != ele[35][21];
    ele[14][22] != ele[14][23];
    ele[14][22] != ele[14][24];
    ele[14][22] != ele[14][25];
    ele[14][22] != ele[14][26];
    ele[14][22] != ele[14][27];
    ele[14][22] != ele[14][28];
    ele[14][22] != ele[14][29];
    ele[14][22] != ele[14][30];
    ele[14][22] != ele[14][31];
    ele[14][22] != ele[14][32];
    ele[14][22] != ele[14][33];
    ele[14][22] != ele[14][34];
    ele[14][22] != ele[14][35];
    ele[14][22] != ele[15][18];
    ele[14][22] != ele[15][19];
    ele[14][22] != ele[15][20];
    ele[14][22] != ele[15][21];
    ele[14][22] != ele[15][22];
    ele[14][22] != ele[15][23];
    ele[14][22] != ele[16][18];
    ele[14][22] != ele[16][19];
    ele[14][22] != ele[16][20];
    ele[14][22] != ele[16][21];
    ele[14][22] != ele[16][22];
    ele[14][22] != ele[16][23];
    ele[14][22] != ele[17][18];
    ele[14][22] != ele[17][19];
    ele[14][22] != ele[17][20];
    ele[14][22] != ele[17][21];
    ele[14][22] != ele[17][22];
    ele[14][22] != ele[17][23];
    ele[14][22] != ele[18][22];
    ele[14][22] != ele[19][22];
    ele[14][22] != ele[20][22];
    ele[14][22] != ele[21][22];
    ele[14][22] != ele[22][22];
    ele[14][22] != ele[23][22];
    ele[14][22] != ele[24][22];
    ele[14][22] != ele[25][22];
    ele[14][22] != ele[26][22];
    ele[14][22] != ele[27][22];
    ele[14][22] != ele[28][22];
    ele[14][22] != ele[29][22];
    ele[14][22] != ele[30][22];
    ele[14][22] != ele[31][22];
    ele[14][22] != ele[32][22];
    ele[14][22] != ele[33][22];
    ele[14][22] != ele[34][22];
    ele[14][22] != ele[35][22];
    ele[14][23] != ele[14][24];
    ele[14][23] != ele[14][25];
    ele[14][23] != ele[14][26];
    ele[14][23] != ele[14][27];
    ele[14][23] != ele[14][28];
    ele[14][23] != ele[14][29];
    ele[14][23] != ele[14][30];
    ele[14][23] != ele[14][31];
    ele[14][23] != ele[14][32];
    ele[14][23] != ele[14][33];
    ele[14][23] != ele[14][34];
    ele[14][23] != ele[14][35];
    ele[14][23] != ele[15][18];
    ele[14][23] != ele[15][19];
    ele[14][23] != ele[15][20];
    ele[14][23] != ele[15][21];
    ele[14][23] != ele[15][22];
    ele[14][23] != ele[15][23];
    ele[14][23] != ele[16][18];
    ele[14][23] != ele[16][19];
    ele[14][23] != ele[16][20];
    ele[14][23] != ele[16][21];
    ele[14][23] != ele[16][22];
    ele[14][23] != ele[16][23];
    ele[14][23] != ele[17][18];
    ele[14][23] != ele[17][19];
    ele[14][23] != ele[17][20];
    ele[14][23] != ele[17][21];
    ele[14][23] != ele[17][22];
    ele[14][23] != ele[17][23];
    ele[14][23] != ele[18][23];
    ele[14][23] != ele[19][23];
    ele[14][23] != ele[20][23];
    ele[14][23] != ele[21][23];
    ele[14][23] != ele[22][23];
    ele[14][23] != ele[23][23];
    ele[14][23] != ele[24][23];
    ele[14][23] != ele[25][23];
    ele[14][23] != ele[26][23];
    ele[14][23] != ele[27][23];
    ele[14][23] != ele[28][23];
    ele[14][23] != ele[29][23];
    ele[14][23] != ele[30][23];
    ele[14][23] != ele[31][23];
    ele[14][23] != ele[32][23];
    ele[14][23] != ele[33][23];
    ele[14][23] != ele[34][23];
    ele[14][23] != ele[35][23];
    ele[14][24] != ele[14][25];
    ele[14][24] != ele[14][26];
    ele[14][24] != ele[14][27];
    ele[14][24] != ele[14][28];
    ele[14][24] != ele[14][29];
    ele[14][24] != ele[14][30];
    ele[14][24] != ele[14][31];
    ele[14][24] != ele[14][32];
    ele[14][24] != ele[14][33];
    ele[14][24] != ele[14][34];
    ele[14][24] != ele[14][35];
    ele[14][24] != ele[15][24];
    ele[14][24] != ele[15][25];
    ele[14][24] != ele[15][26];
    ele[14][24] != ele[15][27];
    ele[14][24] != ele[15][28];
    ele[14][24] != ele[15][29];
    ele[14][24] != ele[16][24];
    ele[14][24] != ele[16][25];
    ele[14][24] != ele[16][26];
    ele[14][24] != ele[16][27];
    ele[14][24] != ele[16][28];
    ele[14][24] != ele[16][29];
    ele[14][24] != ele[17][24];
    ele[14][24] != ele[17][25];
    ele[14][24] != ele[17][26];
    ele[14][24] != ele[17][27];
    ele[14][24] != ele[17][28];
    ele[14][24] != ele[17][29];
    ele[14][24] != ele[18][24];
    ele[14][24] != ele[19][24];
    ele[14][24] != ele[20][24];
    ele[14][24] != ele[21][24];
    ele[14][24] != ele[22][24];
    ele[14][24] != ele[23][24];
    ele[14][24] != ele[24][24];
    ele[14][24] != ele[25][24];
    ele[14][24] != ele[26][24];
    ele[14][24] != ele[27][24];
    ele[14][24] != ele[28][24];
    ele[14][24] != ele[29][24];
    ele[14][24] != ele[30][24];
    ele[14][24] != ele[31][24];
    ele[14][24] != ele[32][24];
    ele[14][24] != ele[33][24];
    ele[14][24] != ele[34][24];
    ele[14][24] != ele[35][24];
    ele[14][25] != ele[14][26];
    ele[14][25] != ele[14][27];
    ele[14][25] != ele[14][28];
    ele[14][25] != ele[14][29];
    ele[14][25] != ele[14][30];
    ele[14][25] != ele[14][31];
    ele[14][25] != ele[14][32];
    ele[14][25] != ele[14][33];
    ele[14][25] != ele[14][34];
    ele[14][25] != ele[14][35];
    ele[14][25] != ele[15][24];
    ele[14][25] != ele[15][25];
    ele[14][25] != ele[15][26];
    ele[14][25] != ele[15][27];
    ele[14][25] != ele[15][28];
    ele[14][25] != ele[15][29];
    ele[14][25] != ele[16][24];
    ele[14][25] != ele[16][25];
    ele[14][25] != ele[16][26];
    ele[14][25] != ele[16][27];
    ele[14][25] != ele[16][28];
    ele[14][25] != ele[16][29];
    ele[14][25] != ele[17][24];
    ele[14][25] != ele[17][25];
    ele[14][25] != ele[17][26];
    ele[14][25] != ele[17][27];
    ele[14][25] != ele[17][28];
    ele[14][25] != ele[17][29];
    ele[14][25] != ele[18][25];
    ele[14][25] != ele[19][25];
    ele[14][25] != ele[20][25];
    ele[14][25] != ele[21][25];
    ele[14][25] != ele[22][25];
    ele[14][25] != ele[23][25];
    ele[14][25] != ele[24][25];
    ele[14][25] != ele[25][25];
    ele[14][25] != ele[26][25];
    ele[14][25] != ele[27][25];
    ele[14][25] != ele[28][25];
    ele[14][25] != ele[29][25];
    ele[14][25] != ele[30][25];
    ele[14][25] != ele[31][25];
    ele[14][25] != ele[32][25];
    ele[14][25] != ele[33][25];
    ele[14][25] != ele[34][25];
    ele[14][25] != ele[35][25];
    ele[14][26] != ele[14][27];
    ele[14][26] != ele[14][28];
    ele[14][26] != ele[14][29];
    ele[14][26] != ele[14][30];
    ele[14][26] != ele[14][31];
    ele[14][26] != ele[14][32];
    ele[14][26] != ele[14][33];
    ele[14][26] != ele[14][34];
    ele[14][26] != ele[14][35];
    ele[14][26] != ele[15][24];
    ele[14][26] != ele[15][25];
    ele[14][26] != ele[15][26];
    ele[14][26] != ele[15][27];
    ele[14][26] != ele[15][28];
    ele[14][26] != ele[15][29];
    ele[14][26] != ele[16][24];
    ele[14][26] != ele[16][25];
    ele[14][26] != ele[16][26];
    ele[14][26] != ele[16][27];
    ele[14][26] != ele[16][28];
    ele[14][26] != ele[16][29];
    ele[14][26] != ele[17][24];
    ele[14][26] != ele[17][25];
    ele[14][26] != ele[17][26];
    ele[14][26] != ele[17][27];
    ele[14][26] != ele[17][28];
    ele[14][26] != ele[17][29];
    ele[14][26] != ele[18][26];
    ele[14][26] != ele[19][26];
    ele[14][26] != ele[20][26];
    ele[14][26] != ele[21][26];
    ele[14][26] != ele[22][26];
    ele[14][26] != ele[23][26];
    ele[14][26] != ele[24][26];
    ele[14][26] != ele[25][26];
    ele[14][26] != ele[26][26];
    ele[14][26] != ele[27][26];
    ele[14][26] != ele[28][26];
    ele[14][26] != ele[29][26];
    ele[14][26] != ele[30][26];
    ele[14][26] != ele[31][26];
    ele[14][26] != ele[32][26];
    ele[14][26] != ele[33][26];
    ele[14][26] != ele[34][26];
    ele[14][26] != ele[35][26];
    ele[14][27] != ele[14][28];
    ele[14][27] != ele[14][29];
    ele[14][27] != ele[14][30];
    ele[14][27] != ele[14][31];
    ele[14][27] != ele[14][32];
    ele[14][27] != ele[14][33];
    ele[14][27] != ele[14][34];
    ele[14][27] != ele[14][35];
    ele[14][27] != ele[15][24];
    ele[14][27] != ele[15][25];
    ele[14][27] != ele[15][26];
    ele[14][27] != ele[15][27];
    ele[14][27] != ele[15][28];
    ele[14][27] != ele[15][29];
    ele[14][27] != ele[16][24];
    ele[14][27] != ele[16][25];
    ele[14][27] != ele[16][26];
    ele[14][27] != ele[16][27];
    ele[14][27] != ele[16][28];
    ele[14][27] != ele[16][29];
    ele[14][27] != ele[17][24];
    ele[14][27] != ele[17][25];
    ele[14][27] != ele[17][26];
    ele[14][27] != ele[17][27];
    ele[14][27] != ele[17][28];
    ele[14][27] != ele[17][29];
    ele[14][27] != ele[18][27];
    ele[14][27] != ele[19][27];
    ele[14][27] != ele[20][27];
    ele[14][27] != ele[21][27];
    ele[14][27] != ele[22][27];
    ele[14][27] != ele[23][27];
    ele[14][27] != ele[24][27];
    ele[14][27] != ele[25][27];
    ele[14][27] != ele[26][27];
    ele[14][27] != ele[27][27];
    ele[14][27] != ele[28][27];
    ele[14][27] != ele[29][27];
    ele[14][27] != ele[30][27];
    ele[14][27] != ele[31][27];
    ele[14][27] != ele[32][27];
    ele[14][27] != ele[33][27];
    ele[14][27] != ele[34][27];
    ele[14][27] != ele[35][27];
    ele[14][28] != ele[14][29];
    ele[14][28] != ele[14][30];
    ele[14][28] != ele[14][31];
    ele[14][28] != ele[14][32];
    ele[14][28] != ele[14][33];
    ele[14][28] != ele[14][34];
    ele[14][28] != ele[14][35];
    ele[14][28] != ele[15][24];
    ele[14][28] != ele[15][25];
    ele[14][28] != ele[15][26];
    ele[14][28] != ele[15][27];
    ele[14][28] != ele[15][28];
    ele[14][28] != ele[15][29];
    ele[14][28] != ele[16][24];
    ele[14][28] != ele[16][25];
    ele[14][28] != ele[16][26];
    ele[14][28] != ele[16][27];
    ele[14][28] != ele[16][28];
    ele[14][28] != ele[16][29];
    ele[14][28] != ele[17][24];
    ele[14][28] != ele[17][25];
    ele[14][28] != ele[17][26];
    ele[14][28] != ele[17][27];
    ele[14][28] != ele[17][28];
    ele[14][28] != ele[17][29];
    ele[14][28] != ele[18][28];
    ele[14][28] != ele[19][28];
    ele[14][28] != ele[20][28];
    ele[14][28] != ele[21][28];
    ele[14][28] != ele[22][28];
    ele[14][28] != ele[23][28];
    ele[14][28] != ele[24][28];
    ele[14][28] != ele[25][28];
    ele[14][28] != ele[26][28];
    ele[14][28] != ele[27][28];
    ele[14][28] != ele[28][28];
    ele[14][28] != ele[29][28];
    ele[14][28] != ele[30][28];
    ele[14][28] != ele[31][28];
    ele[14][28] != ele[32][28];
    ele[14][28] != ele[33][28];
    ele[14][28] != ele[34][28];
    ele[14][28] != ele[35][28];
    ele[14][29] != ele[14][30];
    ele[14][29] != ele[14][31];
    ele[14][29] != ele[14][32];
    ele[14][29] != ele[14][33];
    ele[14][29] != ele[14][34];
    ele[14][29] != ele[14][35];
    ele[14][29] != ele[15][24];
    ele[14][29] != ele[15][25];
    ele[14][29] != ele[15][26];
    ele[14][29] != ele[15][27];
    ele[14][29] != ele[15][28];
    ele[14][29] != ele[15][29];
    ele[14][29] != ele[16][24];
    ele[14][29] != ele[16][25];
    ele[14][29] != ele[16][26];
    ele[14][29] != ele[16][27];
    ele[14][29] != ele[16][28];
    ele[14][29] != ele[16][29];
    ele[14][29] != ele[17][24];
    ele[14][29] != ele[17][25];
    ele[14][29] != ele[17][26];
    ele[14][29] != ele[17][27];
    ele[14][29] != ele[17][28];
    ele[14][29] != ele[17][29];
    ele[14][29] != ele[18][29];
    ele[14][29] != ele[19][29];
    ele[14][29] != ele[20][29];
    ele[14][29] != ele[21][29];
    ele[14][29] != ele[22][29];
    ele[14][29] != ele[23][29];
    ele[14][29] != ele[24][29];
    ele[14][29] != ele[25][29];
    ele[14][29] != ele[26][29];
    ele[14][29] != ele[27][29];
    ele[14][29] != ele[28][29];
    ele[14][29] != ele[29][29];
    ele[14][29] != ele[30][29];
    ele[14][29] != ele[31][29];
    ele[14][29] != ele[32][29];
    ele[14][29] != ele[33][29];
    ele[14][29] != ele[34][29];
    ele[14][29] != ele[35][29];
    ele[14][3] != ele[14][10];
    ele[14][3] != ele[14][11];
    ele[14][3] != ele[14][12];
    ele[14][3] != ele[14][13];
    ele[14][3] != ele[14][14];
    ele[14][3] != ele[14][15];
    ele[14][3] != ele[14][16];
    ele[14][3] != ele[14][17];
    ele[14][3] != ele[14][18];
    ele[14][3] != ele[14][19];
    ele[14][3] != ele[14][20];
    ele[14][3] != ele[14][21];
    ele[14][3] != ele[14][22];
    ele[14][3] != ele[14][23];
    ele[14][3] != ele[14][24];
    ele[14][3] != ele[14][25];
    ele[14][3] != ele[14][26];
    ele[14][3] != ele[14][27];
    ele[14][3] != ele[14][28];
    ele[14][3] != ele[14][29];
    ele[14][3] != ele[14][30];
    ele[14][3] != ele[14][31];
    ele[14][3] != ele[14][32];
    ele[14][3] != ele[14][33];
    ele[14][3] != ele[14][34];
    ele[14][3] != ele[14][35];
    ele[14][3] != ele[14][4];
    ele[14][3] != ele[14][5];
    ele[14][3] != ele[14][6];
    ele[14][3] != ele[14][7];
    ele[14][3] != ele[14][8];
    ele[14][3] != ele[14][9];
    ele[14][3] != ele[15][0];
    ele[14][3] != ele[15][1];
    ele[14][3] != ele[15][2];
    ele[14][3] != ele[15][3];
    ele[14][3] != ele[15][4];
    ele[14][3] != ele[15][5];
    ele[14][3] != ele[16][0];
    ele[14][3] != ele[16][1];
    ele[14][3] != ele[16][2];
    ele[14][3] != ele[16][3];
    ele[14][3] != ele[16][4];
    ele[14][3] != ele[16][5];
    ele[14][3] != ele[17][0];
    ele[14][3] != ele[17][1];
    ele[14][3] != ele[17][2];
    ele[14][3] != ele[17][3];
    ele[14][3] != ele[17][4];
    ele[14][3] != ele[17][5];
    ele[14][3] != ele[18][3];
    ele[14][3] != ele[19][3];
    ele[14][3] != ele[20][3];
    ele[14][3] != ele[21][3];
    ele[14][3] != ele[22][3];
    ele[14][3] != ele[23][3];
    ele[14][3] != ele[24][3];
    ele[14][3] != ele[25][3];
    ele[14][3] != ele[26][3];
    ele[14][3] != ele[27][3];
    ele[14][3] != ele[28][3];
    ele[14][3] != ele[29][3];
    ele[14][3] != ele[30][3];
    ele[14][3] != ele[31][3];
    ele[14][3] != ele[32][3];
    ele[14][3] != ele[33][3];
    ele[14][3] != ele[34][3];
    ele[14][3] != ele[35][3];
    ele[14][30] != ele[14][31];
    ele[14][30] != ele[14][32];
    ele[14][30] != ele[14][33];
    ele[14][30] != ele[14][34];
    ele[14][30] != ele[14][35];
    ele[14][30] != ele[15][30];
    ele[14][30] != ele[15][31];
    ele[14][30] != ele[15][32];
    ele[14][30] != ele[15][33];
    ele[14][30] != ele[15][34];
    ele[14][30] != ele[15][35];
    ele[14][30] != ele[16][30];
    ele[14][30] != ele[16][31];
    ele[14][30] != ele[16][32];
    ele[14][30] != ele[16][33];
    ele[14][30] != ele[16][34];
    ele[14][30] != ele[16][35];
    ele[14][30] != ele[17][30];
    ele[14][30] != ele[17][31];
    ele[14][30] != ele[17][32];
    ele[14][30] != ele[17][33];
    ele[14][30] != ele[17][34];
    ele[14][30] != ele[17][35];
    ele[14][30] != ele[18][30];
    ele[14][30] != ele[19][30];
    ele[14][30] != ele[20][30];
    ele[14][30] != ele[21][30];
    ele[14][30] != ele[22][30];
    ele[14][30] != ele[23][30];
    ele[14][30] != ele[24][30];
    ele[14][30] != ele[25][30];
    ele[14][30] != ele[26][30];
    ele[14][30] != ele[27][30];
    ele[14][30] != ele[28][30];
    ele[14][30] != ele[29][30];
    ele[14][30] != ele[30][30];
    ele[14][30] != ele[31][30];
    ele[14][30] != ele[32][30];
    ele[14][30] != ele[33][30];
    ele[14][30] != ele[34][30];
    ele[14][30] != ele[35][30];
    ele[14][31] != ele[14][32];
    ele[14][31] != ele[14][33];
    ele[14][31] != ele[14][34];
    ele[14][31] != ele[14][35];
    ele[14][31] != ele[15][30];
    ele[14][31] != ele[15][31];
    ele[14][31] != ele[15][32];
    ele[14][31] != ele[15][33];
    ele[14][31] != ele[15][34];
    ele[14][31] != ele[15][35];
    ele[14][31] != ele[16][30];
    ele[14][31] != ele[16][31];
    ele[14][31] != ele[16][32];
    ele[14][31] != ele[16][33];
    ele[14][31] != ele[16][34];
    ele[14][31] != ele[16][35];
    ele[14][31] != ele[17][30];
    ele[14][31] != ele[17][31];
    ele[14][31] != ele[17][32];
    ele[14][31] != ele[17][33];
    ele[14][31] != ele[17][34];
    ele[14][31] != ele[17][35];
    ele[14][31] != ele[18][31];
    ele[14][31] != ele[19][31];
    ele[14][31] != ele[20][31];
    ele[14][31] != ele[21][31];
    ele[14][31] != ele[22][31];
    ele[14][31] != ele[23][31];
    ele[14][31] != ele[24][31];
    ele[14][31] != ele[25][31];
    ele[14][31] != ele[26][31];
    ele[14][31] != ele[27][31];
    ele[14][31] != ele[28][31];
    ele[14][31] != ele[29][31];
    ele[14][31] != ele[30][31];
    ele[14][31] != ele[31][31];
    ele[14][31] != ele[32][31];
    ele[14][31] != ele[33][31];
    ele[14][31] != ele[34][31];
    ele[14][31] != ele[35][31];
    ele[14][32] != ele[14][33];
    ele[14][32] != ele[14][34];
    ele[14][32] != ele[14][35];
    ele[14][32] != ele[15][30];
    ele[14][32] != ele[15][31];
    ele[14][32] != ele[15][32];
    ele[14][32] != ele[15][33];
    ele[14][32] != ele[15][34];
    ele[14][32] != ele[15][35];
    ele[14][32] != ele[16][30];
    ele[14][32] != ele[16][31];
    ele[14][32] != ele[16][32];
    ele[14][32] != ele[16][33];
    ele[14][32] != ele[16][34];
    ele[14][32] != ele[16][35];
    ele[14][32] != ele[17][30];
    ele[14][32] != ele[17][31];
    ele[14][32] != ele[17][32];
    ele[14][32] != ele[17][33];
    ele[14][32] != ele[17][34];
    ele[14][32] != ele[17][35];
    ele[14][32] != ele[18][32];
    ele[14][32] != ele[19][32];
    ele[14][32] != ele[20][32];
    ele[14][32] != ele[21][32];
    ele[14][32] != ele[22][32];
    ele[14][32] != ele[23][32];
    ele[14][32] != ele[24][32];
    ele[14][32] != ele[25][32];
    ele[14][32] != ele[26][32];
    ele[14][32] != ele[27][32];
    ele[14][32] != ele[28][32];
    ele[14][32] != ele[29][32];
    ele[14][32] != ele[30][32];
    ele[14][32] != ele[31][32];
    ele[14][32] != ele[32][32];
    ele[14][32] != ele[33][32];
    ele[14][32] != ele[34][32];
    ele[14][32] != ele[35][32];
    ele[14][33] != ele[14][34];
    ele[14][33] != ele[14][35];
    ele[14][33] != ele[15][30];
    ele[14][33] != ele[15][31];
    ele[14][33] != ele[15][32];
    ele[14][33] != ele[15][33];
    ele[14][33] != ele[15][34];
    ele[14][33] != ele[15][35];
    ele[14][33] != ele[16][30];
    ele[14][33] != ele[16][31];
    ele[14][33] != ele[16][32];
    ele[14][33] != ele[16][33];
    ele[14][33] != ele[16][34];
    ele[14][33] != ele[16][35];
    ele[14][33] != ele[17][30];
    ele[14][33] != ele[17][31];
    ele[14][33] != ele[17][32];
    ele[14][33] != ele[17][33];
    ele[14][33] != ele[17][34];
    ele[14][33] != ele[17][35];
    ele[14][33] != ele[18][33];
    ele[14][33] != ele[19][33];
    ele[14][33] != ele[20][33];
    ele[14][33] != ele[21][33];
    ele[14][33] != ele[22][33];
    ele[14][33] != ele[23][33];
    ele[14][33] != ele[24][33];
    ele[14][33] != ele[25][33];
    ele[14][33] != ele[26][33];
    ele[14][33] != ele[27][33];
    ele[14][33] != ele[28][33];
    ele[14][33] != ele[29][33];
    ele[14][33] != ele[30][33];
    ele[14][33] != ele[31][33];
    ele[14][33] != ele[32][33];
    ele[14][33] != ele[33][33];
    ele[14][33] != ele[34][33];
    ele[14][33] != ele[35][33];
    ele[14][34] != ele[14][35];
    ele[14][34] != ele[15][30];
    ele[14][34] != ele[15][31];
    ele[14][34] != ele[15][32];
    ele[14][34] != ele[15][33];
    ele[14][34] != ele[15][34];
    ele[14][34] != ele[15][35];
    ele[14][34] != ele[16][30];
    ele[14][34] != ele[16][31];
    ele[14][34] != ele[16][32];
    ele[14][34] != ele[16][33];
    ele[14][34] != ele[16][34];
    ele[14][34] != ele[16][35];
    ele[14][34] != ele[17][30];
    ele[14][34] != ele[17][31];
    ele[14][34] != ele[17][32];
    ele[14][34] != ele[17][33];
    ele[14][34] != ele[17][34];
    ele[14][34] != ele[17][35];
    ele[14][34] != ele[18][34];
    ele[14][34] != ele[19][34];
    ele[14][34] != ele[20][34];
    ele[14][34] != ele[21][34];
    ele[14][34] != ele[22][34];
    ele[14][34] != ele[23][34];
    ele[14][34] != ele[24][34];
    ele[14][34] != ele[25][34];
    ele[14][34] != ele[26][34];
    ele[14][34] != ele[27][34];
    ele[14][34] != ele[28][34];
    ele[14][34] != ele[29][34];
    ele[14][34] != ele[30][34];
    ele[14][34] != ele[31][34];
    ele[14][34] != ele[32][34];
    ele[14][34] != ele[33][34];
    ele[14][34] != ele[34][34];
    ele[14][34] != ele[35][34];
    ele[14][35] != ele[15][30];
    ele[14][35] != ele[15][31];
    ele[14][35] != ele[15][32];
    ele[14][35] != ele[15][33];
    ele[14][35] != ele[15][34];
    ele[14][35] != ele[15][35];
    ele[14][35] != ele[16][30];
    ele[14][35] != ele[16][31];
    ele[14][35] != ele[16][32];
    ele[14][35] != ele[16][33];
    ele[14][35] != ele[16][34];
    ele[14][35] != ele[16][35];
    ele[14][35] != ele[17][30];
    ele[14][35] != ele[17][31];
    ele[14][35] != ele[17][32];
    ele[14][35] != ele[17][33];
    ele[14][35] != ele[17][34];
    ele[14][35] != ele[17][35];
    ele[14][35] != ele[18][35];
    ele[14][35] != ele[19][35];
    ele[14][35] != ele[20][35];
    ele[14][35] != ele[21][35];
    ele[14][35] != ele[22][35];
    ele[14][35] != ele[23][35];
    ele[14][35] != ele[24][35];
    ele[14][35] != ele[25][35];
    ele[14][35] != ele[26][35];
    ele[14][35] != ele[27][35];
    ele[14][35] != ele[28][35];
    ele[14][35] != ele[29][35];
    ele[14][35] != ele[30][35];
    ele[14][35] != ele[31][35];
    ele[14][35] != ele[32][35];
    ele[14][35] != ele[33][35];
    ele[14][35] != ele[34][35];
    ele[14][35] != ele[35][35];
    ele[14][4] != ele[14][10];
    ele[14][4] != ele[14][11];
    ele[14][4] != ele[14][12];
    ele[14][4] != ele[14][13];
    ele[14][4] != ele[14][14];
    ele[14][4] != ele[14][15];
    ele[14][4] != ele[14][16];
    ele[14][4] != ele[14][17];
    ele[14][4] != ele[14][18];
    ele[14][4] != ele[14][19];
    ele[14][4] != ele[14][20];
    ele[14][4] != ele[14][21];
    ele[14][4] != ele[14][22];
    ele[14][4] != ele[14][23];
    ele[14][4] != ele[14][24];
    ele[14][4] != ele[14][25];
    ele[14][4] != ele[14][26];
    ele[14][4] != ele[14][27];
    ele[14][4] != ele[14][28];
    ele[14][4] != ele[14][29];
    ele[14][4] != ele[14][30];
    ele[14][4] != ele[14][31];
    ele[14][4] != ele[14][32];
    ele[14][4] != ele[14][33];
    ele[14][4] != ele[14][34];
    ele[14][4] != ele[14][35];
    ele[14][4] != ele[14][5];
    ele[14][4] != ele[14][6];
    ele[14][4] != ele[14][7];
    ele[14][4] != ele[14][8];
    ele[14][4] != ele[14][9];
    ele[14][4] != ele[15][0];
    ele[14][4] != ele[15][1];
    ele[14][4] != ele[15][2];
    ele[14][4] != ele[15][3];
    ele[14][4] != ele[15][4];
    ele[14][4] != ele[15][5];
    ele[14][4] != ele[16][0];
    ele[14][4] != ele[16][1];
    ele[14][4] != ele[16][2];
    ele[14][4] != ele[16][3];
    ele[14][4] != ele[16][4];
    ele[14][4] != ele[16][5];
    ele[14][4] != ele[17][0];
    ele[14][4] != ele[17][1];
    ele[14][4] != ele[17][2];
    ele[14][4] != ele[17][3];
    ele[14][4] != ele[17][4];
    ele[14][4] != ele[17][5];
    ele[14][4] != ele[18][4];
    ele[14][4] != ele[19][4];
    ele[14][4] != ele[20][4];
    ele[14][4] != ele[21][4];
    ele[14][4] != ele[22][4];
    ele[14][4] != ele[23][4];
    ele[14][4] != ele[24][4];
    ele[14][4] != ele[25][4];
    ele[14][4] != ele[26][4];
    ele[14][4] != ele[27][4];
    ele[14][4] != ele[28][4];
    ele[14][4] != ele[29][4];
    ele[14][4] != ele[30][4];
    ele[14][4] != ele[31][4];
    ele[14][4] != ele[32][4];
    ele[14][4] != ele[33][4];
    ele[14][4] != ele[34][4];
    ele[14][4] != ele[35][4];
    ele[14][5] != ele[14][10];
    ele[14][5] != ele[14][11];
    ele[14][5] != ele[14][12];
    ele[14][5] != ele[14][13];
    ele[14][5] != ele[14][14];
    ele[14][5] != ele[14][15];
    ele[14][5] != ele[14][16];
    ele[14][5] != ele[14][17];
    ele[14][5] != ele[14][18];
    ele[14][5] != ele[14][19];
    ele[14][5] != ele[14][20];
    ele[14][5] != ele[14][21];
    ele[14][5] != ele[14][22];
    ele[14][5] != ele[14][23];
    ele[14][5] != ele[14][24];
    ele[14][5] != ele[14][25];
    ele[14][5] != ele[14][26];
    ele[14][5] != ele[14][27];
    ele[14][5] != ele[14][28];
    ele[14][5] != ele[14][29];
    ele[14][5] != ele[14][30];
    ele[14][5] != ele[14][31];
    ele[14][5] != ele[14][32];
    ele[14][5] != ele[14][33];
    ele[14][5] != ele[14][34];
    ele[14][5] != ele[14][35];
    ele[14][5] != ele[14][6];
    ele[14][5] != ele[14][7];
    ele[14][5] != ele[14][8];
    ele[14][5] != ele[14][9];
    ele[14][5] != ele[15][0];
    ele[14][5] != ele[15][1];
    ele[14][5] != ele[15][2];
    ele[14][5] != ele[15][3];
    ele[14][5] != ele[15][4];
    ele[14][5] != ele[15][5];
    ele[14][5] != ele[16][0];
    ele[14][5] != ele[16][1];
    ele[14][5] != ele[16][2];
    ele[14][5] != ele[16][3];
    ele[14][5] != ele[16][4];
    ele[14][5] != ele[16][5];
    ele[14][5] != ele[17][0];
    ele[14][5] != ele[17][1];
    ele[14][5] != ele[17][2];
    ele[14][5] != ele[17][3];
    ele[14][5] != ele[17][4];
    ele[14][5] != ele[17][5];
    ele[14][5] != ele[18][5];
    ele[14][5] != ele[19][5];
    ele[14][5] != ele[20][5];
    ele[14][5] != ele[21][5];
    ele[14][5] != ele[22][5];
    ele[14][5] != ele[23][5];
    ele[14][5] != ele[24][5];
    ele[14][5] != ele[25][5];
    ele[14][5] != ele[26][5];
    ele[14][5] != ele[27][5];
    ele[14][5] != ele[28][5];
    ele[14][5] != ele[29][5];
    ele[14][5] != ele[30][5];
    ele[14][5] != ele[31][5];
    ele[14][5] != ele[32][5];
    ele[14][5] != ele[33][5];
    ele[14][5] != ele[34][5];
    ele[14][5] != ele[35][5];
    ele[14][6] != ele[14][10];
    ele[14][6] != ele[14][11];
    ele[14][6] != ele[14][12];
    ele[14][6] != ele[14][13];
    ele[14][6] != ele[14][14];
    ele[14][6] != ele[14][15];
    ele[14][6] != ele[14][16];
    ele[14][6] != ele[14][17];
    ele[14][6] != ele[14][18];
    ele[14][6] != ele[14][19];
    ele[14][6] != ele[14][20];
    ele[14][6] != ele[14][21];
    ele[14][6] != ele[14][22];
    ele[14][6] != ele[14][23];
    ele[14][6] != ele[14][24];
    ele[14][6] != ele[14][25];
    ele[14][6] != ele[14][26];
    ele[14][6] != ele[14][27];
    ele[14][6] != ele[14][28];
    ele[14][6] != ele[14][29];
    ele[14][6] != ele[14][30];
    ele[14][6] != ele[14][31];
    ele[14][6] != ele[14][32];
    ele[14][6] != ele[14][33];
    ele[14][6] != ele[14][34];
    ele[14][6] != ele[14][35];
    ele[14][6] != ele[14][7];
    ele[14][6] != ele[14][8];
    ele[14][6] != ele[14][9];
    ele[14][6] != ele[15][10];
    ele[14][6] != ele[15][11];
    ele[14][6] != ele[15][6];
    ele[14][6] != ele[15][7];
    ele[14][6] != ele[15][8];
    ele[14][6] != ele[15][9];
    ele[14][6] != ele[16][10];
    ele[14][6] != ele[16][11];
    ele[14][6] != ele[16][6];
    ele[14][6] != ele[16][7];
    ele[14][6] != ele[16][8];
    ele[14][6] != ele[16][9];
    ele[14][6] != ele[17][10];
    ele[14][6] != ele[17][11];
    ele[14][6] != ele[17][6];
    ele[14][6] != ele[17][7];
    ele[14][6] != ele[17][8];
    ele[14][6] != ele[17][9];
    ele[14][6] != ele[18][6];
    ele[14][6] != ele[19][6];
    ele[14][6] != ele[20][6];
    ele[14][6] != ele[21][6];
    ele[14][6] != ele[22][6];
    ele[14][6] != ele[23][6];
    ele[14][6] != ele[24][6];
    ele[14][6] != ele[25][6];
    ele[14][6] != ele[26][6];
    ele[14][6] != ele[27][6];
    ele[14][6] != ele[28][6];
    ele[14][6] != ele[29][6];
    ele[14][6] != ele[30][6];
    ele[14][6] != ele[31][6];
    ele[14][6] != ele[32][6];
    ele[14][6] != ele[33][6];
    ele[14][6] != ele[34][6];
    ele[14][6] != ele[35][6];
    ele[14][7] != ele[14][10];
    ele[14][7] != ele[14][11];
    ele[14][7] != ele[14][12];
    ele[14][7] != ele[14][13];
    ele[14][7] != ele[14][14];
    ele[14][7] != ele[14][15];
    ele[14][7] != ele[14][16];
    ele[14][7] != ele[14][17];
    ele[14][7] != ele[14][18];
    ele[14][7] != ele[14][19];
    ele[14][7] != ele[14][20];
    ele[14][7] != ele[14][21];
    ele[14][7] != ele[14][22];
    ele[14][7] != ele[14][23];
    ele[14][7] != ele[14][24];
    ele[14][7] != ele[14][25];
    ele[14][7] != ele[14][26];
    ele[14][7] != ele[14][27];
    ele[14][7] != ele[14][28];
    ele[14][7] != ele[14][29];
    ele[14][7] != ele[14][30];
    ele[14][7] != ele[14][31];
    ele[14][7] != ele[14][32];
    ele[14][7] != ele[14][33];
    ele[14][7] != ele[14][34];
    ele[14][7] != ele[14][35];
    ele[14][7] != ele[14][8];
    ele[14][7] != ele[14][9];
    ele[14][7] != ele[15][10];
    ele[14][7] != ele[15][11];
    ele[14][7] != ele[15][6];
    ele[14][7] != ele[15][7];
    ele[14][7] != ele[15][8];
    ele[14][7] != ele[15][9];
    ele[14][7] != ele[16][10];
    ele[14][7] != ele[16][11];
    ele[14][7] != ele[16][6];
    ele[14][7] != ele[16][7];
    ele[14][7] != ele[16][8];
    ele[14][7] != ele[16][9];
    ele[14][7] != ele[17][10];
    ele[14][7] != ele[17][11];
    ele[14][7] != ele[17][6];
    ele[14][7] != ele[17][7];
    ele[14][7] != ele[17][8];
    ele[14][7] != ele[17][9];
    ele[14][7] != ele[18][7];
    ele[14][7] != ele[19][7];
    ele[14][7] != ele[20][7];
    ele[14][7] != ele[21][7];
    ele[14][7] != ele[22][7];
    ele[14][7] != ele[23][7];
    ele[14][7] != ele[24][7];
    ele[14][7] != ele[25][7];
    ele[14][7] != ele[26][7];
    ele[14][7] != ele[27][7];
    ele[14][7] != ele[28][7];
    ele[14][7] != ele[29][7];
    ele[14][7] != ele[30][7];
    ele[14][7] != ele[31][7];
    ele[14][7] != ele[32][7];
    ele[14][7] != ele[33][7];
    ele[14][7] != ele[34][7];
    ele[14][7] != ele[35][7];
    ele[14][8] != ele[14][10];
    ele[14][8] != ele[14][11];
    ele[14][8] != ele[14][12];
    ele[14][8] != ele[14][13];
    ele[14][8] != ele[14][14];
    ele[14][8] != ele[14][15];
    ele[14][8] != ele[14][16];
    ele[14][8] != ele[14][17];
    ele[14][8] != ele[14][18];
    ele[14][8] != ele[14][19];
    ele[14][8] != ele[14][20];
    ele[14][8] != ele[14][21];
    ele[14][8] != ele[14][22];
    ele[14][8] != ele[14][23];
    ele[14][8] != ele[14][24];
    ele[14][8] != ele[14][25];
    ele[14][8] != ele[14][26];
    ele[14][8] != ele[14][27];
    ele[14][8] != ele[14][28];
    ele[14][8] != ele[14][29];
    ele[14][8] != ele[14][30];
    ele[14][8] != ele[14][31];
    ele[14][8] != ele[14][32];
    ele[14][8] != ele[14][33];
    ele[14][8] != ele[14][34];
    ele[14][8] != ele[14][35];
    ele[14][8] != ele[14][9];
    ele[14][8] != ele[15][10];
    ele[14][8] != ele[15][11];
    ele[14][8] != ele[15][6];
    ele[14][8] != ele[15][7];
    ele[14][8] != ele[15][8];
    ele[14][8] != ele[15][9];
    ele[14][8] != ele[16][10];
    ele[14][8] != ele[16][11];
    ele[14][8] != ele[16][6];
    ele[14][8] != ele[16][7];
    ele[14][8] != ele[16][8];
    ele[14][8] != ele[16][9];
    ele[14][8] != ele[17][10];
    ele[14][8] != ele[17][11];
    ele[14][8] != ele[17][6];
    ele[14][8] != ele[17][7];
    ele[14][8] != ele[17][8];
    ele[14][8] != ele[17][9];
    ele[14][8] != ele[18][8];
    ele[14][8] != ele[19][8];
    ele[14][8] != ele[20][8];
    ele[14][8] != ele[21][8];
    ele[14][8] != ele[22][8];
    ele[14][8] != ele[23][8];
    ele[14][8] != ele[24][8];
    ele[14][8] != ele[25][8];
    ele[14][8] != ele[26][8];
    ele[14][8] != ele[27][8];
    ele[14][8] != ele[28][8];
    ele[14][8] != ele[29][8];
    ele[14][8] != ele[30][8];
    ele[14][8] != ele[31][8];
    ele[14][8] != ele[32][8];
    ele[14][8] != ele[33][8];
    ele[14][8] != ele[34][8];
    ele[14][8] != ele[35][8];
    ele[14][9] != ele[14][10];
    ele[14][9] != ele[14][11];
    ele[14][9] != ele[14][12];
    ele[14][9] != ele[14][13];
    ele[14][9] != ele[14][14];
    ele[14][9] != ele[14][15];
    ele[14][9] != ele[14][16];
    ele[14][9] != ele[14][17];
    ele[14][9] != ele[14][18];
    ele[14][9] != ele[14][19];
    ele[14][9] != ele[14][20];
    ele[14][9] != ele[14][21];
    ele[14][9] != ele[14][22];
    ele[14][9] != ele[14][23];
    ele[14][9] != ele[14][24];
    ele[14][9] != ele[14][25];
    ele[14][9] != ele[14][26];
    ele[14][9] != ele[14][27];
    ele[14][9] != ele[14][28];
    ele[14][9] != ele[14][29];
    ele[14][9] != ele[14][30];
    ele[14][9] != ele[14][31];
    ele[14][9] != ele[14][32];
    ele[14][9] != ele[14][33];
    ele[14][9] != ele[14][34];
    ele[14][9] != ele[14][35];
    ele[14][9] != ele[15][10];
    ele[14][9] != ele[15][11];
    ele[14][9] != ele[15][6];
    ele[14][9] != ele[15][7];
    ele[14][9] != ele[15][8];
    ele[14][9] != ele[15][9];
    ele[14][9] != ele[16][10];
    ele[14][9] != ele[16][11];
    ele[14][9] != ele[16][6];
    ele[14][9] != ele[16][7];
    ele[14][9] != ele[16][8];
    ele[14][9] != ele[16][9];
    ele[14][9] != ele[17][10];
    ele[14][9] != ele[17][11];
    ele[14][9] != ele[17][6];
    ele[14][9] != ele[17][7];
    ele[14][9] != ele[17][8];
    ele[14][9] != ele[17][9];
    ele[14][9] != ele[18][9];
    ele[14][9] != ele[19][9];
    ele[14][9] != ele[20][9];
    ele[14][9] != ele[21][9];
    ele[14][9] != ele[22][9];
    ele[14][9] != ele[23][9];
    ele[14][9] != ele[24][9];
    ele[14][9] != ele[25][9];
    ele[14][9] != ele[26][9];
    ele[14][9] != ele[27][9];
    ele[14][9] != ele[28][9];
    ele[14][9] != ele[29][9];
    ele[14][9] != ele[30][9];
    ele[14][9] != ele[31][9];
    ele[14][9] != ele[32][9];
    ele[14][9] != ele[33][9];
    ele[14][9] != ele[34][9];
    ele[14][9] != ele[35][9];
    ele[15][0] != ele[15][1];
    ele[15][0] != ele[15][10];
    ele[15][0] != ele[15][11];
    ele[15][0] != ele[15][12];
    ele[15][0] != ele[15][13];
    ele[15][0] != ele[15][14];
    ele[15][0] != ele[15][15];
    ele[15][0] != ele[15][16];
    ele[15][0] != ele[15][17];
    ele[15][0] != ele[15][18];
    ele[15][0] != ele[15][19];
    ele[15][0] != ele[15][2];
    ele[15][0] != ele[15][20];
    ele[15][0] != ele[15][21];
    ele[15][0] != ele[15][22];
    ele[15][0] != ele[15][23];
    ele[15][0] != ele[15][24];
    ele[15][0] != ele[15][25];
    ele[15][0] != ele[15][26];
    ele[15][0] != ele[15][27];
    ele[15][0] != ele[15][28];
    ele[15][0] != ele[15][29];
    ele[15][0] != ele[15][3];
    ele[15][0] != ele[15][30];
    ele[15][0] != ele[15][31];
    ele[15][0] != ele[15][32];
    ele[15][0] != ele[15][33];
    ele[15][0] != ele[15][34];
    ele[15][0] != ele[15][35];
    ele[15][0] != ele[15][4];
    ele[15][0] != ele[15][5];
    ele[15][0] != ele[15][6];
    ele[15][0] != ele[15][7];
    ele[15][0] != ele[15][8];
    ele[15][0] != ele[15][9];
    ele[15][0] != ele[16][0];
    ele[15][0] != ele[16][1];
    ele[15][0] != ele[16][2];
    ele[15][0] != ele[16][3];
    ele[15][0] != ele[16][4];
    ele[15][0] != ele[16][5];
    ele[15][0] != ele[17][0];
    ele[15][0] != ele[17][1];
    ele[15][0] != ele[17][2];
    ele[15][0] != ele[17][3];
    ele[15][0] != ele[17][4];
    ele[15][0] != ele[17][5];
    ele[15][0] != ele[18][0];
    ele[15][0] != ele[19][0];
    ele[15][0] != ele[20][0];
    ele[15][0] != ele[21][0];
    ele[15][0] != ele[22][0];
    ele[15][0] != ele[23][0];
    ele[15][0] != ele[24][0];
    ele[15][0] != ele[25][0];
    ele[15][0] != ele[26][0];
    ele[15][0] != ele[27][0];
    ele[15][0] != ele[28][0];
    ele[15][0] != ele[29][0];
    ele[15][0] != ele[30][0];
    ele[15][0] != ele[31][0];
    ele[15][0] != ele[32][0];
    ele[15][0] != ele[33][0];
    ele[15][0] != ele[34][0];
    ele[15][0] != ele[35][0];
    ele[15][1] != ele[15][10];
    ele[15][1] != ele[15][11];
    ele[15][1] != ele[15][12];
    ele[15][1] != ele[15][13];
    ele[15][1] != ele[15][14];
    ele[15][1] != ele[15][15];
    ele[15][1] != ele[15][16];
    ele[15][1] != ele[15][17];
    ele[15][1] != ele[15][18];
    ele[15][1] != ele[15][19];
    ele[15][1] != ele[15][2];
    ele[15][1] != ele[15][20];
    ele[15][1] != ele[15][21];
    ele[15][1] != ele[15][22];
    ele[15][1] != ele[15][23];
    ele[15][1] != ele[15][24];
    ele[15][1] != ele[15][25];
    ele[15][1] != ele[15][26];
    ele[15][1] != ele[15][27];
    ele[15][1] != ele[15][28];
    ele[15][1] != ele[15][29];
    ele[15][1] != ele[15][3];
    ele[15][1] != ele[15][30];
    ele[15][1] != ele[15][31];
    ele[15][1] != ele[15][32];
    ele[15][1] != ele[15][33];
    ele[15][1] != ele[15][34];
    ele[15][1] != ele[15][35];
    ele[15][1] != ele[15][4];
    ele[15][1] != ele[15][5];
    ele[15][1] != ele[15][6];
    ele[15][1] != ele[15][7];
    ele[15][1] != ele[15][8];
    ele[15][1] != ele[15][9];
    ele[15][1] != ele[16][0];
    ele[15][1] != ele[16][1];
    ele[15][1] != ele[16][2];
    ele[15][1] != ele[16][3];
    ele[15][1] != ele[16][4];
    ele[15][1] != ele[16][5];
    ele[15][1] != ele[17][0];
    ele[15][1] != ele[17][1];
    ele[15][1] != ele[17][2];
    ele[15][1] != ele[17][3];
    ele[15][1] != ele[17][4];
    ele[15][1] != ele[17][5];
    ele[15][1] != ele[18][1];
    ele[15][1] != ele[19][1];
    ele[15][1] != ele[20][1];
    ele[15][1] != ele[21][1];
    ele[15][1] != ele[22][1];
    ele[15][1] != ele[23][1];
    ele[15][1] != ele[24][1];
    ele[15][1] != ele[25][1];
    ele[15][1] != ele[26][1];
    ele[15][1] != ele[27][1];
    ele[15][1] != ele[28][1];
    ele[15][1] != ele[29][1];
    ele[15][1] != ele[30][1];
    ele[15][1] != ele[31][1];
    ele[15][1] != ele[32][1];
    ele[15][1] != ele[33][1];
    ele[15][1] != ele[34][1];
    ele[15][1] != ele[35][1];
    ele[15][10] != ele[15][11];
    ele[15][10] != ele[15][12];
    ele[15][10] != ele[15][13];
    ele[15][10] != ele[15][14];
    ele[15][10] != ele[15][15];
    ele[15][10] != ele[15][16];
    ele[15][10] != ele[15][17];
    ele[15][10] != ele[15][18];
    ele[15][10] != ele[15][19];
    ele[15][10] != ele[15][20];
    ele[15][10] != ele[15][21];
    ele[15][10] != ele[15][22];
    ele[15][10] != ele[15][23];
    ele[15][10] != ele[15][24];
    ele[15][10] != ele[15][25];
    ele[15][10] != ele[15][26];
    ele[15][10] != ele[15][27];
    ele[15][10] != ele[15][28];
    ele[15][10] != ele[15][29];
    ele[15][10] != ele[15][30];
    ele[15][10] != ele[15][31];
    ele[15][10] != ele[15][32];
    ele[15][10] != ele[15][33];
    ele[15][10] != ele[15][34];
    ele[15][10] != ele[15][35];
    ele[15][10] != ele[16][10];
    ele[15][10] != ele[16][11];
    ele[15][10] != ele[16][6];
    ele[15][10] != ele[16][7];
    ele[15][10] != ele[16][8];
    ele[15][10] != ele[16][9];
    ele[15][10] != ele[17][10];
    ele[15][10] != ele[17][11];
    ele[15][10] != ele[17][6];
    ele[15][10] != ele[17][7];
    ele[15][10] != ele[17][8];
    ele[15][10] != ele[17][9];
    ele[15][10] != ele[18][10];
    ele[15][10] != ele[19][10];
    ele[15][10] != ele[20][10];
    ele[15][10] != ele[21][10];
    ele[15][10] != ele[22][10];
    ele[15][10] != ele[23][10];
    ele[15][10] != ele[24][10];
    ele[15][10] != ele[25][10];
    ele[15][10] != ele[26][10];
    ele[15][10] != ele[27][10];
    ele[15][10] != ele[28][10];
    ele[15][10] != ele[29][10];
    ele[15][10] != ele[30][10];
    ele[15][10] != ele[31][10];
    ele[15][10] != ele[32][10];
    ele[15][10] != ele[33][10];
    ele[15][10] != ele[34][10];
    ele[15][10] != ele[35][10];
    ele[15][11] != ele[15][12];
    ele[15][11] != ele[15][13];
    ele[15][11] != ele[15][14];
    ele[15][11] != ele[15][15];
    ele[15][11] != ele[15][16];
    ele[15][11] != ele[15][17];
    ele[15][11] != ele[15][18];
    ele[15][11] != ele[15][19];
    ele[15][11] != ele[15][20];
    ele[15][11] != ele[15][21];
    ele[15][11] != ele[15][22];
    ele[15][11] != ele[15][23];
    ele[15][11] != ele[15][24];
    ele[15][11] != ele[15][25];
    ele[15][11] != ele[15][26];
    ele[15][11] != ele[15][27];
    ele[15][11] != ele[15][28];
    ele[15][11] != ele[15][29];
    ele[15][11] != ele[15][30];
    ele[15][11] != ele[15][31];
    ele[15][11] != ele[15][32];
    ele[15][11] != ele[15][33];
    ele[15][11] != ele[15][34];
    ele[15][11] != ele[15][35];
    ele[15][11] != ele[16][10];
    ele[15][11] != ele[16][11];
    ele[15][11] != ele[16][6];
    ele[15][11] != ele[16][7];
    ele[15][11] != ele[16][8];
    ele[15][11] != ele[16][9];
    ele[15][11] != ele[17][10];
    ele[15][11] != ele[17][11];
    ele[15][11] != ele[17][6];
    ele[15][11] != ele[17][7];
    ele[15][11] != ele[17][8];
    ele[15][11] != ele[17][9];
    ele[15][11] != ele[18][11];
    ele[15][11] != ele[19][11];
    ele[15][11] != ele[20][11];
    ele[15][11] != ele[21][11];
    ele[15][11] != ele[22][11];
    ele[15][11] != ele[23][11];
    ele[15][11] != ele[24][11];
    ele[15][11] != ele[25][11];
    ele[15][11] != ele[26][11];
    ele[15][11] != ele[27][11];
    ele[15][11] != ele[28][11];
    ele[15][11] != ele[29][11];
    ele[15][11] != ele[30][11];
    ele[15][11] != ele[31][11];
    ele[15][11] != ele[32][11];
    ele[15][11] != ele[33][11];
    ele[15][11] != ele[34][11];
    ele[15][11] != ele[35][11];
    ele[15][12] != ele[15][13];
    ele[15][12] != ele[15][14];
    ele[15][12] != ele[15][15];
    ele[15][12] != ele[15][16];
    ele[15][12] != ele[15][17];
    ele[15][12] != ele[15][18];
    ele[15][12] != ele[15][19];
    ele[15][12] != ele[15][20];
    ele[15][12] != ele[15][21];
    ele[15][12] != ele[15][22];
    ele[15][12] != ele[15][23];
    ele[15][12] != ele[15][24];
    ele[15][12] != ele[15][25];
    ele[15][12] != ele[15][26];
    ele[15][12] != ele[15][27];
    ele[15][12] != ele[15][28];
    ele[15][12] != ele[15][29];
    ele[15][12] != ele[15][30];
    ele[15][12] != ele[15][31];
    ele[15][12] != ele[15][32];
    ele[15][12] != ele[15][33];
    ele[15][12] != ele[15][34];
    ele[15][12] != ele[15][35];
    ele[15][12] != ele[16][12];
    ele[15][12] != ele[16][13];
    ele[15][12] != ele[16][14];
    ele[15][12] != ele[16][15];
    ele[15][12] != ele[16][16];
    ele[15][12] != ele[16][17];
    ele[15][12] != ele[17][12];
    ele[15][12] != ele[17][13];
    ele[15][12] != ele[17][14];
    ele[15][12] != ele[17][15];
    ele[15][12] != ele[17][16];
    ele[15][12] != ele[17][17];
    ele[15][12] != ele[18][12];
    ele[15][12] != ele[19][12];
    ele[15][12] != ele[20][12];
    ele[15][12] != ele[21][12];
    ele[15][12] != ele[22][12];
    ele[15][12] != ele[23][12];
    ele[15][12] != ele[24][12];
    ele[15][12] != ele[25][12];
    ele[15][12] != ele[26][12];
    ele[15][12] != ele[27][12];
    ele[15][12] != ele[28][12];
    ele[15][12] != ele[29][12];
    ele[15][12] != ele[30][12];
    ele[15][12] != ele[31][12];
    ele[15][12] != ele[32][12];
    ele[15][12] != ele[33][12];
    ele[15][12] != ele[34][12];
    ele[15][12] != ele[35][12];
    ele[15][13] != ele[15][14];
    ele[15][13] != ele[15][15];
    ele[15][13] != ele[15][16];
    ele[15][13] != ele[15][17];
    ele[15][13] != ele[15][18];
    ele[15][13] != ele[15][19];
    ele[15][13] != ele[15][20];
    ele[15][13] != ele[15][21];
    ele[15][13] != ele[15][22];
    ele[15][13] != ele[15][23];
    ele[15][13] != ele[15][24];
    ele[15][13] != ele[15][25];
    ele[15][13] != ele[15][26];
    ele[15][13] != ele[15][27];
    ele[15][13] != ele[15][28];
    ele[15][13] != ele[15][29];
    ele[15][13] != ele[15][30];
    ele[15][13] != ele[15][31];
    ele[15][13] != ele[15][32];
    ele[15][13] != ele[15][33];
    ele[15][13] != ele[15][34];
    ele[15][13] != ele[15][35];
    ele[15][13] != ele[16][12];
    ele[15][13] != ele[16][13];
    ele[15][13] != ele[16][14];
    ele[15][13] != ele[16][15];
    ele[15][13] != ele[16][16];
    ele[15][13] != ele[16][17];
    ele[15][13] != ele[17][12];
    ele[15][13] != ele[17][13];
    ele[15][13] != ele[17][14];
    ele[15][13] != ele[17][15];
    ele[15][13] != ele[17][16];
    ele[15][13] != ele[17][17];
    ele[15][13] != ele[18][13];
    ele[15][13] != ele[19][13];
    ele[15][13] != ele[20][13];
    ele[15][13] != ele[21][13];
    ele[15][13] != ele[22][13];
    ele[15][13] != ele[23][13];
    ele[15][13] != ele[24][13];
    ele[15][13] != ele[25][13];
    ele[15][13] != ele[26][13];
    ele[15][13] != ele[27][13];
    ele[15][13] != ele[28][13];
    ele[15][13] != ele[29][13];
    ele[15][13] != ele[30][13];
    ele[15][13] != ele[31][13];
    ele[15][13] != ele[32][13];
    ele[15][13] != ele[33][13];
    ele[15][13] != ele[34][13];
    ele[15][13] != ele[35][13];
    ele[15][14] != ele[15][15];
    ele[15][14] != ele[15][16];
    ele[15][14] != ele[15][17];
    ele[15][14] != ele[15][18];
    ele[15][14] != ele[15][19];
    ele[15][14] != ele[15][20];
    ele[15][14] != ele[15][21];
    ele[15][14] != ele[15][22];
    ele[15][14] != ele[15][23];
    ele[15][14] != ele[15][24];
    ele[15][14] != ele[15][25];
    ele[15][14] != ele[15][26];
    ele[15][14] != ele[15][27];
    ele[15][14] != ele[15][28];
    ele[15][14] != ele[15][29];
    ele[15][14] != ele[15][30];
    ele[15][14] != ele[15][31];
    ele[15][14] != ele[15][32];
    ele[15][14] != ele[15][33];
    ele[15][14] != ele[15][34];
    ele[15][14] != ele[15][35];
    ele[15][14] != ele[16][12];
    ele[15][14] != ele[16][13];
    ele[15][14] != ele[16][14];
    ele[15][14] != ele[16][15];
    ele[15][14] != ele[16][16];
    ele[15][14] != ele[16][17];
    ele[15][14] != ele[17][12];
    ele[15][14] != ele[17][13];
    ele[15][14] != ele[17][14];
    ele[15][14] != ele[17][15];
    ele[15][14] != ele[17][16];
    ele[15][14] != ele[17][17];
    ele[15][14] != ele[18][14];
    ele[15][14] != ele[19][14];
    ele[15][14] != ele[20][14];
    ele[15][14] != ele[21][14];
    ele[15][14] != ele[22][14];
    ele[15][14] != ele[23][14];
    ele[15][14] != ele[24][14];
    ele[15][14] != ele[25][14];
    ele[15][14] != ele[26][14];
    ele[15][14] != ele[27][14];
    ele[15][14] != ele[28][14];
    ele[15][14] != ele[29][14];
    ele[15][14] != ele[30][14];
    ele[15][14] != ele[31][14];
    ele[15][14] != ele[32][14];
    ele[15][14] != ele[33][14];
    ele[15][14] != ele[34][14];
    ele[15][14] != ele[35][14];
    ele[15][15] != ele[15][16];
    ele[15][15] != ele[15][17];
    ele[15][15] != ele[15][18];
    ele[15][15] != ele[15][19];
    ele[15][15] != ele[15][20];
    ele[15][15] != ele[15][21];
    ele[15][15] != ele[15][22];
    ele[15][15] != ele[15][23];
    ele[15][15] != ele[15][24];
    ele[15][15] != ele[15][25];
    ele[15][15] != ele[15][26];
    ele[15][15] != ele[15][27];
    ele[15][15] != ele[15][28];
    ele[15][15] != ele[15][29];
    ele[15][15] != ele[15][30];
    ele[15][15] != ele[15][31];
    ele[15][15] != ele[15][32];
    ele[15][15] != ele[15][33];
    ele[15][15] != ele[15][34];
    ele[15][15] != ele[15][35];
    ele[15][15] != ele[16][12];
    ele[15][15] != ele[16][13];
    ele[15][15] != ele[16][14];
    ele[15][15] != ele[16][15];
    ele[15][15] != ele[16][16];
    ele[15][15] != ele[16][17];
    ele[15][15] != ele[17][12];
    ele[15][15] != ele[17][13];
    ele[15][15] != ele[17][14];
    ele[15][15] != ele[17][15];
    ele[15][15] != ele[17][16];
    ele[15][15] != ele[17][17];
    ele[15][15] != ele[18][15];
    ele[15][15] != ele[19][15];
    ele[15][15] != ele[20][15];
    ele[15][15] != ele[21][15];
    ele[15][15] != ele[22][15];
    ele[15][15] != ele[23][15];
    ele[15][15] != ele[24][15];
    ele[15][15] != ele[25][15];
    ele[15][15] != ele[26][15];
    ele[15][15] != ele[27][15];
    ele[15][15] != ele[28][15];
    ele[15][15] != ele[29][15];
    ele[15][15] != ele[30][15];
    ele[15][15] != ele[31][15];
    ele[15][15] != ele[32][15];
    ele[15][15] != ele[33][15];
    ele[15][15] != ele[34][15];
    ele[15][15] != ele[35][15];
    ele[15][16] != ele[15][17];
    ele[15][16] != ele[15][18];
    ele[15][16] != ele[15][19];
    ele[15][16] != ele[15][20];
    ele[15][16] != ele[15][21];
    ele[15][16] != ele[15][22];
    ele[15][16] != ele[15][23];
    ele[15][16] != ele[15][24];
    ele[15][16] != ele[15][25];
    ele[15][16] != ele[15][26];
    ele[15][16] != ele[15][27];
    ele[15][16] != ele[15][28];
    ele[15][16] != ele[15][29];
    ele[15][16] != ele[15][30];
    ele[15][16] != ele[15][31];
    ele[15][16] != ele[15][32];
    ele[15][16] != ele[15][33];
    ele[15][16] != ele[15][34];
    ele[15][16] != ele[15][35];
    ele[15][16] != ele[16][12];
    ele[15][16] != ele[16][13];
    ele[15][16] != ele[16][14];
    ele[15][16] != ele[16][15];
    ele[15][16] != ele[16][16];
    ele[15][16] != ele[16][17];
    ele[15][16] != ele[17][12];
    ele[15][16] != ele[17][13];
    ele[15][16] != ele[17][14];
    ele[15][16] != ele[17][15];
    ele[15][16] != ele[17][16];
    ele[15][16] != ele[17][17];
    ele[15][16] != ele[18][16];
    ele[15][16] != ele[19][16];
    ele[15][16] != ele[20][16];
    ele[15][16] != ele[21][16];
    ele[15][16] != ele[22][16];
    ele[15][16] != ele[23][16];
    ele[15][16] != ele[24][16];
    ele[15][16] != ele[25][16];
    ele[15][16] != ele[26][16];
    ele[15][16] != ele[27][16];
    ele[15][16] != ele[28][16];
    ele[15][16] != ele[29][16];
    ele[15][16] != ele[30][16];
    ele[15][16] != ele[31][16];
    ele[15][16] != ele[32][16];
    ele[15][16] != ele[33][16];
    ele[15][16] != ele[34][16];
    ele[15][16] != ele[35][16];
    ele[15][17] != ele[15][18];
    ele[15][17] != ele[15][19];
    ele[15][17] != ele[15][20];
    ele[15][17] != ele[15][21];
    ele[15][17] != ele[15][22];
    ele[15][17] != ele[15][23];
    ele[15][17] != ele[15][24];
    ele[15][17] != ele[15][25];
    ele[15][17] != ele[15][26];
    ele[15][17] != ele[15][27];
    ele[15][17] != ele[15][28];
    ele[15][17] != ele[15][29];
    ele[15][17] != ele[15][30];
    ele[15][17] != ele[15][31];
    ele[15][17] != ele[15][32];
    ele[15][17] != ele[15][33];
    ele[15][17] != ele[15][34];
    ele[15][17] != ele[15][35];
    ele[15][17] != ele[16][12];
    ele[15][17] != ele[16][13];
    ele[15][17] != ele[16][14];
    ele[15][17] != ele[16][15];
    ele[15][17] != ele[16][16];
    ele[15][17] != ele[16][17];
    ele[15][17] != ele[17][12];
    ele[15][17] != ele[17][13];
    ele[15][17] != ele[17][14];
    ele[15][17] != ele[17][15];
    ele[15][17] != ele[17][16];
    ele[15][17] != ele[17][17];
    ele[15][17] != ele[18][17];
    ele[15][17] != ele[19][17];
    ele[15][17] != ele[20][17];
    ele[15][17] != ele[21][17];
    ele[15][17] != ele[22][17];
    ele[15][17] != ele[23][17];
    ele[15][17] != ele[24][17];
    ele[15][17] != ele[25][17];
    ele[15][17] != ele[26][17];
    ele[15][17] != ele[27][17];
    ele[15][17] != ele[28][17];
    ele[15][17] != ele[29][17];
    ele[15][17] != ele[30][17];
    ele[15][17] != ele[31][17];
    ele[15][17] != ele[32][17];
    ele[15][17] != ele[33][17];
    ele[15][17] != ele[34][17];
    ele[15][17] != ele[35][17];
    ele[15][18] != ele[15][19];
    ele[15][18] != ele[15][20];
    ele[15][18] != ele[15][21];
    ele[15][18] != ele[15][22];
    ele[15][18] != ele[15][23];
    ele[15][18] != ele[15][24];
    ele[15][18] != ele[15][25];
    ele[15][18] != ele[15][26];
    ele[15][18] != ele[15][27];
    ele[15][18] != ele[15][28];
    ele[15][18] != ele[15][29];
    ele[15][18] != ele[15][30];
    ele[15][18] != ele[15][31];
    ele[15][18] != ele[15][32];
    ele[15][18] != ele[15][33];
    ele[15][18] != ele[15][34];
    ele[15][18] != ele[15][35];
    ele[15][18] != ele[16][18];
    ele[15][18] != ele[16][19];
    ele[15][18] != ele[16][20];
    ele[15][18] != ele[16][21];
    ele[15][18] != ele[16][22];
    ele[15][18] != ele[16][23];
    ele[15][18] != ele[17][18];
    ele[15][18] != ele[17][19];
    ele[15][18] != ele[17][20];
    ele[15][18] != ele[17][21];
    ele[15][18] != ele[17][22];
    ele[15][18] != ele[17][23];
    ele[15][18] != ele[18][18];
    ele[15][18] != ele[19][18];
    ele[15][18] != ele[20][18];
    ele[15][18] != ele[21][18];
    ele[15][18] != ele[22][18];
    ele[15][18] != ele[23][18];
    ele[15][18] != ele[24][18];
    ele[15][18] != ele[25][18];
    ele[15][18] != ele[26][18];
    ele[15][18] != ele[27][18];
    ele[15][18] != ele[28][18];
    ele[15][18] != ele[29][18];
    ele[15][18] != ele[30][18];
    ele[15][18] != ele[31][18];
    ele[15][18] != ele[32][18];
    ele[15][18] != ele[33][18];
    ele[15][18] != ele[34][18];
    ele[15][18] != ele[35][18];
    ele[15][19] != ele[15][20];
    ele[15][19] != ele[15][21];
    ele[15][19] != ele[15][22];
    ele[15][19] != ele[15][23];
    ele[15][19] != ele[15][24];
    ele[15][19] != ele[15][25];
    ele[15][19] != ele[15][26];
    ele[15][19] != ele[15][27];
    ele[15][19] != ele[15][28];
    ele[15][19] != ele[15][29];
    ele[15][19] != ele[15][30];
    ele[15][19] != ele[15][31];
    ele[15][19] != ele[15][32];
    ele[15][19] != ele[15][33];
    ele[15][19] != ele[15][34];
    ele[15][19] != ele[15][35];
    ele[15][19] != ele[16][18];
    ele[15][19] != ele[16][19];
    ele[15][19] != ele[16][20];
    ele[15][19] != ele[16][21];
    ele[15][19] != ele[16][22];
    ele[15][19] != ele[16][23];
    ele[15][19] != ele[17][18];
    ele[15][19] != ele[17][19];
    ele[15][19] != ele[17][20];
    ele[15][19] != ele[17][21];
    ele[15][19] != ele[17][22];
    ele[15][19] != ele[17][23];
    ele[15][19] != ele[18][19];
    ele[15][19] != ele[19][19];
    ele[15][19] != ele[20][19];
    ele[15][19] != ele[21][19];
    ele[15][19] != ele[22][19];
    ele[15][19] != ele[23][19];
    ele[15][19] != ele[24][19];
    ele[15][19] != ele[25][19];
    ele[15][19] != ele[26][19];
    ele[15][19] != ele[27][19];
    ele[15][19] != ele[28][19];
    ele[15][19] != ele[29][19];
    ele[15][19] != ele[30][19];
    ele[15][19] != ele[31][19];
    ele[15][19] != ele[32][19];
    ele[15][19] != ele[33][19];
    ele[15][19] != ele[34][19];
    ele[15][19] != ele[35][19];
    ele[15][2] != ele[15][10];
    ele[15][2] != ele[15][11];
    ele[15][2] != ele[15][12];
    ele[15][2] != ele[15][13];
    ele[15][2] != ele[15][14];
    ele[15][2] != ele[15][15];
    ele[15][2] != ele[15][16];
    ele[15][2] != ele[15][17];
    ele[15][2] != ele[15][18];
    ele[15][2] != ele[15][19];
    ele[15][2] != ele[15][20];
    ele[15][2] != ele[15][21];
    ele[15][2] != ele[15][22];
    ele[15][2] != ele[15][23];
    ele[15][2] != ele[15][24];
    ele[15][2] != ele[15][25];
    ele[15][2] != ele[15][26];
    ele[15][2] != ele[15][27];
    ele[15][2] != ele[15][28];
    ele[15][2] != ele[15][29];
    ele[15][2] != ele[15][3];
    ele[15][2] != ele[15][30];
    ele[15][2] != ele[15][31];
    ele[15][2] != ele[15][32];
    ele[15][2] != ele[15][33];
    ele[15][2] != ele[15][34];
    ele[15][2] != ele[15][35];
    ele[15][2] != ele[15][4];
    ele[15][2] != ele[15][5];
    ele[15][2] != ele[15][6];
    ele[15][2] != ele[15][7];
    ele[15][2] != ele[15][8];
    ele[15][2] != ele[15][9];
    ele[15][2] != ele[16][0];
    ele[15][2] != ele[16][1];
    ele[15][2] != ele[16][2];
    ele[15][2] != ele[16][3];
    ele[15][2] != ele[16][4];
    ele[15][2] != ele[16][5];
    ele[15][2] != ele[17][0];
    ele[15][2] != ele[17][1];
    ele[15][2] != ele[17][2];
    ele[15][2] != ele[17][3];
    ele[15][2] != ele[17][4];
    ele[15][2] != ele[17][5];
    ele[15][2] != ele[18][2];
    ele[15][2] != ele[19][2];
    ele[15][2] != ele[20][2];
    ele[15][2] != ele[21][2];
    ele[15][2] != ele[22][2];
    ele[15][2] != ele[23][2];
    ele[15][2] != ele[24][2];
    ele[15][2] != ele[25][2];
    ele[15][2] != ele[26][2];
    ele[15][2] != ele[27][2];
    ele[15][2] != ele[28][2];
    ele[15][2] != ele[29][2];
    ele[15][2] != ele[30][2];
    ele[15][2] != ele[31][2];
    ele[15][2] != ele[32][2];
    ele[15][2] != ele[33][2];
    ele[15][2] != ele[34][2];
    ele[15][2] != ele[35][2];
    ele[15][20] != ele[15][21];
    ele[15][20] != ele[15][22];
    ele[15][20] != ele[15][23];
    ele[15][20] != ele[15][24];
    ele[15][20] != ele[15][25];
    ele[15][20] != ele[15][26];
    ele[15][20] != ele[15][27];
    ele[15][20] != ele[15][28];
    ele[15][20] != ele[15][29];
    ele[15][20] != ele[15][30];
    ele[15][20] != ele[15][31];
    ele[15][20] != ele[15][32];
    ele[15][20] != ele[15][33];
    ele[15][20] != ele[15][34];
    ele[15][20] != ele[15][35];
    ele[15][20] != ele[16][18];
    ele[15][20] != ele[16][19];
    ele[15][20] != ele[16][20];
    ele[15][20] != ele[16][21];
    ele[15][20] != ele[16][22];
    ele[15][20] != ele[16][23];
    ele[15][20] != ele[17][18];
    ele[15][20] != ele[17][19];
    ele[15][20] != ele[17][20];
    ele[15][20] != ele[17][21];
    ele[15][20] != ele[17][22];
    ele[15][20] != ele[17][23];
    ele[15][20] != ele[18][20];
    ele[15][20] != ele[19][20];
    ele[15][20] != ele[20][20];
    ele[15][20] != ele[21][20];
    ele[15][20] != ele[22][20];
    ele[15][20] != ele[23][20];
    ele[15][20] != ele[24][20];
    ele[15][20] != ele[25][20];
    ele[15][20] != ele[26][20];
    ele[15][20] != ele[27][20];
    ele[15][20] != ele[28][20];
    ele[15][20] != ele[29][20];
    ele[15][20] != ele[30][20];
    ele[15][20] != ele[31][20];
    ele[15][20] != ele[32][20];
    ele[15][20] != ele[33][20];
    ele[15][20] != ele[34][20];
    ele[15][20] != ele[35][20];
    ele[15][21] != ele[15][22];
    ele[15][21] != ele[15][23];
    ele[15][21] != ele[15][24];
    ele[15][21] != ele[15][25];
    ele[15][21] != ele[15][26];
    ele[15][21] != ele[15][27];
    ele[15][21] != ele[15][28];
    ele[15][21] != ele[15][29];
    ele[15][21] != ele[15][30];
    ele[15][21] != ele[15][31];
    ele[15][21] != ele[15][32];
    ele[15][21] != ele[15][33];
    ele[15][21] != ele[15][34];
    ele[15][21] != ele[15][35];
    ele[15][21] != ele[16][18];
    ele[15][21] != ele[16][19];
    ele[15][21] != ele[16][20];
    ele[15][21] != ele[16][21];
    ele[15][21] != ele[16][22];
    ele[15][21] != ele[16][23];
    ele[15][21] != ele[17][18];
    ele[15][21] != ele[17][19];
    ele[15][21] != ele[17][20];
    ele[15][21] != ele[17][21];
    ele[15][21] != ele[17][22];
    ele[15][21] != ele[17][23];
    ele[15][21] != ele[18][21];
    ele[15][21] != ele[19][21];
    ele[15][21] != ele[20][21];
    ele[15][21] != ele[21][21];
    ele[15][21] != ele[22][21];
    ele[15][21] != ele[23][21];
    ele[15][21] != ele[24][21];
    ele[15][21] != ele[25][21];
    ele[15][21] != ele[26][21];
    ele[15][21] != ele[27][21];
    ele[15][21] != ele[28][21];
    ele[15][21] != ele[29][21];
    ele[15][21] != ele[30][21];
    ele[15][21] != ele[31][21];
    ele[15][21] != ele[32][21];
    ele[15][21] != ele[33][21];
    ele[15][21] != ele[34][21];
    ele[15][21] != ele[35][21];
    ele[15][22] != ele[15][23];
    ele[15][22] != ele[15][24];
    ele[15][22] != ele[15][25];
    ele[15][22] != ele[15][26];
    ele[15][22] != ele[15][27];
    ele[15][22] != ele[15][28];
    ele[15][22] != ele[15][29];
    ele[15][22] != ele[15][30];
    ele[15][22] != ele[15][31];
    ele[15][22] != ele[15][32];
    ele[15][22] != ele[15][33];
    ele[15][22] != ele[15][34];
    ele[15][22] != ele[15][35];
    ele[15][22] != ele[16][18];
    ele[15][22] != ele[16][19];
    ele[15][22] != ele[16][20];
    ele[15][22] != ele[16][21];
    ele[15][22] != ele[16][22];
    ele[15][22] != ele[16][23];
    ele[15][22] != ele[17][18];
    ele[15][22] != ele[17][19];
    ele[15][22] != ele[17][20];
    ele[15][22] != ele[17][21];
    ele[15][22] != ele[17][22];
    ele[15][22] != ele[17][23];
    ele[15][22] != ele[18][22];
    ele[15][22] != ele[19][22];
    ele[15][22] != ele[20][22];
    ele[15][22] != ele[21][22];
    ele[15][22] != ele[22][22];
    ele[15][22] != ele[23][22];
    ele[15][22] != ele[24][22];
    ele[15][22] != ele[25][22];
    ele[15][22] != ele[26][22];
    ele[15][22] != ele[27][22];
    ele[15][22] != ele[28][22];
    ele[15][22] != ele[29][22];
    ele[15][22] != ele[30][22];
    ele[15][22] != ele[31][22];
    ele[15][22] != ele[32][22];
    ele[15][22] != ele[33][22];
    ele[15][22] != ele[34][22];
    ele[15][22] != ele[35][22];
    ele[15][23] != ele[15][24];
    ele[15][23] != ele[15][25];
    ele[15][23] != ele[15][26];
    ele[15][23] != ele[15][27];
    ele[15][23] != ele[15][28];
    ele[15][23] != ele[15][29];
    ele[15][23] != ele[15][30];
    ele[15][23] != ele[15][31];
    ele[15][23] != ele[15][32];
    ele[15][23] != ele[15][33];
    ele[15][23] != ele[15][34];
    ele[15][23] != ele[15][35];
    ele[15][23] != ele[16][18];
    ele[15][23] != ele[16][19];
    ele[15][23] != ele[16][20];
    ele[15][23] != ele[16][21];
    ele[15][23] != ele[16][22];
    ele[15][23] != ele[16][23];
    ele[15][23] != ele[17][18];
    ele[15][23] != ele[17][19];
    ele[15][23] != ele[17][20];
    ele[15][23] != ele[17][21];
    ele[15][23] != ele[17][22];
    ele[15][23] != ele[17][23];
    ele[15][23] != ele[18][23];
    ele[15][23] != ele[19][23];
    ele[15][23] != ele[20][23];
    ele[15][23] != ele[21][23];
    ele[15][23] != ele[22][23];
    ele[15][23] != ele[23][23];
    ele[15][23] != ele[24][23];
    ele[15][23] != ele[25][23];
    ele[15][23] != ele[26][23];
    ele[15][23] != ele[27][23];
    ele[15][23] != ele[28][23];
    ele[15][23] != ele[29][23];
    ele[15][23] != ele[30][23];
    ele[15][23] != ele[31][23];
    ele[15][23] != ele[32][23];
    ele[15][23] != ele[33][23];
    ele[15][23] != ele[34][23];
    ele[15][23] != ele[35][23];
    ele[15][24] != ele[15][25];
    ele[15][24] != ele[15][26];
    ele[15][24] != ele[15][27];
    ele[15][24] != ele[15][28];
    ele[15][24] != ele[15][29];
    ele[15][24] != ele[15][30];
    ele[15][24] != ele[15][31];
    ele[15][24] != ele[15][32];
    ele[15][24] != ele[15][33];
    ele[15][24] != ele[15][34];
    ele[15][24] != ele[15][35];
    ele[15][24] != ele[16][24];
    ele[15][24] != ele[16][25];
    ele[15][24] != ele[16][26];
    ele[15][24] != ele[16][27];
    ele[15][24] != ele[16][28];
    ele[15][24] != ele[16][29];
    ele[15][24] != ele[17][24];
    ele[15][24] != ele[17][25];
    ele[15][24] != ele[17][26];
    ele[15][24] != ele[17][27];
    ele[15][24] != ele[17][28];
    ele[15][24] != ele[17][29];
    ele[15][24] != ele[18][24];
    ele[15][24] != ele[19][24];
    ele[15][24] != ele[20][24];
    ele[15][24] != ele[21][24];
    ele[15][24] != ele[22][24];
    ele[15][24] != ele[23][24];
    ele[15][24] != ele[24][24];
    ele[15][24] != ele[25][24];
    ele[15][24] != ele[26][24];
    ele[15][24] != ele[27][24];
    ele[15][24] != ele[28][24];
    ele[15][24] != ele[29][24];
    ele[15][24] != ele[30][24];
    ele[15][24] != ele[31][24];
    ele[15][24] != ele[32][24];
    ele[15][24] != ele[33][24];
    ele[15][24] != ele[34][24];
    ele[15][24] != ele[35][24];
    ele[15][25] != ele[15][26];
    ele[15][25] != ele[15][27];
    ele[15][25] != ele[15][28];
    ele[15][25] != ele[15][29];
    ele[15][25] != ele[15][30];
    ele[15][25] != ele[15][31];
    ele[15][25] != ele[15][32];
    ele[15][25] != ele[15][33];
    ele[15][25] != ele[15][34];
    ele[15][25] != ele[15][35];
    ele[15][25] != ele[16][24];
    ele[15][25] != ele[16][25];
    ele[15][25] != ele[16][26];
    ele[15][25] != ele[16][27];
    ele[15][25] != ele[16][28];
    ele[15][25] != ele[16][29];
    ele[15][25] != ele[17][24];
    ele[15][25] != ele[17][25];
    ele[15][25] != ele[17][26];
    ele[15][25] != ele[17][27];
    ele[15][25] != ele[17][28];
    ele[15][25] != ele[17][29];
    ele[15][25] != ele[18][25];
    ele[15][25] != ele[19][25];
    ele[15][25] != ele[20][25];
    ele[15][25] != ele[21][25];
    ele[15][25] != ele[22][25];
    ele[15][25] != ele[23][25];
    ele[15][25] != ele[24][25];
    ele[15][25] != ele[25][25];
    ele[15][25] != ele[26][25];
    ele[15][25] != ele[27][25];
    ele[15][25] != ele[28][25];
    ele[15][25] != ele[29][25];
    ele[15][25] != ele[30][25];
    ele[15][25] != ele[31][25];
    ele[15][25] != ele[32][25];
    ele[15][25] != ele[33][25];
    ele[15][25] != ele[34][25];
    ele[15][25] != ele[35][25];
    ele[15][26] != ele[15][27];
    ele[15][26] != ele[15][28];
    ele[15][26] != ele[15][29];
    ele[15][26] != ele[15][30];
    ele[15][26] != ele[15][31];
    ele[15][26] != ele[15][32];
    ele[15][26] != ele[15][33];
    ele[15][26] != ele[15][34];
    ele[15][26] != ele[15][35];
    ele[15][26] != ele[16][24];
    ele[15][26] != ele[16][25];
    ele[15][26] != ele[16][26];
    ele[15][26] != ele[16][27];
    ele[15][26] != ele[16][28];
    ele[15][26] != ele[16][29];
    ele[15][26] != ele[17][24];
    ele[15][26] != ele[17][25];
    ele[15][26] != ele[17][26];
    ele[15][26] != ele[17][27];
    ele[15][26] != ele[17][28];
    ele[15][26] != ele[17][29];
    ele[15][26] != ele[18][26];
    ele[15][26] != ele[19][26];
    ele[15][26] != ele[20][26];
    ele[15][26] != ele[21][26];
    ele[15][26] != ele[22][26];
    ele[15][26] != ele[23][26];
    ele[15][26] != ele[24][26];
    ele[15][26] != ele[25][26];
    ele[15][26] != ele[26][26];
    ele[15][26] != ele[27][26];
    ele[15][26] != ele[28][26];
    ele[15][26] != ele[29][26];
    ele[15][26] != ele[30][26];
    ele[15][26] != ele[31][26];
    ele[15][26] != ele[32][26];
    ele[15][26] != ele[33][26];
    ele[15][26] != ele[34][26];
    ele[15][26] != ele[35][26];
    ele[15][27] != ele[15][28];
    ele[15][27] != ele[15][29];
    ele[15][27] != ele[15][30];
    ele[15][27] != ele[15][31];
    ele[15][27] != ele[15][32];
    ele[15][27] != ele[15][33];
    ele[15][27] != ele[15][34];
    ele[15][27] != ele[15][35];
    ele[15][27] != ele[16][24];
    ele[15][27] != ele[16][25];
    ele[15][27] != ele[16][26];
    ele[15][27] != ele[16][27];
    ele[15][27] != ele[16][28];
    ele[15][27] != ele[16][29];
    ele[15][27] != ele[17][24];
    ele[15][27] != ele[17][25];
    ele[15][27] != ele[17][26];
    ele[15][27] != ele[17][27];
    ele[15][27] != ele[17][28];
    ele[15][27] != ele[17][29];
    ele[15][27] != ele[18][27];
    ele[15][27] != ele[19][27];
    ele[15][27] != ele[20][27];
    ele[15][27] != ele[21][27];
    ele[15][27] != ele[22][27];
    ele[15][27] != ele[23][27];
    ele[15][27] != ele[24][27];
    ele[15][27] != ele[25][27];
    ele[15][27] != ele[26][27];
    ele[15][27] != ele[27][27];
    ele[15][27] != ele[28][27];
    ele[15][27] != ele[29][27];
    ele[15][27] != ele[30][27];
    ele[15][27] != ele[31][27];
    ele[15][27] != ele[32][27];
    ele[15][27] != ele[33][27];
    ele[15][27] != ele[34][27];
    ele[15][27] != ele[35][27];
    ele[15][28] != ele[15][29];
    ele[15][28] != ele[15][30];
    ele[15][28] != ele[15][31];
    ele[15][28] != ele[15][32];
    ele[15][28] != ele[15][33];
    ele[15][28] != ele[15][34];
    ele[15][28] != ele[15][35];
    ele[15][28] != ele[16][24];
    ele[15][28] != ele[16][25];
    ele[15][28] != ele[16][26];
    ele[15][28] != ele[16][27];
    ele[15][28] != ele[16][28];
    ele[15][28] != ele[16][29];
    ele[15][28] != ele[17][24];
    ele[15][28] != ele[17][25];
    ele[15][28] != ele[17][26];
    ele[15][28] != ele[17][27];
    ele[15][28] != ele[17][28];
    ele[15][28] != ele[17][29];
    ele[15][28] != ele[18][28];
    ele[15][28] != ele[19][28];
    ele[15][28] != ele[20][28];
    ele[15][28] != ele[21][28];
    ele[15][28] != ele[22][28];
    ele[15][28] != ele[23][28];
    ele[15][28] != ele[24][28];
    ele[15][28] != ele[25][28];
    ele[15][28] != ele[26][28];
    ele[15][28] != ele[27][28];
    ele[15][28] != ele[28][28];
    ele[15][28] != ele[29][28];
    ele[15][28] != ele[30][28];
    ele[15][28] != ele[31][28];
    ele[15][28] != ele[32][28];
    ele[15][28] != ele[33][28];
    ele[15][28] != ele[34][28];
    ele[15][28] != ele[35][28];
    ele[15][29] != ele[15][30];
    ele[15][29] != ele[15][31];
    ele[15][29] != ele[15][32];
    ele[15][29] != ele[15][33];
    ele[15][29] != ele[15][34];
    ele[15][29] != ele[15][35];
    ele[15][29] != ele[16][24];
    ele[15][29] != ele[16][25];
    ele[15][29] != ele[16][26];
    ele[15][29] != ele[16][27];
    ele[15][29] != ele[16][28];
    ele[15][29] != ele[16][29];
    ele[15][29] != ele[17][24];
    ele[15][29] != ele[17][25];
    ele[15][29] != ele[17][26];
    ele[15][29] != ele[17][27];
    ele[15][29] != ele[17][28];
    ele[15][29] != ele[17][29];
    ele[15][29] != ele[18][29];
    ele[15][29] != ele[19][29];
    ele[15][29] != ele[20][29];
    ele[15][29] != ele[21][29];
    ele[15][29] != ele[22][29];
    ele[15][29] != ele[23][29];
    ele[15][29] != ele[24][29];
    ele[15][29] != ele[25][29];
    ele[15][29] != ele[26][29];
    ele[15][29] != ele[27][29];
    ele[15][29] != ele[28][29];
    ele[15][29] != ele[29][29];
    ele[15][29] != ele[30][29];
    ele[15][29] != ele[31][29];
    ele[15][29] != ele[32][29];
    ele[15][29] != ele[33][29];
    ele[15][29] != ele[34][29];
    ele[15][29] != ele[35][29];
    ele[15][3] != ele[15][10];
    ele[15][3] != ele[15][11];
    ele[15][3] != ele[15][12];
    ele[15][3] != ele[15][13];
    ele[15][3] != ele[15][14];
    ele[15][3] != ele[15][15];
    ele[15][3] != ele[15][16];
    ele[15][3] != ele[15][17];
    ele[15][3] != ele[15][18];
    ele[15][3] != ele[15][19];
    ele[15][3] != ele[15][20];
    ele[15][3] != ele[15][21];
    ele[15][3] != ele[15][22];
    ele[15][3] != ele[15][23];
    ele[15][3] != ele[15][24];
    ele[15][3] != ele[15][25];
    ele[15][3] != ele[15][26];
    ele[15][3] != ele[15][27];
    ele[15][3] != ele[15][28];
    ele[15][3] != ele[15][29];
    ele[15][3] != ele[15][30];
    ele[15][3] != ele[15][31];
    ele[15][3] != ele[15][32];
    ele[15][3] != ele[15][33];
    ele[15][3] != ele[15][34];
    ele[15][3] != ele[15][35];
    ele[15][3] != ele[15][4];
    ele[15][3] != ele[15][5];
    ele[15][3] != ele[15][6];
    ele[15][3] != ele[15][7];
    ele[15][3] != ele[15][8];
    ele[15][3] != ele[15][9];
    ele[15][3] != ele[16][0];
    ele[15][3] != ele[16][1];
    ele[15][3] != ele[16][2];
    ele[15][3] != ele[16][3];
    ele[15][3] != ele[16][4];
    ele[15][3] != ele[16][5];
    ele[15][3] != ele[17][0];
    ele[15][3] != ele[17][1];
    ele[15][3] != ele[17][2];
    ele[15][3] != ele[17][3];
    ele[15][3] != ele[17][4];
    ele[15][3] != ele[17][5];
    ele[15][3] != ele[18][3];
    ele[15][3] != ele[19][3];
    ele[15][3] != ele[20][3];
    ele[15][3] != ele[21][3];
    ele[15][3] != ele[22][3];
    ele[15][3] != ele[23][3];
    ele[15][3] != ele[24][3];
    ele[15][3] != ele[25][3];
    ele[15][3] != ele[26][3];
    ele[15][3] != ele[27][3];
    ele[15][3] != ele[28][3];
    ele[15][3] != ele[29][3];
    ele[15][3] != ele[30][3];
    ele[15][3] != ele[31][3];
    ele[15][3] != ele[32][3];
    ele[15][3] != ele[33][3];
    ele[15][3] != ele[34][3];
    ele[15][3] != ele[35][3];
    ele[15][30] != ele[15][31];
    ele[15][30] != ele[15][32];
    ele[15][30] != ele[15][33];
    ele[15][30] != ele[15][34];
    ele[15][30] != ele[15][35];
    ele[15][30] != ele[16][30];
    ele[15][30] != ele[16][31];
    ele[15][30] != ele[16][32];
    ele[15][30] != ele[16][33];
    ele[15][30] != ele[16][34];
    ele[15][30] != ele[16][35];
    ele[15][30] != ele[17][30];
    ele[15][30] != ele[17][31];
    ele[15][30] != ele[17][32];
    ele[15][30] != ele[17][33];
    ele[15][30] != ele[17][34];
    ele[15][30] != ele[17][35];
    ele[15][30] != ele[18][30];
    ele[15][30] != ele[19][30];
    ele[15][30] != ele[20][30];
    ele[15][30] != ele[21][30];
    ele[15][30] != ele[22][30];
    ele[15][30] != ele[23][30];
    ele[15][30] != ele[24][30];
    ele[15][30] != ele[25][30];
    ele[15][30] != ele[26][30];
    ele[15][30] != ele[27][30];
    ele[15][30] != ele[28][30];
    ele[15][30] != ele[29][30];
    ele[15][30] != ele[30][30];
    ele[15][30] != ele[31][30];
    ele[15][30] != ele[32][30];
    ele[15][30] != ele[33][30];
    ele[15][30] != ele[34][30];
    ele[15][30] != ele[35][30];
    ele[15][31] != ele[15][32];
    ele[15][31] != ele[15][33];
    ele[15][31] != ele[15][34];
    ele[15][31] != ele[15][35];
    ele[15][31] != ele[16][30];
    ele[15][31] != ele[16][31];
    ele[15][31] != ele[16][32];
    ele[15][31] != ele[16][33];
    ele[15][31] != ele[16][34];
    ele[15][31] != ele[16][35];
    ele[15][31] != ele[17][30];
    ele[15][31] != ele[17][31];
    ele[15][31] != ele[17][32];
    ele[15][31] != ele[17][33];
    ele[15][31] != ele[17][34];
    ele[15][31] != ele[17][35];
    ele[15][31] != ele[18][31];
    ele[15][31] != ele[19][31];
    ele[15][31] != ele[20][31];
    ele[15][31] != ele[21][31];
    ele[15][31] != ele[22][31];
    ele[15][31] != ele[23][31];
    ele[15][31] != ele[24][31];
    ele[15][31] != ele[25][31];
    ele[15][31] != ele[26][31];
    ele[15][31] != ele[27][31];
    ele[15][31] != ele[28][31];
    ele[15][31] != ele[29][31];
    ele[15][31] != ele[30][31];
    ele[15][31] != ele[31][31];
    ele[15][31] != ele[32][31];
    ele[15][31] != ele[33][31];
    ele[15][31] != ele[34][31];
    ele[15][31] != ele[35][31];
    ele[15][32] != ele[15][33];
    ele[15][32] != ele[15][34];
    ele[15][32] != ele[15][35];
    ele[15][32] != ele[16][30];
    ele[15][32] != ele[16][31];
    ele[15][32] != ele[16][32];
    ele[15][32] != ele[16][33];
    ele[15][32] != ele[16][34];
    ele[15][32] != ele[16][35];
    ele[15][32] != ele[17][30];
    ele[15][32] != ele[17][31];
    ele[15][32] != ele[17][32];
    ele[15][32] != ele[17][33];
    ele[15][32] != ele[17][34];
    ele[15][32] != ele[17][35];
    ele[15][32] != ele[18][32];
    ele[15][32] != ele[19][32];
    ele[15][32] != ele[20][32];
    ele[15][32] != ele[21][32];
    ele[15][32] != ele[22][32];
    ele[15][32] != ele[23][32];
    ele[15][32] != ele[24][32];
    ele[15][32] != ele[25][32];
    ele[15][32] != ele[26][32];
    ele[15][32] != ele[27][32];
    ele[15][32] != ele[28][32];
    ele[15][32] != ele[29][32];
    ele[15][32] != ele[30][32];
    ele[15][32] != ele[31][32];
    ele[15][32] != ele[32][32];
    ele[15][32] != ele[33][32];
    ele[15][32] != ele[34][32];
    ele[15][32] != ele[35][32];
    ele[15][33] != ele[15][34];
    ele[15][33] != ele[15][35];
    ele[15][33] != ele[16][30];
    ele[15][33] != ele[16][31];
    ele[15][33] != ele[16][32];
    ele[15][33] != ele[16][33];
    ele[15][33] != ele[16][34];
    ele[15][33] != ele[16][35];
    ele[15][33] != ele[17][30];
    ele[15][33] != ele[17][31];
    ele[15][33] != ele[17][32];
    ele[15][33] != ele[17][33];
    ele[15][33] != ele[17][34];
    ele[15][33] != ele[17][35];
    ele[15][33] != ele[18][33];
    ele[15][33] != ele[19][33];
    ele[15][33] != ele[20][33];
    ele[15][33] != ele[21][33];
    ele[15][33] != ele[22][33];
    ele[15][33] != ele[23][33];
    ele[15][33] != ele[24][33];
    ele[15][33] != ele[25][33];
    ele[15][33] != ele[26][33];
    ele[15][33] != ele[27][33];
    ele[15][33] != ele[28][33];
    ele[15][33] != ele[29][33];
    ele[15][33] != ele[30][33];
    ele[15][33] != ele[31][33];
    ele[15][33] != ele[32][33];
    ele[15][33] != ele[33][33];
    ele[15][33] != ele[34][33];
    ele[15][33] != ele[35][33];
    ele[15][34] != ele[15][35];
    ele[15][34] != ele[16][30];
    ele[15][34] != ele[16][31];
    ele[15][34] != ele[16][32];
    ele[15][34] != ele[16][33];
    ele[15][34] != ele[16][34];
    ele[15][34] != ele[16][35];
    ele[15][34] != ele[17][30];
    ele[15][34] != ele[17][31];
    ele[15][34] != ele[17][32];
    ele[15][34] != ele[17][33];
    ele[15][34] != ele[17][34];
    ele[15][34] != ele[17][35];
    ele[15][34] != ele[18][34];
    ele[15][34] != ele[19][34];
    ele[15][34] != ele[20][34];
    ele[15][34] != ele[21][34];
    ele[15][34] != ele[22][34];
    ele[15][34] != ele[23][34];
    ele[15][34] != ele[24][34];
    ele[15][34] != ele[25][34];
    ele[15][34] != ele[26][34];
    ele[15][34] != ele[27][34];
    ele[15][34] != ele[28][34];
    ele[15][34] != ele[29][34];
    ele[15][34] != ele[30][34];
    ele[15][34] != ele[31][34];
    ele[15][34] != ele[32][34];
    ele[15][34] != ele[33][34];
    ele[15][34] != ele[34][34];
    ele[15][34] != ele[35][34];
    ele[15][35] != ele[16][30];
    ele[15][35] != ele[16][31];
    ele[15][35] != ele[16][32];
    ele[15][35] != ele[16][33];
    ele[15][35] != ele[16][34];
    ele[15][35] != ele[16][35];
    ele[15][35] != ele[17][30];
    ele[15][35] != ele[17][31];
    ele[15][35] != ele[17][32];
    ele[15][35] != ele[17][33];
    ele[15][35] != ele[17][34];
    ele[15][35] != ele[17][35];
    ele[15][35] != ele[18][35];
    ele[15][35] != ele[19][35];
    ele[15][35] != ele[20][35];
    ele[15][35] != ele[21][35];
    ele[15][35] != ele[22][35];
    ele[15][35] != ele[23][35];
    ele[15][35] != ele[24][35];
    ele[15][35] != ele[25][35];
    ele[15][35] != ele[26][35];
    ele[15][35] != ele[27][35];
    ele[15][35] != ele[28][35];
    ele[15][35] != ele[29][35];
    ele[15][35] != ele[30][35];
    ele[15][35] != ele[31][35];
    ele[15][35] != ele[32][35];
    ele[15][35] != ele[33][35];
    ele[15][35] != ele[34][35];
    ele[15][35] != ele[35][35];
    ele[15][4] != ele[15][10];
    ele[15][4] != ele[15][11];
    ele[15][4] != ele[15][12];
    ele[15][4] != ele[15][13];
    ele[15][4] != ele[15][14];
    ele[15][4] != ele[15][15];
    ele[15][4] != ele[15][16];
    ele[15][4] != ele[15][17];
    ele[15][4] != ele[15][18];
    ele[15][4] != ele[15][19];
    ele[15][4] != ele[15][20];
    ele[15][4] != ele[15][21];
    ele[15][4] != ele[15][22];
    ele[15][4] != ele[15][23];
    ele[15][4] != ele[15][24];
    ele[15][4] != ele[15][25];
    ele[15][4] != ele[15][26];
    ele[15][4] != ele[15][27];
    ele[15][4] != ele[15][28];
    ele[15][4] != ele[15][29];
    ele[15][4] != ele[15][30];
    ele[15][4] != ele[15][31];
    ele[15][4] != ele[15][32];
    ele[15][4] != ele[15][33];
    ele[15][4] != ele[15][34];
    ele[15][4] != ele[15][35];
    ele[15][4] != ele[15][5];
    ele[15][4] != ele[15][6];
    ele[15][4] != ele[15][7];
    ele[15][4] != ele[15][8];
    ele[15][4] != ele[15][9];
    ele[15][4] != ele[16][0];
    ele[15][4] != ele[16][1];
    ele[15][4] != ele[16][2];
    ele[15][4] != ele[16][3];
    ele[15][4] != ele[16][4];
    ele[15][4] != ele[16][5];
    ele[15][4] != ele[17][0];
    ele[15][4] != ele[17][1];
    ele[15][4] != ele[17][2];
    ele[15][4] != ele[17][3];
    ele[15][4] != ele[17][4];
    ele[15][4] != ele[17][5];
    ele[15][4] != ele[18][4];
    ele[15][4] != ele[19][4];
    ele[15][4] != ele[20][4];
    ele[15][4] != ele[21][4];
    ele[15][4] != ele[22][4];
    ele[15][4] != ele[23][4];
    ele[15][4] != ele[24][4];
    ele[15][4] != ele[25][4];
    ele[15][4] != ele[26][4];
    ele[15][4] != ele[27][4];
    ele[15][4] != ele[28][4];
    ele[15][4] != ele[29][4];
    ele[15][4] != ele[30][4];
    ele[15][4] != ele[31][4];
    ele[15][4] != ele[32][4];
    ele[15][4] != ele[33][4];
    ele[15][4] != ele[34][4];
    ele[15][4] != ele[35][4];
    ele[15][5] != ele[15][10];
    ele[15][5] != ele[15][11];
    ele[15][5] != ele[15][12];
    ele[15][5] != ele[15][13];
    ele[15][5] != ele[15][14];
    ele[15][5] != ele[15][15];
    ele[15][5] != ele[15][16];
    ele[15][5] != ele[15][17];
    ele[15][5] != ele[15][18];
    ele[15][5] != ele[15][19];
    ele[15][5] != ele[15][20];
    ele[15][5] != ele[15][21];
    ele[15][5] != ele[15][22];
    ele[15][5] != ele[15][23];
    ele[15][5] != ele[15][24];
    ele[15][5] != ele[15][25];
    ele[15][5] != ele[15][26];
    ele[15][5] != ele[15][27];
    ele[15][5] != ele[15][28];
    ele[15][5] != ele[15][29];
    ele[15][5] != ele[15][30];
    ele[15][5] != ele[15][31];
    ele[15][5] != ele[15][32];
    ele[15][5] != ele[15][33];
    ele[15][5] != ele[15][34];
    ele[15][5] != ele[15][35];
    ele[15][5] != ele[15][6];
    ele[15][5] != ele[15][7];
    ele[15][5] != ele[15][8];
    ele[15][5] != ele[15][9];
    ele[15][5] != ele[16][0];
    ele[15][5] != ele[16][1];
    ele[15][5] != ele[16][2];
    ele[15][5] != ele[16][3];
    ele[15][5] != ele[16][4];
    ele[15][5] != ele[16][5];
    ele[15][5] != ele[17][0];
    ele[15][5] != ele[17][1];
    ele[15][5] != ele[17][2];
    ele[15][5] != ele[17][3];
    ele[15][5] != ele[17][4];
    ele[15][5] != ele[17][5];
    ele[15][5] != ele[18][5];
    ele[15][5] != ele[19][5];
    ele[15][5] != ele[20][5];
    ele[15][5] != ele[21][5];
    ele[15][5] != ele[22][5];
    ele[15][5] != ele[23][5];
    ele[15][5] != ele[24][5];
    ele[15][5] != ele[25][5];
    ele[15][5] != ele[26][5];
    ele[15][5] != ele[27][5];
    ele[15][5] != ele[28][5];
    ele[15][5] != ele[29][5];
    ele[15][5] != ele[30][5];
    ele[15][5] != ele[31][5];
    ele[15][5] != ele[32][5];
    ele[15][5] != ele[33][5];
    ele[15][5] != ele[34][5];
    ele[15][5] != ele[35][5];
    ele[15][6] != ele[15][10];
    ele[15][6] != ele[15][11];
    ele[15][6] != ele[15][12];
    ele[15][6] != ele[15][13];
    ele[15][6] != ele[15][14];
    ele[15][6] != ele[15][15];
    ele[15][6] != ele[15][16];
    ele[15][6] != ele[15][17];
    ele[15][6] != ele[15][18];
    ele[15][6] != ele[15][19];
    ele[15][6] != ele[15][20];
    ele[15][6] != ele[15][21];
    ele[15][6] != ele[15][22];
    ele[15][6] != ele[15][23];
    ele[15][6] != ele[15][24];
    ele[15][6] != ele[15][25];
    ele[15][6] != ele[15][26];
    ele[15][6] != ele[15][27];
    ele[15][6] != ele[15][28];
    ele[15][6] != ele[15][29];
    ele[15][6] != ele[15][30];
    ele[15][6] != ele[15][31];
    ele[15][6] != ele[15][32];
    ele[15][6] != ele[15][33];
    ele[15][6] != ele[15][34];
    ele[15][6] != ele[15][35];
    ele[15][6] != ele[15][7];
    ele[15][6] != ele[15][8];
    ele[15][6] != ele[15][9];
    ele[15][6] != ele[16][10];
    ele[15][6] != ele[16][11];
    ele[15][6] != ele[16][6];
    ele[15][6] != ele[16][7];
    ele[15][6] != ele[16][8];
    ele[15][6] != ele[16][9];
    ele[15][6] != ele[17][10];
    ele[15][6] != ele[17][11];
    ele[15][6] != ele[17][6];
    ele[15][6] != ele[17][7];
    ele[15][6] != ele[17][8];
    ele[15][6] != ele[17][9];
    ele[15][6] != ele[18][6];
    ele[15][6] != ele[19][6];
    ele[15][6] != ele[20][6];
    ele[15][6] != ele[21][6];
    ele[15][6] != ele[22][6];
    ele[15][6] != ele[23][6];
    ele[15][6] != ele[24][6];
    ele[15][6] != ele[25][6];
    ele[15][6] != ele[26][6];
    ele[15][6] != ele[27][6];
    ele[15][6] != ele[28][6];
    ele[15][6] != ele[29][6];
    ele[15][6] != ele[30][6];
    ele[15][6] != ele[31][6];
    ele[15][6] != ele[32][6];
    ele[15][6] != ele[33][6];
    ele[15][6] != ele[34][6];
    ele[15][6] != ele[35][6];
    ele[15][7] != ele[15][10];
    ele[15][7] != ele[15][11];
    ele[15][7] != ele[15][12];
    ele[15][7] != ele[15][13];
    ele[15][7] != ele[15][14];
    ele[15][7] != ele[15][15];
    ele[15][7] != ele[15][16];
    ele[15][7] != ele[15][17];
    ele[15][7] != ele[15][18];
    ele[15][7] != ele[15][19];
    ele[15][7] != ele[15][20];
    ele[15][7] != ele[15][21];
    ele[15][7] != ele[15][22];
    ele[15][7] != ele[15][23];
    ele[15][7] != ele[15][24];
    ele[15][7] != ele[15][25];
    ele[15][7] != ele[15][26];
    ele[15][7] != ele[15][27];
    ele[15][7] != ele[15][28];
    ele[15][7] != ele[15][29];
    ele[15][7] != ele[15][30];
    ele[15][7] != ele[15][31];
    ele[15][7] != ele[15][32];
    ele[15][7] != ele[15][33];
    ele[15][7] != ele[15][34];
    ele[15][7] != ele[15][35];
    ele[15][7] != ele[15][8];
    ele[15][7] != ele[15][9];
    ele[15][7] != ele[16][10];
    ele[15][7] != ele[16][11];
    ele[15][7] != ele[16][6];
    ele[15][7] != ele[16][7];
    ele[15][7] != ele[16][8];
    ele[15][7] != ele[16][9];
    ele[15][7] != ele[17][10];
    ele[15][7] != ele[17][11];
    ele[15][7] != ele[17][6];
    ele[15][7] != ele[17][7];
    ele[15][7] != ele[17][8];
    ele[15][7] != ele[17][9];
    ele[15][7] != ele[18][7];
    ele[15][7] != ele[19][7];
    ele[15][7] != ele[20][7];
    ele[15][7] != ele[21][7];
    ele[15][7] != ele[22][7];
    ele[15][7] != ele[23][7];
    ele[15][7] != ele[24][7];
    ele[15][7] != ele[25][7];
    ele[15][7] != ele[26][7];
    ele[15][7] != ele[27][7];
    ele[15][7] != ele[28][7];
    ele[15][7] != ele[29][7];
    ele[15][7] != ele[30][7];
    ele[15][7] != ele[31][7];
    ele[15][7] != ele[32][7];
    ele[15][7] != ele[33][7];
    ele[15][7] != ele[34][7];
    ele[15][7] != ele[35][7];
    ele[15][8] != ele[15][10];
    ele[15][8] != ele[15][11];
    ele[15][8] != ele[15][12];
    ele[15][8] != ele[15][13];
    ele[15][8] != ele[15][14];
    ele[15][8] != ele[15][15];
    ele[15][8] != ele[15][16];
    ele[15][8] != ele[15][17];
    ele[15][8] != ele[15][18];
    ele[15][8] != ele[15][19];
    ele[15][8] != ele[15][20];
    ele[15][8] != ele[15][21];
    ele[15][8] != ele[15][22];
    ele[15][8] != ele[15][23];
    ele[15][8] != ele[15][24];
    ele[15][8] != ele[15][25];
    ele[15][8] != ele[15][26];
    ele[15][8] != ele[15][27];
    ele[15][8] != ele[15][28];
    ele[15][8] != ele[15][29];
    ele[15][8] != ele[15][30];
    ele[15][8] != ele[15][31];
    ele[15][8] != ele[15][32];
    ele[15][8] != ele[15][33];
    ele[15][8] != ele[15][34];
    ele[15][8] != ele[15][35];
    ele[15][8] != ele[15][9];
    ele[15][8] != ele[16][10];
    ele[15][8] != ele[16][11];
    ele[15][8] != ele[16][6];
    ele[15][8] != ele[16][7];
    ele[15][8] != ele[16][8];
    ele[15][8] != ele[16][9];
    ele[15][8] != ele[17][10];
    ele[15][8] != ele[17][11];
    ele[15][8] != ele[17][6];
    ele[15][8] != ele[17][7];
    ele[15][8] != ele[17][8];
    ele[15][8] != ele[17][9];
    ele[15][8] != ele[18][8];
    ele[15][8] != ele[19][8];
    ele[15][8] != ele[20][8];
    ele[15][8] != ele[21][8];
    ele[15][8] != ele[22][8];
    ele[15][8] != ele[23][8];
    ele[15][8] != ele[24][8];
    ele[15][8] != ele[25][8];
    ele[15][8] != ele[26][8];
    ele[15][8] != ele[27][8];
    ele[15][8] != ele[28][8];
    ele[15][8] != ele[29][8];
    ele[15][8] != ele[30][8];
    ele[15][8] != ele[31][8];
    ele[15][8] != ele[32][8];
    ele[15][8] != ele[33][8];
    ele[15][8] != ele[34][8];
    ele[15][8] != ele[35][8];
    ele[15][9] != ele[15][10];
    ele[15][9] != ele[15][11];
    ele[15][9] != ele[15][12];
    ele[15][9] != ele[15][13];
    ele[15][9] != ele[15][14];
    ele[15][9] != ele[15][15];
    ele[15][9] != ele[15][16];
    ele[15][9] != ele[15][17];
    ele[15][9] != ele[15][18];
    ele[15][9] != ele[15][19];
    ele[15][9] != ele[15][20];
    ele[15][9] != ele[15][21];
    ele[15][9] != ele[15][22];
    ele[15][9] != ele[15][23];
    ele[15][9] != ele[15][24];
    ele[15][9] != ele[15][25];
    ele[15][9] != ele[15][26];
    ele[15][9] != ele[15][27];
    ele[15][9] != ele[15][28];
    ele[15][9] != ele[15][29];
    ele[15][9] != ele[15][30];
    ele[15][9] != ele[15][31];
    ele[15][9] != ele[15][32];
    ele[15][9] != ele[15][33];
    ele[15][9] != ele[15][34];
    ele[15][9] != ele[15][35];
    ele[15][9] != ele[16][10];
    ele[15][9] != ele[16][11];
    ele[15][9] != ele[16][6];
    ele[15][9] != ele[16][7];
    ele[15][9] != ele[16][8];
    ele[15][9] != ele[16][9];
    ele[15][9] != ele[17][10];
    ele[15][9] != ele[17][11];
    ele[15][9] != ele[17][6];
    ele[15][9] != ele[17][7];
    ele[15][9] != ele[17][8];
    ele[15][9] != ele[17][9];
    ele[15][9] != ele[18][9];
    ele[15][9] != ele[19][9];
    ele[15][9] != ele[20][9];
    ele[15][9] != ele[21][9];
    ele[15][9] != ele[22][9];
    ele[15][9] != ele[23][9];
    ele[15][9] != ele[24][9];
    ele[15][9] != ele[25][9];
    ele[15][9] != ele[26][9];
    ele[15][9] != ele[27][9];
    ele[15][9] != ele[28][9];
    ele[15][9] != ele[29][9];
    ele[15][9] != ele[30][9];
    ele[15][9] != ele[31][9];
    ele[15][9] != ele[32][9];
    ele[15][9] != ele[33][9];
    ele[15][9] != ele[34][9];
    ele[15][9] != ele[35][9];
    ele[16][0] != ele[16][1];
    ele[16][0] != ele[16][10];
    ele[16][0] != ele[16][11];
    ele[16][0] != ele[16][12];
    ele[16][0] != ele[16][13];
    ele[16][0] != ele[16][14];
    ele[16][0] != ele[16][15];
    ele[16][0] != ele[16][16];
    ele[16][0] != ele[16][17];
    ele[16][0] != ele[16][18];
    ele[16][0] != ele[16][19];
    ele[16][0] != ele[16][2];
    ele[16][0] != ele[16][20];
    ele[16][0] != ele[16][21];
    ele[16][0] != ele[16][22];
    ele[16][0] != ele[16][23];
    ele[16][0] != ele[16][24];
    ele[16][0] != ele[16][25];
    ele[16][0] != ele[16][26];
    ele[16][0] != ele[16][27];
    ele[16][0] != ele[16][28];
    ele[16][0] != ele[16][29];
    ele[16][0] != ele[16][3];
    ele[16][0] != ele[16][30];
    ele[16][0] != ele[16][31];
    ele[16][0] != ele[16][32];
    ele[16][0] != ele[16][33];
    ele[16][0] != ele[16][34];
    ele[16][0] != ele[16][35];
    ele[16][0] != ele[16][4];
    ele[16][0] != ele[16][5];
    ele[16][0] != ele[16][6];
    ele[16][0] != ele[16][7];
    ele[16][0] != ele[16][8];
    ele[16][0] != ele[16][9];
    ele[16][0] != ele[17][0];
    ele[16][0] != ele[17][1];
    ele[16][0] != ele[17][2];
    ele[16][0] != ele[17][3];
    ele[16][0] != ele[17][4];
    ele[16][0] != ele[17][5];
    ele[16][0] != ele[18][0];
    ele[16][0] != ele[19][0];
    ele[16][0] != ele[20][0];
    ele[16][0] != ele[21][0];
    ele[16][0] != ele[22][0];
    ele[16][0] != ele[23][0];
    ele[16][0] != ele[24][0];
    ele[16][0] != ele[25][0];
    ele[16][0] != ele[26][0];
    ele[16][0] != ele[27][0];
    ele[16][0] != ele[28][0];
    ele[16][0] != ele[29][0];
    ele[16][0] != ele[30][0];
    ele[16][0] != ele[31][0];
    ele[16][0] != ele[32][0];
    ele[16][0] != ele[33][0];
    ele[16][0] != ele[34][0];
    ele[16][0] != ele[35][0];
    ele[16][1] != ele[16][10];
    ele[16][1] != ele[16][11];
    ele[16][1] != ele[16][12];
    ele[16][1] != ele[16][13];
    ele[16][1] != ele[16][14];
    ele[16][1] != ele[16][15];
    ele[16][1] != ele[16][16];
    ele[16][1] != ele[16][17];
    ele[16][1] != ele[16][18];
    ele[16][1] != ele[16][19];
    ele[16][1] != ele[16][2];
    ele[16][1] != ele[16][20];
    ele[16][1] != ele[16][21];
    ele[16][1] != ele[16][22];
    ele[16][1] != ele[16][23];
    ele[16][1] != ele[16][24];
    ele[16][1] != ele[16][25];
    ele[16][1] != ele[16][26];
    ele[16][1] != ele[16][27];
    ele[16][1] != ele[16][28];
    ele[16][1] != ele[16][29];
    ele[16][1] != ele[16][3];
    ele[16][1] != ele[16][30];
    ele[16][1] != ele[16][31];
    ele[16][1] != ele[16][32];
    ele[16][1] != ele[16][33];
    ele[16][1] != ele[16][34];
    ele[16][1] != ele[16][35];
    ele[16][1] != ele[16][4];
    ele[16][1] != ele[16][5];
    ele[16][1] != ele[16][6];
    ele[16][1] != ele[16][7];
    ele[16][1] != ele[16][8];
    ele[16][1] != ele[16][9];
    ele[16][1] != ele[17][0];
    ele[16][1] != ele[17][1];
    ele[16][1] != ele[17][2];
    ele[16][1] != ele[17][3];
    ele[16][1] != ele[17][4];
    ele[16][1] != ele[17][5];
    ele[16][1] != ele[18][1];
    ele[16][1] != ele[19][1];
    ele[16][1] != ele[20][1];
    ele[16][1] != ele[21][1];
    ele[16][1] != ele[22][1];
    ele[16][1] != ele[23][1];
    ele[16][1] != ele[24][1];
    ele[16][1] != ele[25][1];
    ele[16][1] != ele[26][1];
    ele[16][1] != ele[27][1];
    ele[16][1] != ele[28][1];
    ele[16][1] != ele[29][1];
    ele[16][1] != ele[30][1];
    ele[16][1] != ele[31][1];
    ele[16][1] != ele[32][1];
    ele[16][1] != ele[33][1];
    ele[16][1] != ele[34][1];
    ele[16][1] != ele[35][1];
    ele[16][10] != ele[16][11];
    ele[16][10] != ele[16][12];
    ele[16][10] != ele[16][13];
    ele[16][10] != ele[16][14];
    ele[16][10] != ele[16][15];
    ele[16][10] != ele[16][16];
    ele[16][10] != ele[16][17];
    ele[16][10] != ele[16][18];
    ele[16][10] != ele[16][19];
    ele[16][10] != ele[16][20];
    ele[16][10] != ele[16][21];
    ele[16][10] != ele[16][22];
    ele[16][10] != ele[16][23];
    ele[16][10] != ele[16][24];
    ele[16][10] != ele[16][25];
    ele[16][10] != ele[16][26];
    ele[16][10] != ele[16][27];
    ele[16][10] != ele[16][28];
    ele[16][10] != ele[16][29];
    ele[16][10] != ele[16][30];
    ele[16][10] != ele[16][31];
    ele[16][10] != ele[16][32];
    ele[16][10] != ele[16][33];
    ele[16][10] != ele[16][34];
    ele[16][10] != ele[16][35];
    ele[16][10] != ele[17][10];
    ele[16][10] != ele[17][11];
    ele[16][10] != ele[17][6];
    ele[16][10] != ele[17][7];
    ele[16][10] != ele[17][8];
    ele[16][10] != ele[17][9];
    ele[16][10] != ele[18][10];
    ele[16][10] != ele[19][10];
    ele[16][10] != ele[20][10];
    ele[16][10] != ele[21][10];
    ele[16][10] != ele[22][10];
    ele[16][10] != ele[23][10];
    ele[16][10] != ele[24][10];
    ele[16][10] != ele[25][10];
    ele[16][10] != ele[26][10];
    ele[16][10] != ele[27][10];
    ele[16][10] != ele[28][10];
    ele[16][10] != ele[29][10];
    ele[16][10] != ele[30][10];
    ele[16][10] != ele[31][10];
    ele[16][10] != ele[32][10];
    ele[16][10] != ele[33][10];
    ele[16][10] != ele[34][10];
    ele[16][10] != ele[35][10];
    ele[16][11] != ele[16][12];
    ele[16][11] != ele[16][13];
    ele[16][11] != ele[16][14];
    ele[16][11] != ele[16][15];
    ele[16][11] != ele[16][16];
    ele[16][11] != ele[16][17];
    ele[16][11] != ele[16][18];
    ele[16][11] != ele[16][19];
    ele[16][11] != ele[16][20];
    ele[16][11] != ele[16][21];
    ele[16][11] != ele[16][22];
    ele[16][11] != ele[16][23];
    ele[16][11] != ele[16][24];
    ele[16][11] != ele[16][25];
    ele[16][11] != ele[16][26];
    ele[16][11] != ele[16][27];
    ele[16][11] != ele[16][28];
    ele[16][11] != ele[16][29];
    ele[16][11] != ele[16][30];
    ele[16][11] != ele[16][31];
    ele[16][11] != ele[16][32];
    ele[16][11] != ele[16][33];
    ele[16][11] != ele[16][34];
    ele[16][11] != ele[16][35];
    ele[16][11] != ele[17][10];
    ele[16][11] != ele[17][11];
    ele[16][11] != ele[17][6];
    ele[16][11] != ele[17][7];
    ele[16][11] != ele[17][8];
    ele[16][11] != ele[17][9];
    ele[16][11] != ele[18][11];
    ele[16][11] != ele[19][11];
    ele[16][11] != ele[20][11];
    ele[16][11] != ele[21][11];
    ele[16][11] != ele[22][11];
    ele[16][11] != ele[23][11];
    ele[16][11] != ele[24][11];
    ele[16][11] != ele[25][11];
    ele[16][11] != ele[26][11];
    ele[16][11] != ele[27][11];
    ele[16][11] != ele[28][11];
    ele[16][11] != ele[29][11];
    ele[16][11] != ele[30][11];
    ele[16][11] != ele[31][11];
    ele[16][11] != ele[32][11];
    ele[16][11] != ele[33][11];
    ele[16][11] != ele[34][11];
    ele[16][11] != ele[35][11];
    ele[16][12] != ele[16][13];
    ele[16][12] != ele[16][14];
    ele[16][12] != ele[16][15];
    ele[16][12] != ele[16][16];
    ele[16][12] != ele[16][17];
    ele[16][12] != ele[16][18];
    ele[16][12] != ele[16][19];
    ele[16][12] != ele[16][20];
    ele[16][12] != ele[16][21];
    ele[16][12] != ele[16][22];
    ele[16][12] != ele[16][23];
    ele[16][12] != ele[16][24];
    ele[16][12] != ele[16][25];
    ele[16][12] != ele[16][26];
    ele[16][12] != ele[16][27];
    ele[16][12] != ele[16][28];
    ele[16][12] != ele[16][29];
    ele[16][12] != ele[16][30];
    ele[16][12] != ele[16][31];
    ele[16][12] != ele[16][32];
    ele[16][12] != ele[16][33];
    ele[16][12] != ele[16][34];
    ele[16][12] != ele[16][35];
    ele[16][12] != ele[17][12];
    ele[16][12] != ele[17][13];
    ele[16][12] != ele[17][14];
    ele[16][12] != ele[17][15];
    ele[16][12] != ele[17][16];
    ele[16][12] != ele[17][17];
    ele[16][12] != ele[18][12];
    ele[16][12] != ele[19][12];
    ele[16][12] != ele[20][12];
    ele[16][12] != ele[21][12];
    ele[16][12] != ele[22][12];
    ele[16][12] != ele[23][12];
    ele[16][12] != ele[24][12];
    ele[16][12] != ele[25][12];
    ele[16][12] != ele[26][12];
    ele[16][12] != ele[27][12];
    ele[16][12] != ele[28][12];
    ele[16][12] != ele[29][12];
    ele[16][12] != ele[30][12];
    ele[16][12] != ele[31][12];
    ele[16][12] != ele[32][12];
    ele[16][12] != ele[33][12];
    ele[16][12] != ele[34][12];
    ele[16][12] != ele[35][12];
    ele[16][13] != ele[16][14];
    ele[16][13] != ele[16][15];
    ele[16][13] != ele[16][16];
    ele[16][13] != ele[16][17];
    ele[16][13] != ele[16][18];
    ele[16][13] != ele[16][19];
    ele[16][13] != ele[16][20];
    ele[16][13] != ele[16][21];
    ele[16][13] != ele[16][22];
    ele[16][13] != ele[16][23];
    ele[16][13] != ele[16][24];
    ele[16][13] != ele[16][25];
    ele[16][13] != ele[16][26];
    ele[16][13] != ele[16][27];
    ele[16][13] != ele[16][28];
    ele[16][13] != ele[16][29];
    ele[16][13] != ele[16][30];
    ele[16][13] != ele[16][31];
    ele[16][13] != ele[16][32];
    ele[16][13] != ele[16][33];
    ele[16][13] != ele[16][34];
    ele[16][13] != ele[16][35];
    ele[16][13] != ele[17][12];
    ele[16][13] != ele[17][13];
    ele[16][13] != ele[17][14];
    ele[16][13] != ele[17][15];
    ele[16][13] != ele[17][16];
    ele[16][13] != ele[17][17];
    ele[16][13] != ele[18][13];
    ele[16][13] != ele[19][13];
    ele[16][13] != ele[20][13];
    ele[16][13] != ele[21][13];
    ele[16][13] != ele[22][13];
    ele[16][13] != ele[23][13];
    ele[16][13] != ele[24][13];
    ele[16][13] != ele[25][13];
    ele[16][13] != ele[26][13];
    ele[16][13] != ele[27][13];
    ele[16][13] != ele[28][13];
    ele[16][13] != ele[29][13];
    ele[16][13] != ele[30][13];
    ele[16][13] != ele[31][13];
    ele[16][13] != ele[32][13];
    ele[16][13] != ele[33][13];
    ele[16][13] != ele[34][13];
    ele[16][13] != ele[35][13];
    ele[16][14] != ele[16][15];
    ele[16][14] != ele[16][16];
    ele[16][14] != ele[16][17];
    ele[16][14] != ele[16][18];
    ele[16][14] != ele[16][19];
    ele[16][14] != ele[16][20];
    ele[16][14] != ele[16][21];
    ele[16][14] != ele[16][22];
    ele[16][14] != ele[16][23];
    ele[16][14] != ele[16][24];
    ele[16][14] != ele[16][25];
    ele[16][14] != ele[16][26];
    ele[16][14] != ele[16][27];
    ele[16][14] != ele[16][28];
    ele[16][14] != ele[16][29];
    ele[16][14] != ele[16][30];
    ele[16][14] != ele[16][31];
    ele[16][14] != ele[16][32];
    ele[16][14] != ele[16][33];
    ele[16][14] != ele[16][34];
    ele[16][14] != ele[16][35];
    ele[16][14] != ele[17][12];
    ele[16][14] != ele[17][13];
    ele[16][14] != ele[17][14];
    ele[16][14] != ele[17][15];
    ele[16][14] != ele[17][16];
    ele[16][14] != ele[17][17];
    ele[16][14] != ele[18][14];
    ele[16][14] != ele[19][14];
    ele[16][14] != ele[20][14];
    ele[16][14] != ele[21][14];
    ele[16][14] != ele[22][14];
    ele[16][14] != ele[23][14];
    ele[16][14] != ele[24][14];
    ele[16][14] != ele[25][14];
    ele[16][14] != ele[26][14];
    ele[16][14] != ele[27][14];
    ele[16][14] != ele[28][14];
    ele[16][14] != ele[29][14];
    ele[16][14] != ele[30][14];
    ele[16][14] != ele[31][14];
    ele[16][14] != ele[32][14];
    ele[16][14] != ele[33][14];
    ele[16][14] != ele[34][14];
    ele[16][14] != ele[35][14];
    ele[16][15] != ele[16][16];
    ele[16][15] != ele[16][17];
    ele[16][15] != ele[16][18];
    ele[16][15] != ele[16][19];
    ele[16][15] != ele[16][20];
    ele[16][15] != ele[16][21];
    ele[16][15] != ele[16][22];
    ele[16][15] != ele[16][23];
    ele[16][15] != ele[16][24];
    ele[16][15] != ele[16][25];
    ele[16][15] != ele[16][26];
    ele[16][15] != ele[16][27];
    ele[16][15] != ele[16][28];
    ele[16][15] != ele[16][29];
    ele[16][15] != ele[16][30];
    ele[16][15] != ele[16][31];
    ele[16][15] != ele[16][32];
    ele[16][15] != ele[16][33];
    ele[16][15] != ele[16][34];
    ele[16][15] != ele[16][35];
    ele[16][15] != ele[17][12];
    ele[16][15] != ele[17][13];
    ele[16][15] != ele[17][14];
    ele[16][15] != ele[17][15];
    ele[16][15] != ele[17][16];
    ele[16][15] != ele[17][17];
    ele[16][15] != ele[18][15];
    ele[16][15] != ele[19][15];
    ele[16][15] != ele[20][15];
    ele[16][15] != ele[21][15];
    ele[16][15] != ele[22][15];
    ele[16][15] != ele[23][15];
    ele[16][15] != ele[24][15];
    ele[16][15] != ele[25][15];
    ele[16][15] != ele[26][15];
    ele[16][15] != ele[27][15];
    ele[16][15] != ele[28][15];
    ele[16][15] != ele[29][15];
    ele[16][15] != ele[30][15];
    ele[16][15] != ele[31][15];
    ele[16][15] != ele[32][15];
    ele[16][15] != ele[33][15];
    ele[16][15] != ele[34][15];
    ele[16][15] != ele[35][15];
    ele[16][16] != ele[16][17];
    ele[16][16] != ele[16][18];
    ele[16][16] != ele[16][19];
    ele[16][16] != ele[16][20];
    ele[16][16] != ele[16][21];
    ele[16][16] != ele[16][22];
    ele[16][16] != ele[16][23];
    ele[16][16] != ele[16][24];
    ele[16][16] != ele[16][25];
    ele[16][16] != ele[16][26];
    ele[16][16] != ele[16][27];
    ele[16][16] != ele[16][28];
    ele[16][16] != ele[16][29];
    ele[16][16] != ele[16][30];
    ele[16][16] != ele[16][31];
    ele[16][16] != ele[16][32];
    ele[16][16] != ele[16][33];
    ele[16][16] != ele[16][34];
    ele[16][16] != ele[16][35];
    ele[16][16] != ele[17][12];
    ele[16][16] != ele[17][13];
    ele[16][16] != ele[17][14];
    ele[16][16] != ele[17][15];
    ele[16][16] != ele[17][16];
    ele[16][16] != ele[17][17];
    ele[16][16] != ele[18][16];
    ele[16][16] != ele[19][16];
    ele[16][16] != ele[20][16];
    ele[16][16] != ele[21][16];
    ele[16][16] != ele[22][16];
    ele[16][16] != ele[23][16];
    ele[16][16] != ele[24][16];
    ele[16][16] != ele[25][16];
    ele[16][16] != ele[26][16];
    ele[16][16] != ele[27][16];
    ele[16][16] != ele[28][16];
    ele[16][16] != ele[29][16];
    ele[16][16] != ele[30][16];
    ele[16][16] != ele[31][16];
    ele[16][16] != ele[32][16];
    ele[16][16] != ele[33][16];
    ele[16][16] != ele[34][16];
    ele[16][16] != ele[35][16];
    ele[16][17] != ele[16][18];
    ele[16][17] != ele[16][19];
    ele[16][17] != ele[16][20];
    ele[16][17] != ele[16][21];
    ele[16][17] != ele[16][22];
    ele[16][17] != ele[16][23];
    ele[16][17] != ele[16][24];
    ele[16][17] != ele[16][25];
    ele[16][17] != ele[16][26];
    ele[16][17] != ele[16][27];
    ele[16][17] != ele[16][28];
    ele[16][17] != ele[16][29];
    ele[16][17] != ele[16][30];
    ele[16][17] != ele[16][31];
    ele[16][17] != ele[16][32];
    ele[16][17] != ele[16][33];
    ele[16][17] != ele[16][34];
    ele[16][17] != ele[16][35];
    ele[16][17] != ele[17][12];
    ele[16][17] != ele[17][13];
    ele[16][17] != ele[17][14];
    ele[16][17] != ele[17][15];
    ele[16][17] != ele[17][16];
    ele[16][17] != ele[17][17];
    ele[16][17] != ele[18][17];
    ele[16][17] != ele[19][17];
    ele[16][17] != ele[20][17];
    ele[16][17] != ele[21][17];
    ele[16][17] != ele[22][17];
    ele[16][17] != ele[23][17];
    ele[16][17] != ele[24][17];
    ele[16][17] != ele[25][17];
    ele[16][17] != ele[26][17];
    ele[16][17] != ele[27][17];
    ele[16][17] != ele[28][17];
    ele[16][17] != ele[29][17];
    ele[16][17] != ele[30][17];
    ele[16][17] != ele[31][17];
    ele[16][17] != ele[32][17];
    ele[16][17] != ele[33][17];
    ele[16][17] != ele[34][17];
    ele[16][17] != ele[35][17];
    ele[16][18] != ele[16][19];
    ele[16][18] != ele[16][20];
    ele[16][18] != ele[16][21];
    ele[16][18] != ele[16][22];
    ele[16][18] != ele[16][23];
    ele[16][18] != ele[16][24];
    ele[16][18] != ele[16][25];
    ele[16][18] != ele[16][26];
    ele[16][18] != ele[16][27];
    ele[16][18] != ele[16][28];
    ele[16][18] != ele[16][29];
    ele[16][18] != ele[16][30];
    ele[16][18] != ele[16][31];
    ele[16][18] != ele[16][32];
    ele[16][18] != ele[16][33];
    ele[16][18] != ele[16][34];
    ele[16][18] != ele[16][35];
    ele[16][18] != ele[17][18];
    ele[16][18] != ele[17][19];
    ele[16][18] != ele[17][20];
    ele[16][18] != ele[17][21];
    ele[16][18] != ele[17][22];
    ele[16][18] != ele[17][23];
    ele[16][18] != ele[18][18];
    ele[16][18] != ele[19][18];
    ele[16][18] != ele[20][18];
    ele[16][18] != ele[21][18];
    ele[16][18] != ele[22][18];
    ele[16][18] != ele[23][18];
    ele[16][18] != ele[24][18];
    ele[16][18] != ele[25][18];
    ele[16][18] != ele[26][18];
    ele[16][18] != ele[27][18];
    ele[16][18] != ele[28][18];
    ele[16][18] != ele[29][18];
    ele[16][18] != ele[30][18];
    ele[16][18] != ele[31][18];
    ele[16][18] != ele[32][18];
    ele[16][18] != ele[33][18];
    ele[16][18] != ele[34][18];
    ele[16][18] != ele[35][18];
    ele[16][19] != ele[16][20];
    ele[16][19] != ele[16][21];
    ele[16][19] != ele[16][22];
    ele[16][19] != ele[16][23];
    ele[16][19] != ele[16][24];
    ele[16][19] != ele[16][25];
    ele[16][19] != ele[16][26];
    ele[16][19] != ele[16][27];
    ele[16][19] != ele[16][28];
    ele[16][19] != ele[16][29];
    ele[16][19] != ele[16][30];
    ele[16][19] != ele[16][31];
    ele[16][19] != ele[16][32];
    ele[16][19] != ele[16][33];
    ele[16][19] != ele[16][34];
    ele[16][19] != ele[16][35];
    ele[16][19] != ele[17][18];
    ele[16][19] != ele[17][19];
    ele[16][19] != ele[17][20];
    ele[16][19] != ele[17][21];
    ele[16][19] != ele[17][22];
    ele[16][19] != ele[17][23];
    ele[16][19] != ele[18][19];
    ele[16][19] != ele[19][19];
    ele[16][19] != ele[20][19];
    ele[16][19] != ele[21][19];
    ele[16][19] != ele[22][19];
    ele[16][19] != ele[23][19];
    ele[16][19] != ele[24][19];
    ele[16][19] != ele[25][19];
    ele[16][19] != ele[26][19];
    ele[16][19] != ele[27][19];
    ele[16][19] != ele[28][19];
    ele[16][19] != ele[29][19];
    ele[16][19] != ele[30][19];
    ele[16][19] != ele[31][19];
    ele[16][19] != ele[32][19];
    ele[16][19] != ele[33][19];
    ele[16][19] != ele[34][19];
    ele[16][19] != ele[35][19];
    ele[16][2] != ele[16][10];
    ele[16][2] != ele[16][11];
    ele[16][2] != ele[16][12];
    ele[16][2] != ele[16][13];
    ele[16][2] != ele[16][14];
    ele[16][2] != ele[16][15];
    ele[16][2] != ele[16][16];
    ele[16][2] != ele[16][17];
    ele[16][2] != ele[16][18];
    ele[16][2] != ele[16][19];
    ele[16][2] != ele[16][20];
    ele[16][2] != ele[16][21];
    ele[16][2] != ele[16][22];
    ele[16][2] != ele[16][23];
    ele[16][2] != ele[16][24];
    ele[16][2] != ele[16][25];
    ele[16][2] != ele[16][26];
    ele[16][2] != ele[16][27];
    ele[16][2] != ele[16][28];
    ele[16][2] != ele[16][29];
    ele[16][2] != ele[16][3];
    ele[16][2] != ele[16][30];
    ele[16][2] != ele[16][31];
    ele[16][2] != ele[16][32];
    ele[16][2] != ele[16][33];
    ele[16][2] != ele[16][34];
    ele[16][2] != ele[16][35];
    ele[16][2] != ele[16][4];
    ele[16][2] != ele[16][5];
    ele[16][2] != ele[16][6];
    ele[16][2] != ele[16][7];
    ele[16][2] != ele[16][8];
    ele[16][2] != ele[16][9];
    ele[16][2] != ele[17][0];
    ele[16][2] != ele[17][1];
    ele[16][2] != ele[17][2];
    ele[16][2] != ele[17][3];
    ele[16][2] != ele[17][4];
    ele[16][2] != ele[17][5];
    ele[16][2] != ele[18][2];
    ele[16][2] != ele[19][2];
    ele[16][2] != ele[20][2];
    ele[16][2] != ele[21][2];
    ele[16][2] != ele[22][2];
    ele[16][2] != ele[23][2];
    ele[16][2] != ele[24][2];
    ele[16][2] != ele[25][2];
    ele[16][2] != ele[26][2];
    ele[16][2] != ele[27][2];
    ele[16][2] != ele[28][2];
    ele[16][2] != ele[29][2];
    ele[16][2] != ele[30][2];
    ele[16][2] != ele[31][2];
    ele[16][2] != ele[32][2];
    ele[16][2] != ele[33][2];
    ele[16][2] != ele[34][2];
    ele[16][2] != ele[35][2];
    ele[16][20] != ele[16][21];
    ele[16][20] != ele[16][22];
    ele[16][20] != ele[16][23];
    ele[16][20] != ele[16][24];
    ele[16][20] != ele[16][25];
    ele[16][20] != ele[16][26];
    ele[16][20] != ele[16][27];
    ele[16][20] != ele[16][28];
    ele[16][20] != ele[16][29];
    ele[16][20] != ele[16][30];
    ele[16][20] != ele[16][31];
    ele[16][20] != ele[16][32];
    ele[16][20] != ele[16][33];
    ele[16][20] != ele[16][34];
    ele[16][20] != ele[16][35];
    ele[16][20] != ele[17][18];
    ele[16][20] != ele[17][19];
    ele[16][20] != ele[17][20];
    ele[16][20] != ele[17][21];
    ele[16][20] != ele[17][22];
    ele[16][20] != ele[17][23];
    ele[16][20] != ele[18][20];
    ele[16][20] != ele[19][20];
    ele[16][20] != ele[20][20];
    ele[16][20] != ele[21][20];
    ele[16][20] != ele[22][20];
    ele[16][20] != ele[23][20];
    ele[16][20] != ele[24][20];
    ele[16][20] != ele[25][20];
    ele[16][20] != ele[26][20];
    ele[16][20] != ele[27][20];
    ele[16][20] != ele[28][20];
    ele[16][20] != ele[29][20];
    ele[16][20] != ele[30][20];
    ele[16][20] != ele[31][20];
    ele[16][20] != ele[32][20];
    ele[16][20] != ele[33][20];
    ele[16][20] != ele[34][20];
    ele[16][20] != ele[35][20];
    ele[16][21] != ele[16][22];
    ele[16][21] != ele[16][23];
    ele[16][21] != ele[16][24];
    ele[16][21] != ele[16][25];
    ele[16][21] != ele[16][26];
    ele[16][21] != ele[16][27];
    ele[16][21] != ele[16][28];
    ele[16][21] != ele[16][29];
    ele[16][21] != ele[16][30];
    ele[16][21] != ele[16][31];
    ele[16][21] != ele[16][32];
    ele[16][21] != ele[16][33];
    ele[16][21] != ele[16][34];
    ele[16][21] != ele[16][35];
    ele[16][21] != ele[17][18];
    ele[16][21] != ele[17][19];
    ele[16][21] != ele[17][20];
    ele[16][21] != ele[17][21];
    ele[16][21] != ele[17][22];
    ele[16][21] != ele[17][23];
    ele[16][21] != ele[18][21];
    ele[16][21] != ele[19][21];
    ele[16][21] != ele[20][21];
    ele[16][21] != ele[21][21];
    ele[16][21] != ele[22][21];
    ele[16][21] != ele[23][21];
    ele[16][21] != ele[24][21];
    ele[16][21] != ele[25][21];
    ele[16][21] != ele[26][21];
    ele[16][21] != ele[27][21];
    ele[16][21] != ele[28][21];
    ele[16][21] != ele[29][21];
    ele[16][21] != ele[30][21];
    ele[16][21] != ele[31][21];
    ele[16][21] != ele[32][21];
    ele[16][21] != ele[33][21];
    ele[16][21] != ele[34][21];
    ele[16][21] != ele[35][21];
    ele[16][22] != ele[16][23];
    ele[16][22] != ele[16][24];
    ele[16][22] != ele[16][25];
    ele[16][22] != ele[16][26];
    ele[16][22] != ele[16][27];
    ele[16][22] != ele[16][28];
    ele[16][22] != ele[16][29];
    ele[16][22] != ele[16][30];
    ele[16][22] != ele[16][31];
    ele[16][22] != ele[16][32];
    ele[16][22] != ele[16][33];
    ele[16][22] != ele[16][34];
    ele[16][22] != ele[16][35];
    ele[16][22] != ele[17][18];
    ele[16][22] != ele[17][19];
    ele[16][22] != ele[17][20];
    ele[16][22] != ele[17][21];
    ele[16][22] != ele[17][22];
    ele[16][22] != ele[17][23];
    ele[16][22] != ele[18][22];
    ele[16][22] != ele[19][22];
    ele[16][22] != ele[20][22];
    ele[16][22] != ele[21][22];
    ele[16][22] != ele[22][22];
    ele[16][22] != ele[23][22];
    ele[16][22] != ele[24][22];
    ele[16][22] != ele[25][22];
    ele[16][22] != ele[26][22];
    ele[16][22] != ele[27][22];
    ele[16][22] != ele[28][22];
    ele[16][22] != ele[29][22];
    ele[16][22] != ele[30][22];
    ele[16][22] != ele[31][22];
    ele[16][22] != ele[32][22];
    ele[16][22] != ele[33][22];
    ele[16][22] != ele[34][22];
    ele[16][22] != ele[35][22];
    ele[16][23] != ele[16][24];
    ele[16][23] != ele[16][25];
    ele[16][23] != ele[16][26];
    ele[16][23] != ele[16][27];
    ele[16][23] != ele[16][28];
    ele[16][23] != ele[16][29];
    ele[16][23] != ele[16][30];
    ele[16][23] != ele[16][31];
    ele[16][23] != ele[16][32];
    ele[16][23] != ele[16][33];
    ele[16][23] != ele[16][34];
    ele[16][23] != ele[16][35];
    ele[16][23] != ele[17][18];
    ele[16][23] != ele[17][19];
    ele[16][23] != ele[17][20];
    ele[16][23] != ele[17][21];
    ele[16][23] != ele[17][22];
    ele[16][23] != ele[17][23];
    ele[16][23] != ele[18][23];
    ele[16][23] != ele[19][23];
    ele[16][23] != ele[20][23];
    ele[16][23] != ele[21][23];
    ele[16][23] != ele[22][23];
    ele[16][23] != ele[23][23];
    ele[16][23] != ele[24][23];
    ele[16][23] != ele[25][23];
    ele[16][23] != ele[26][23];
    ele[16][23] != ele[27][23];
    ele[16][23] != ele[28][23];
    ele[16][23] != ele[29][23];
    ele[16][23] != ele[30][23];
    ele[16][23] != ele[31][23];
    ele[16][23] != ele[32][23];
    ele[16][23] != ele[33][23];
    ele[16][23] != ele[34][23];
    ele[16][23] != ele[35][23];
    ele[16][24] != ele[16][25];
    ele[16][24] != ele[16][26];
    ele[16][24] != ele[16][27];
    ele[16][24] != ele[16][28];
    ele[16][24] != ele[16][29];
    ele[16][24] != ele[16][30];
    ele[16][24] != ele[16][31];
    ele[16][24] != ele[16][32];
    ele[16][24] != ele[16][33];
    ele[16][24] != ele[16][34];
    ele[16][24] != ele[16][35];
    ele[16][24] != ele[17][24];
    ele[16][24] != ele[17][25];
    ele[16][24] != ele[17][26];
    ele[16][24] != ele[17][27];
    ele[16][24] != ele[17][28];
    ele[16][24] != ele[17][29];
    ele[16][24] != ele[18][24];
    ele[16][24] != ele[19][24];
    ele[16][24] != ele[20][24];
    ele[16][24] != ele[21][24];
    ele[16][24] != ele[22][24];
    ele[16][24] != ele[23][24];
    ele[16][24] != ele[24][24];
    ele[16][24] != ele[25][24];
    ele[16][24] != ele[26][24];
    ele[16][24] != ele[27][24];
    ele[16][24] != ele[28][24];
    ele[16][24] != ele[29][24];
    ele[16][24] != ele[30][24];
    ele[16][24] != ele[31][24];
    ele[16][24] != ele[32][24];
    ele[16][24] != ele[33][24];
    ele[16][24] != ele[34][24];
    ele[16][24] != ele[35][24];
    ele[16][25] != ele[16][26];
    ele[16][25] != ele[16][27];
    ele[16][25] != ele[16][28];
    ele[16][25] != ele[16][29];
    ele[16][25] != ele[16][30];
    ele[16][25] != ele[16][31];
    ele[16][25] != ele[16][32];
    ele[16][25] != ele[16][33];
    ele[16][25] != ele[16][34];
    ele[16][25] != ele[16][35];
    ele[16][25] != ele[17][24];
    ele[16][25] != ele[17][25];
    ele[16][25] != ele[17][26];
    ele[16][25] != ele[17][27];
    ele[16][25] != ele[17][28];
    ele[16][25] != ele[17][29];
    ele[16][25] != ele[18][25];
    ele[16][25] != ele[19][25];
    ele[16][25] != ele[20][25];
    ele[16][25] != ele[21][25];
    ele[16][25] != ele[22][25];
    ele[16][25] != ele[23][25];
    ele[16][25] != ele[24][25];
    ele[16][25] != ele[25][25];
    ele[16][25] != ele[26][25];
    ele[16][25] != ele[27][25];
    ele[16][25] != ele[28][25];
    ele[16][25] != ele[29][25];
    ele[16][25] != ele[30][25];
    ele[16][25] != ele[31][25];
    ele[16][25] != ele[32][25];
    ele[16][25] != ele[33][25];
    ele[16][25] != ele[34][25];
    ele[16][25] != ele[35][25];
    ele[16][26] != ele[16][27];
    ele[16][26] != ele[16][28];
    ele[16][26] != ele[16][29];
    ele[16][26] != ele[16][30];
    ele[16][26] != ele[16][31];
    ele[16][26] != ele[16][32];
    ele[16][26] != ele[16][33];
    ele[16][26] != ele[16][34];
    ele[16][26] != ele[16][35];
    ele[16][26] != ele[17][24];
    ele[16][26] != ele[17][25];
    ele[16][26] != ele[17][26];
    ele[16][26] != ele[17][27];
    ele[16][26] != ele[17][28];
    ele[16][26] != ele[17][29];
    ele[16][26] != ele[18][26];
    ele[16][26] != ele[19][26];
    ele[16][26] != ele[20][26];
    ele[16][26] != ele[21][26];
    ele[16][26] != ele[22][26];
    ele[16][26] != ele[23][26];
    ele[16][26] != ele[24][26];
    ele[16][26] != ele[25][26];
    ele[16][26] != ele[26][26];
    ele[16][26] != ele[27][26];
    ele[16][26] != ele[28][26];
    ele[16][26] != ele[29][26];
    ele[16][26] != ele[30][26];
    ele[16][26] != ele[31][26];
    ele[16][26] != ele[32][26];
    ele[16][26] != ele[33][26];
    ele[16][26] != ele[34][26];
    ele[16][26] != ele[35][26];
    ele[16][27] != ele[16][28];
    ele[16][27] != ele[16][29];
    ele[16][27] != ele[16][30];
    ele[16][27] != ele[16][31];
    ele[16][27] != ele[16][32];
    ele[16][27] != ele[16][33];
    ele[16][27] != ele[16][34];
    ele[16][27] != ele[16][35];
    ele[16][27] != ele[17][24];
    ele[16][27] != ele[17][25];
    ele[16][27] != ele[17][26];
    ele[16][27] != ele[17][27];
    ele[16][27] != ele[17][28];
    ele[16][27] != ele[17][29];
    ele[16][27] != ele[18][27];
    ele[16][27] != ele[19][27];
    ele[16][27] != ele[20][27];
    ele[16][27] != ele[21][27];
    ele[16][27] != ele[22][27];
    ele[16][27] != ele[23][27];
    ele[16][27] != ele[24][27];
    ele[16][27] != ele[25][27];
    ele[16][27] != ele[26][27];
    ele[16][27] != ele[27][27];
    ele[16][27] != ele[28][27];
    ele[16][27] != ele[29][27];
    ele[16][27] != ele[30][27];
    ele[16][27] != ele[31][27];
    ele[16][27] != ele[32][27];
    ele[16][27] != ele[33][27];
    ele[16][27] != ele[34][27];
    ele[16][27] != ele[35][27];
    ele[16][28] != ele[16][29];
    ele[16][28] != ele[16][30];
    ele[16][28] != ele[16][31];
    ele[16][28] != ele[16][32];
    ele[16][28] != ele[16][33];
    ele[16][28] != ele[16][34];
    ele[16][28] != ele[16][35];
    ele[16][28] != ele[17][24];
    ele[16][28] != ele[17][25];
    ele[16][28] != ele[17][26];
    ele[16][28] != ele[17][27];
    ele[16][28] != ele[17][28];
    ele[16][28] != ele[17][29];
    ele[16][28] != ele[18][28];
    ele[16][28] != ele[19][28];
    ele[16][28] != ele[20][28];
    ele[16][28] != ele[21][28];
    ele[16][28] != ele[22][28];
    ele[16][28] != ele[23][28];
    ele[16][28] != ele[24][28];
    ele[16][28] != ele[25][28];
    ele[16][28] != ele[26][28];
    ele[16][28] != ele[27][28];
    ele[16][28] != ele[28][28];
    ele[16][28] != ele[29][28];
    ele[16][28] != ele[30][28];
    ele[16][28] != ele[31][28];
    ele[16][28] != ele[32][28];
    ele[16][28] != ele[33][28];
    ele[16][28] != ele[34][28];
    ele[16][28] != ele[35][28];
    ele[16][29] != ele[16][30];
    ele[16][29] != ele[16][31];
    ele[16][29] != ele[16][32];
    ele[16][29] != ele[16][33];
    ele[16][29] != ele[16][34];
    ele[16][29] != ele[16][35];
    ele[16][29] != ele[17][24];
    ele[16][29] != ele[17][25];
    ele[16][29] != ele[17][26];
    ele[16][29] != ele[17][27];
    ele[16][29] != ele[17][28];
    ele[16][29] != ele[17][29];
    ele[16][29] != ele[18][29];
    ele[16][29] != ele[19][29];
    ele[16][29] != ele[20][29];
    ele[16][29] != ele[21][29];
    ele[16][29] != ele[22][29];
    ele[16][29] != ele[23][29];
    ele[16][29] != ele[24][29];
    ele[16][29] != ele[25][29];
    ele[16][29] != ele[26][29];
    ele[16][29] != ele[27][29];
    ele[16][29] != ele[28][29];
    ele[16][29] != ele[29][29];
    ele[16][29] != ele[30][29];
    ele[16][29] != ele[31][29];
    ele[16][29] != ele[32][29];
    ele[16][29] != ele[33][29];
    ele[16][29] != ele[34][29];
    ele[16][29] != ele[35][29];
    ele[16][3] != ele[16][10];
    ele[16][3] != ele[16][11];
    ele[16][3] != ele[16][12];
    ele[16][3] != ele[16][13];
    ele[16][3] != ele[16][14];
    ele[16][3] != ele[16][15];
    ele[16][3] != ele[16][16];
    ele[16][3] != ele[16][17];
    ele[16][3] != ele[16][18];
    ele[16][3] != ele[16][19];
    ele[16][3] != ele[16][20];
    ele[16][3] != ele[16][21];
    ele[16][3] != ele[16][22];
    ele[16][3] != ele[16][23];
    ele[16][3] != ele[16][24];
    ele[16][3] != ele[16][25];
    ele[16][3] != ele[16][26];
    ele[16][3] != ele[16][27];
    ele[16][3] != ele[16][28];
    ele[16][3] != ele[16][29];
    ele[16][3] != ele[16][30];
    ele[16][3] != ele[16][31];
    ele[16][3] != ele[16][32];
    ele[16][3] != ele[16][33];
    ele[16][3] != ele[16][34];
    ele[16][3] != ele[16][35];
    ele[16][3] != ele[16][4];
    ele[16][3] != ele[16][5];
    ele[16][3] != ele[16][6];
    ele[16][3] != ele[16][7];
    ele[16][3] != ele[16][8];
    ele[16][3] != ele[16][9];
    ele[16][3] != ele[17][0];
    ele[16][3] != ele[17][1];
    ele[16][3] != ele[17][2];
    ele[16][3] != ele[17][3];
    ele[16][3] != ele[17][4];
    ele[16][3] != ele[17][5];
    ele[16][3] != ele[18][3];
    ele[16][3] != ele[19][3];
    ele[16][3] != ele[20][3];
    ele[16][3] != ele[21][3];
    ele[16][3] != ele[22][3];
    ele[16][3] != ele[23][3];
    ele[16][3] != ele[24][3];
    ele[16][3] != ele[25][3];
    ele[16][3] != ele[26][3];
    ele[16][3] != ele[27][3];
    ele[16][3] != ele[28][3];
    ele[16][3] != ele[29][3];
    ele[16][3] != ele[30][3];
    ele[16][3] != ele[31][3];
    ele[16][3] != ele[32][3];
    ele[16][3] != ele[33][3];
    ele[16][3] != ele[34][3];
    ele[16][3] != ele[35][3];
    ele[16][30] != ele[16][31];
    ele[16][30] != ele[16][32];
    ele[16][30] != ele[16][33];
    ele[16][30] != ele[16][34];
    ele[16][30] != ele[16][35];
    ele[16][30] != ele[17][30];
    ele[16][30] != ele[17][31];
    ele[16][30] != ele[17][32];
    ele[16][30] != ele[17][33];
    ele[16][30] != ele[17][34];
    ele[16][30] != ele[17][35];
    ele[16][30] != ele[18][30];
    ele[16][30] != ele[19][30];
    ele[16][30] != ele[20][30];
    ele[16][30] != ele[21][30];
    ele[16][30] != ele[22][30];
    ele[16][30] != ele[23][30];
    ele[16][30] != ele[24][30];
    ele[16][30] != ele[25][30];
    ele[16][30] != ele[26][30];
    ele[16][30] != ele[27][30];
    ele[16][30] != ele[28][30];
    ele[16][30] != ele[29][30];
    ele[16][30] != ele[30][30];
    ele[16][30] != ele[31][30];
    ele[16][30] != ele[32][30];
    ele[16][30] != ele[33][30];
    ele[16][30] != ele[34][30];
    ele[16][30] != ele[35][30];
    ele[16][31] != ele[16][32];
    ele[16][31] != ele[16][33];
    ele[16][31] != ele[16][34];
    ele[16][31] != ele[16][35];
    ele[16][31] != ele[17][30];
    ele[16][31] != ele[17][31];
    ele[16][31] != ele[17][32];
    ele[16][31] != ele[17][33];
    ele[16][31] != ele[17][34];
    ele[16][31] != ele[17][35];
    ele[16][31] != ele[18][31];
    ele[16][31] != ele[19][31];
    ele[16][31] != ele[20][31];
    ele[16][31] != ele[21][31];
    ele[16][31] != ele[22][31];
    ele[16][31] != ele[23][31];
    ele[16][31] != ele[24][31];
    ele[16][31] != ele[25][31];
    ele[16][31] != ele[26][31];
    ele[16][31] != ele[27][31];
    ele[16][31] != ele[28][31];
    ele[16][31] != ele[29][31];
    ele[16][31] != ele[30][31];
    ele[16][31] != ele[31][31];
    ele[16][31] != ele[32][31];
    ele[16][31] != ele[33][31];
    ele[16][31] != ele[34][31];
    ele[16][31] != ele[35][31];
    ele[16][32] != ele[16][33];
    ele[16][32] != ele[16][34];
    ele[16][32] != ele[16][35];
    ele[16][32] != ele[17][30];
    ele[16][32] != ele[17][31];
    ele[16][32] != ele[17][32];
    ele[16][32] != ele[17][33];
    ele[16][32] != ele[17][34];
    ele[16][32] != ele[17][35];
    ele[16][32] != ele[18][32];
    ele[16][32] != ele[19][32];
    ele[16][32] != ele[20][32];
    ele[16][32] != ele[21][32];
    ele[16][32] != ele[22][32];
    ele[16][32] != ele[23][32];
    ele[16][32] != ele[24][32];
    ele[16][32] != ele[25][32];
    ele[16][32] != ele[26][32];
    ele[16][32] != ele[27][32];
    ele[16][32] != ele[28][32];
    ele[16][32] != ele[29][32];
    ele[16][32] != ele[30][32];
    ele[16][32] != ele[31][32];
    ele[16][32] != ele[32][32];
    ele[16][32] != ele[33][32];
    ele[16][32] != ele[34][32];
    ele[16][32] != ele[35][32];
    ele[16][33] != ele[16][34];
    ele[16][33] != ele[16][35];
    ele[16][33] != ele[17][30];
    ele[16][33] != ele[17][31];
    ele[16][33] != ele[17][32];
    ele[16][33] != ele[17][33];
    ele[16][33] != ele[17][34];
    ele[16][33] != ele[17][35];
    ele[16][33] != ele[18][33];
    ele[16][33] != ele[19][33];
    ele[16][33] != ele[20][33];
    ele[16][33] != ele[21][33];
    ele[16][33] != ele[22][33];
    ele[16][33] != ele[23][33];
    ele[16][33] != ele[24][33];
    ele[16][33] != ele[25][33];
    ele[16][33] != ele[26][33];
    ele[16][33] != ele[27][33];
    ele[16][33] != ele[28][33];
    ele[16][33] != ele[29][33];
    ele[16][33] != ele[30][33];
    ele[16][33] != ele[31][33];
    ele[16][33] != ele[32][33];
    ele[16][33] != ele[33][33];
    ele[16][33] != ele[34][33];
    ele[16][33] != ele[35][33];
    ele[16][34] != ele[16][35];
    ele[16][34] != ele[17][30];
    ele[16][34] != ele[17][31];
    ele[16][34] != ele[17][32];
    ele[16][34] != ele[17][33];
    ele[16][34] != ele[17][34];
    ele[16][34] != ele[17][35];
    ele[16][34] != ele[18][34];
    ele[16][34] != ele[19][34];
    ele[16][34] != ele[20][34];
    ele[16][34] != ele[21][34];
    ele[16][34] != ele[22][34];
    ele[16][34] != ele[23][34];
    ele[16][34] != ele[24][34];
    ele[16][34] != ele[25][34];
    ele[16][34] != ele[26][34];
    ele[16][34] != ele[27][34];
    ele[16][34] != ele[28][34];
    ele[16][34] != ele[29][34];
    ele[16][34] != ele[30][34];
    ele[16][34] != ele[31][34];
    ele[16][34] != ele[32][34];
    ele[16][34] != ele[33][34];
    ele[16][34] != ele[34][34];
    ele[16][34] != ele[35][34];
    ele[16][35] != ele[17][30];
    ele[16][35] != ele[17][31];
    ele[16][35] != ele[17][32];
    ele[16][35] != ele[17][33];
    ele[16][35] != ele[17][34];
    ele[16][35] != ele[17][35];
    ele[16][35] != ele[18][35];
    ele[16][35] != ele[19][35];
    ele[16][35] != ele[20][35];
    ele[16][35] != ele[21][35];
    ele[16][35] != ele[22][35];
    ele[16][35] != ele[23][35];
    ele[16][35] != ele[24][35];
    ele[16][35] != ele[25][35];
    ele[16][35] != ele[26][35];
    ele[16][35] != ele[27][35];
    ele[16][35] != ele[28][35];
    ele[16][35] != ele[29][35];
    ele[16][35] != ele[30][35];
    ele[16][35] != ele[31][35];
    ele[16][35] != ele[32][35];
    ele[16][35] != ele[33][35];
    ele[16][35] != ele[34][35];
    ele[16][35] != ele[35][35];
    ele[16][4] != ele[16][10];
    ele[16][4] != ele[16][11];
    ele[16][4] != ele[16][12];
    ele[16][4] != ele[16][13];
    ele[16][4] != ele[16][14];
    ele[16][4] != ele[16][15];
    ele[16][4] != ele[16][16];
    ele[16][4] != ele[16][17];
    ele[16][4] != ele[16][18];
    ele[16][4] != ele[16][19];
    ele[16][4] != ele[16][20];
    ele[16][4] != ele[16][21];
    ele[16][4] != ele[16][22];
    ele[16][4] != ele[16][23];
    ele[16][4] != ele[16][24];
    ele[16][4] != ele[16][25];
    ele[16][4] != ele[16][26];
    ele[16][4] != ele[16][27];
    ele[16][4] != ele[16][28];
    ele[16][4] != ele[16][29];
    ele[16][4] != ele[16][30];
    ele[16][4] != ele[16][31];
    ele[16][4] != ele[16][32];
    ele[16][4] != ele[16][33];
    ele[16][4] != ele[16][34];
    ele[16][4] != ele[16][35];
    ele[16][4] != ele[16][5];
    ele[16][4] != ele[16][6];
    ele[16][4] != ele[16][7];
    ele[16][4] != ele[16][8];
    ele[16][4] != ele[16][9];
    ele[16][4] != ele[17][0];
    ele[16][4] != ele[17][1];
    ele[16][4] != ele[17][2];
    ele[16][4] != ele[17][3];
    ele[16][4] != ele[17][4];
    ele[16][4] != ele[17][5];
    ele[16][4] != ele[18][4];
    ele[16][4] != ele[19][4];
    ele[16][4] != ele[20][4];
    ele[16][4] != ele[21][4];
    ele[16][4] != ele[22][4];
    ele[16][4] != ele[23][4];
    ele[16][4] != ele[24][4];
    ele[16][4] != ele[25][4];
    ele[16][4] != ele[26][4];
    ele[16][4] != ele[27][4];
    ele[16][4] != ele[28][4];
    ele[16][4] != ele[29][4];
    ele[16][4] != ele[30][4];
    ele[16][4] != ele[31][4];
    ele[16][4] != ele[32][4];
    ele[16][4] != ele[33][4];
    ele[16][4] != ele[34][4];
    ele[16][4] != ele[35][4];
    ele[16][5] != ele[16][10];
    ele[16][5] != ele[16][11];
    ele[16][5] != ele[16][12];
    ele[16][5] != ele[16][13];
    ele[16][5] != ele[16][14];
    ele[16][5] != ele[16][15];
    ele[16][5] != ele[16][16];
    ele[16][5] != ele[16][17];
    ele[16][5] != ele[16][18];
    ele[16][5] != ele[16][19];
    ele[16][5] != ele[16][20];
    ele[16][5] != ele[16][21];
    ele[16][5] != ele[16][22];
    ele[16][5] != ele[16][23];
    ele[16][5] != ele[16][24];
    ele[16][5] != ele[16][25];
    ele[16][5] != ele[16][26];
    ele[16][5] != ele[16][27];
    ele[16][5] != ele[16][28];
    ele[16][5] != ele[16][29];
    ele[16][5] != ele[16][30];
    ele[16][5] != ele[16][31];
    ele[16][5] != ele[16][32];
    ele[16][5] != ele[16][33];
    ele[16][5] != ele[16][34];
    ele[16][5] != ele[16][35];
    ele[16][5] != ele[16][6];
    ele[16][5] != ele[16][7];
    ele[16][5] != ele[16][8];
    ele[16][5] != ele[16][9];
    ele[16][5] != ele[17][0];
    ele[16][5] != ele[17][1];
    ele[16][5] != ele[17][2];
    ele[16][5] != ele[17][3];
    ele[16][5] != ele[17][4];
    ele[16][5] != ele[17][5];
    ele[16][5] != ele[18][5];
    ele[16][5] != ele[19][5];
    ele[16][5] != ele[20][5];
    ele[16][5] != ele[21][5];
    ele[16][5] != ele[22][5];
    ele[16][5] != ele[23][5];
    ele[16][5] != ele[24][5];
    ele[16][5] != ele[25][5];
    ele[16][5] != ele[26][5];
    ele[16][5] != ele[27][5];
    ele[16][5] != ele[28][5];
    ele[16][5] != ele[29][5];
    ele[16][5] != ele[30][5];
    ele[16][5] != ele[31][5];
    ele[16][5] != ele[32][5];
    ele[16][5] != ele[33][5];
    ele[16][5] != ele[34][5];
    ele[16][5] != ele[35][5];
    ele[16][6] != ele[16][10];
    ele[16][6] != ele[16][11];
    ele[16][6] != ele[16][12];
    ele[16][6] != ele[16][13];
    ele[16][6] != ele[16][14];
    ele[16][6] != ele[16][15];
    ele[16][6] != ele[16][16];
    ele[16][6] != ele[16][17];
    ele[16][6] != ele[16][18];
    ele[16][6] != ele[16][19];
    ele[16][6] != ele[16][20];
    ele[16][6] != ele[16][21];
    ele[16][6] != ele[16][22];
    ele[16][6] != ele[16][23];
    ele[16][6] != ele[16][24];
    ele[16][6] != ele[16][25];
    ele[16][6] != ele[16][26];
    ele[16][6] != ele[16][27];
    ele[16][6] != ele[16][28];
    ele[16][6] != ele[16][29];
    ele[16][6] != ele[16][30];
    ele[16][6] != ele[16][31];
    ele[16][6] != ele[16][32];
    ele[16][6] != ele[16][33];
    ele[16][6] != ele[16][34];
    ele[16][6] != ele[16][35];
    ele[16][6] != ele[16][7];
    ele[16][6] != ele[16][8];
    ele[16][6] != ele[16][9];
    ele[16][6] != ele[17][10];
    ele[16][6] != ele[17][11];
    ele[16][6] != ele[17][6];
    ele[16][6] != ele[17][7];
    ele[16][6] != ele[17][8];
    ele[16][6] != ele[17][9];
    ele[16][6] != ele[18][6];
    ele[16][6] != ele[19][6];
    ele[16][6] != ele[20][6];
    ele[16][6] != ele[21][6];
    ele[16][6] != ele[22][6];
    ele[16][6] != ele[23][6];
    ele[16][6] != ele[24][6];
    ele[16][6] != ele[25][6];
    ele[16][6] != ele[26][6];
    ele[16][6] != ele[27][6];
    ele[16][6] != ele[28][6];
    ele[16][6] != ele[29][6];
    ele[16][6] != ele[30][6];
    ele[16][6] != ele[31][6];
    ele[16][6] != ele[32][6];
    ele[16][6] != ele[33][6];
    ele[16][6] != ele[34][6];
    ele[16][6] != ele[35][6];
    ele[16][7] != ele[16][10];
    ele[16][7] != ele[16][11];
    ele[16][7] != ele[16][12];
    ele[16][7] != ele[16][13];
    ele[16][7] != ele[16][14];
    ele[16][7] != ele[16][15];
    ele[16][7] != ele[16][16];
    ele[16][7] != ele[16][17];
    ele[16][7] != ele[16][18];
    ele[16][7] != ele[16][19];
    ele[16][7] != ele[16][20];
    ele[16][7] != ele[16][21];
    ele[16][7] != ele[16][22];
    ele[16][7] != ele[16][23];
    ele[16][7] != ele[16][24];
    ele[16][7] != ele[16][25];
    ele[16][7] != ele[16][26];
    ele[16][7] != ele[16][27];
    ele[16][7] != ele[16][28];
    ele[16][7] != ele[16][29];
    ele[16][7] != ele[16][30];
    ele[16][7] != ele[16][31];
    ele[16][7] != ele[16][32];
    ele[16][7] != ele[16][33];
    ele[16][7] != ele[16][34];
    ele[16][7] != ele[16][35];
    ele[16][7] != ele[16][8];
    ele[16][7] != ele[16][9];
    ele[16][7] != ele[17][10];
    ele[16][7] != ele[17][11];
    ele[16][7] != ele[17][6];
    ele[16][7] != ele[17][7];
    ele[16][7] != ele[17][8];
    ele[16][7] != ele[17][9];
    ele[16][7] != ele[18][7];
    ele[16][7] != ele[19][7];
    ele[16][7] != ele[20][7];
    ele[16][7] != ele[21][7];
    ele[16][7] != ele[22][7];
    ele[16][7] != ele[23][7];
    ele[16][7] != ele[24][7];
    ele[16][7] != ele[25][7];
    ele[16][7] != ele[26][7];
    ele[16][7] != ele[27][7];
    ele[16][7] != ele[28][7];
    ele[16][7] != ele[29][7];
    ele[16][7] != ele[30][7];
    ele[16][7] != ele[31][7];
    ele[16][7] != ele[32][7];
    ele[16][7] != ele[33][7];
    ele[16][7] != ele[34][7];
    ele[16][7] != ele[35][7];
    ele[16][8] != ele[16][10];
    ele[16][8] != ele[16][11];
    ele[16][8] != ele[16][12];
    ele[16][8] != ele[16][13];
    ele[16][8] != ele[16][14];
    ele[16][8] != ele[16][15];
    ele[16][8] != ele[16][16];
    ele[16][8] != ele[16][17];
    ele[16][8] != ele[16][18];
    ele[16][8] != ele[16][19];
    ele[16][8] != ele[16][20];
    ele[16][8] != ele[16][21];
    ele[16][8] != ele[16][22];
    ele[16][8] != ele[16][23];
    ele[16][8] != ele[16][24];
    ele[16][8] != ele[16][25];
    ele[16][8] != ele[16][26];
    ele[16][8] != ele[16][27];
    ele[16][8] != ele[16][28];
    ele[16][8] != ele[16][29];
    ele[16][8] != ele[16][30];
    ele[16][8] != ele[16][31];
    ele[16][8] != ele[16][32];
    ele[16][8] != ele[16][33];
    ele[16][8] != ele[16][34];
    ele[16][8] != ele[16][35];
    ele[16][8] != ele[16][9];
    ele[16][8] != ele[17][10];
    ele[16][8] != ele[17][11];
    ele[16][8] != ele[17][6];
    ele[16][8] != ele[17][7];
    ele[16][8] != ele[17][8];
    ele[16][8] != ele[17][9];
    ele[16][8] != ele[18][8];
    ele[16][8] != ele[19][8];
    ele[16][8] != ele[20][8];
    ele[16][8] != ele[21][8];
    ele[16][8] != ele[22][8];
    ele[16][8] != ele[23][8];
    ele[16][8] != ele[24][8];
    ele[16][8] != ele[25][8];
    ele[16][8] != ele[26][8];
    ele[16][8] != ele[27][8];
    ele[16][8] != ele[28][8];
    ele[16][8] != ele[29][8];
    ele[16][8] != ele[30][8];
    ele[16][8] != ele[31][8];
    ele[16][8] != ele[32][8];
    ele[16][8] != ele[33][8];
    ele[16][8] != ele[34][8];
    ele[16][8] != ele[35][8];
    ele[16][9] != ele[16][10];
    ele[16][9] != ele[16][11];
    ele[16][9] != ele[16][12];
    ele[16][9] != ele[16][13];
    ele[16][9] != ele[16][14];
    ele[16][9] != ele[16][15];
    ele[16][9] != ele[16][16];
    ele[16][9] != ele[16][17];
    ele[16][9] != ele[16][18];
    ele[16][9] != ele[16][19];
    ele[16][9] != ele[16][20];
    ele[16][9] != ele[16][21];
    ele[16][9] != ele[16][22];
    ele[16][9] != ele[16][23];
    ele[16][9] != ele[16][24];
    ele[16][9] != ele[16][25];
    ele[16][9] != ele[16][26];
    ele[16][9] != ele[16][27];
    ele[16][9] != ele[16][28];
    ele[16][9] != ele[16][29];
    ele[16][9] != ele[16][30];
    ele[16][9] != ele[16][31];
    ele[16][9] != ele[16][32];
    ele[16][9] != ele[16][33];
    ele[16][9] != ele[16][34];
    ele[16][9] != ele[16][35];
    ele[16][9] != ele[17][10];
    ele[16][9] != ele[17][11];
    ele[16][9] != ele[17][6];
    ele[16][9] != ele[17][7];
    ele[16][9] != ele[17][8];
    ele[16][9] != ele[17][9];
    ele[16][9] != ele[18][9];
    ele[16][9] != ele[19][9];
    ele[16][9] != ele[20][9];
    ele[16][9] != ele[21][9];
    ele[16][9] != ele[22][9];
    ele[16][9] != ele[23][9];
    ele[16][9] != ele[24][9];
    ele[16][9] != ele[25][9];
    ele[16][9] != ele[26][9];
    ele[16][9] != ele[27][9];
    ele[16][9] != ele[28][9];
    ele[16][9] != ele[29][9];
    ele[16][9] != ele[30][9];
    ele[16][9] != ele[31][9];
    ele[16][9] != ele[32][9];
    ele[16][9] != ele[33][9];
    ele[16][9] != ele[34][9];
    ele[16][9] != ele[35][9];
    ele[17][0] != ele[17][1];
    ele[17][0] != ele[17][10];
    ele[17][0] != ele[17][11];
    ele[17][0] != ele[17][12];
    ele[17][0] != ele[17][13];
    ele[17][0] != ele[17][14];
    ele[17][0] != ele[17][15];
    ele[17][0] != ele[17][16];
    ele[17][0] != ele[17][17];
    ele[17][0] != ele[17][18];
    ele[17][0] != ele[17][19];
    ele[17][0] != ele[17][2];
    ele[17][0] != ele[17][20];
    ele[17][0] != ele[17][21];
    ele[17][0] != ele[17][22];
    ele[17][0] != ele[17][23];
    ele[17][0] != ele[17][24];
    ele[17][0] != ele[17][25];
    ele[17][0] != ele[17][26];
    ele[17][0] != ele[17][27];
    ele[17][0] != ele[17][28];
    ele[17][0] != ele[17][29];
    ele[17][0] != ele[17][3];
    ele[17][0] != ele[17][30];
    ele[17][0] != ele[17][31];
    ele[17][0] != ele[17][32];
    ele[17][0] != ele[17][33];
    ele[17][0] != ele[17][34];
    ele[17][0] != ele[17][35];
    ele[17][0] != ele[17][4];
    ele[17][0] != ele[17][5];
    ele[17][0] != ele[17][6];
    ele[17][0] != ele[17][7];
    ele[17][0] != ele[17][8];
    ele[17][0] != ele[17][9];
    ele[17][0] != ele[18][0];
    ele[17][0] != ele[19][0];
    ele[17][0] != ele[20][0];
    ele[17][0] != ele[21][0];
    ele[17][0] != ele[22][0];
    ele[17][0] != ele[23][0];
    ele[17][0] != ele[24][0];
    ele[17][0] != ele[25][0];
    ele[17][0] != ele[26][0];
    ele[17][0] != ele[27][0];
    ele[17][0] != ele[28][0];
    ele[17][0] != ele[29][0];
    ele[17][0] != ele[30][0];
    ele[17][0] != ele[31][0];
    ele[17][0] != ele[32][0];
    ele[17][0] != ele[33][0];
    ele[17][0] != ele[34][0];
    ele[17][0] != ele[35][0];
    ele[17][1] != ele[17][10];
    ele[17][1] != ele[17][11];
    ele[17][1] != ele[17][12];
    ele[17][1] != ele[17][13];
    ele[17][1] != ele[17][14];
    ele[17][1] != ele[17][15];
    ele[17][1] != ele[17][16];
    ele[17][1] != ele[17][17];
    ele[17][1] != ele[17][18];
    ele[17][1] != ele[17][19];
    ele[17][1] != ele[17][2];
    ele[17][1] != ele[17][20];
    ele[17][1] != ele[17][21];
    ele[17][1] != ele[17][22];
    ele[17][1] != ele[17][23];
    ele[17][1] != ele[17][24];
    ele[17][1] != ele[17][25];
    ele[17][1] != ele[17][26];
    ele[17][1] != ele[17][27];
    ele[17][1] != ele[17][28];
    ele[17][1] != ele[17][29];
    ele[17][1] != ele[17][3];
    ele[17][1] != ele[17][30];
    ele[17][1] != ele[17][31];
    ele[17][1] != ele[17][32];
    ele[17][1] != ele[17][33];
    ele[17][1] != ele[17][34];
    ele[17][1] != ele[17][35];
    ele[17][1] != ele[17][4];
    ele[17][1] != ele[17][5];
    ele[17][1] != ele[17][6];
    ele[17][1] != ele[17][7];
    ele[17][1] != ele[17][8];
    ele[17][1] != ele[17][9];
    ele[17][1] != ele[18][1];
    ele[17][1] != ele[19][1];
    ele[17][1] != ele[20][1];
    ele[17][1] != ele[21][1];
    ele[17][1] != ele[22][1];
    ele[17][1] != ele[23][1];
    ele[17][1] != ele[24][1];
    ele[17][1] != ele[25][1];
    ele[17][1] != ele[26][1];
    ele[17][1] != ele[27][1];
    ele[17][1] != ele[28][1];
    ele[17][1] != ele[29][1];
    ele[17][1] != ele[30][1];
    ele[17][1] != ele[31][1];
    ele[17][1] != ele[32][1];
    ele[17][1] != ele[33][1];
    ele[17][1] != ele[34][1];
    ele[17][1] != ele[35][1];
    ele[17][10] != ele[17][11];
    ele[17][10] != ele[17][12];
    ele[17][10] != ele[17][13];
    ele[17][10] != ele[17][14];
    ele[17][10] != ele[17][15];
    ele[17][10] != ele[17][16];
    ele[17][10] != ele[17][17];
    ele[17][10] != ele[17][18];
    ele[17][10] != ele[17][19];
    ele[17][10] != ele[17][20];
    ele[17][10] != ele[17][21];
    ele[17][10] != ele[17][22];
    ele[17][10] != ele[17][23];
    ele[17][10] != ele[17][24];
    ele[17][10] != ele[17][25];
    ele[17][10] != ele[17][26];
    ele[17][10] != ele[17][27];
    ele[17][10] != ele[17][28];
    ele[17][10] != ele[17][29];
    ele[17][10] != ele[17][30];
    ele[17][10] != ele[17][31];
    ele[17][10] != ele[17][32];
    ele[17][10] != ele[17][33];
    ele[17][10] != ele[17][34];
    ele[17][10] != ele[17][35];
    ele[17][10] != ele[18][10];
    ele[17][10] != ele[19][10];
    ele[17][10] != ele[20][10];
    ele[17][10] != ele[21][10];
    ele[17][10] != ele[22][10];
    ele[17][10] != ele[23][10];
    ele[17][10] != ele[24][10];
    ele[17][10] != ele[25][10];
    ele[17][10] != ele[26][10];
    ele[17][10] != ele[27][10];
    ele[17][10] != ele[28][10];
    ele[17][10] != ele[29][10];
    ele[17][10] != ele[30][10];
    ele[17][10] != ele[31][10];
    ele[17][10] != ele[32][10];
    ele[17][10] != ele[33][10];
    ele[17][10] != ele[34][10];
    ele[17][10] != ele[35][10];
    ele[17][11] != ele[17][12];
    ele[17][11] != ele[17][13];
    ele[17][11] != ele[17][14];
    ele[17][11] != ele[17][15];
    ele[17][11] != ele[17][16];
    ele[17][11] != ele[17][17];
    ele[17][11] != ele[17][18];
    ele[17][11] != ele[17][19];
    ele[17][11] != ele[17][20];
    ele[17][11] != ele[17][21];
    ele[17][11] != ele[17][22];
    ele[17][11] != ele[17][23];
    ele[17][11] != ele[17][24];
    ele[17][11] != ele[17][25];
    ele[17][11] != ele[17][26];
    ele[17][11] != ele[17][27];
    ele[17][11] != ele[17][28];
    ele[17][11] != ele[17][29];
    ele[17][11] != ele[17][30];
    ele[17][11] != ele[17][31];
    ele[17][11] != ele[17][32];
    ele[17][11] != ele[17][33];
    ele[17][11] != ele[17][34];
    ele[17][11] != ele[17][35];
    ele[17][11] != ele[18][11];
    ele[17][11] != ele[19][11];
    ele[17][11] != ele[20][11];
    ele[17][11] != ele[21][11];
    ele[17][11] != ele[22][11];
    ele[17][11] != ele[23][11];
    ele[17][11] != ele[24][11];
    ele[17][11] != ele[25][11];
    ele[17][11] != ele[26][11];
    ele[17][11] != ele[27][11];
    ele[17][11] != ele[28][11];
    ele[17][11] != ele[29][11];
    ele[17][11] != ele[30][11];
    ele[17][11] != ele[31][11];
    ele[17][11] != ele[32][11];
    ele[17][11] != ele[33][11];
    ele[17][11] != ele[34][11];
    ele[17][11] != ele[35][11];
    ele[17][12] != ele[17][13];
    ele[17][12] != ele[17][14];
    ele[17][12] != ele[17][15];
    ele[17][12] != ele[17][16];
    ele[17][12] != ele[17][17];
    ele[17][12] != ele[17][18];
    ele[17][12] != ele[17][19];
    ele[17][12] != ele[17][20];
    ele[17][12] != ele[17][21];
    ele[17][12] != ele[17][22];
    ele[17][12] != ele[17][23];
    ele[17][12] != ele[17][24];
    ele[17][12] != ele[17][25];
    ele[17][12] != ele[17][26];
    ele[17][12] != ele[17][27];
    ele[17][12] != ele[17][28];
    ele[17][12] != ele[17][29];
    ele[17][12] != ele[17][30];
    ele[17][12] != ele[17][31];
    ele[17][12] != ele[17][32];
    ele[17][12] != ele[17][33];
    ele[17][12] != ele[17][34];
    ele[17][12] != ele[17][35];
    ele[17][12] != ele[18][12];
    ele[17][12] != ele[19][12];
    ele[17][12] != ele[20][12];
    ele[17][12] != ele[21][12];
    ele[17][12] != ele[22][12];
    ele[17][12] != ele[23][12];
    ele[17][12] != ele[24][12];
    ele[17][12] != ele[25][12];
    ele[17][12] != ele[26][12];
    ele[17][12] != ele[27][12];
    ele[17][12] != ele[28][12];
    ele[17][12] != ele[29][12];
    ele[17][12] != ele[30][12];
    ele[17][12] != ele[31][12];
    ele[17][12] != ele[32][12];
    ele[17][12] != ele[33][12];
    ele[17][12] != ele[34][12];
    ele[17][12] != ele[35][12];
    ele[17][13] != ele[17][14];
    ele[17][13] != ele[17][15];
    ele[17][13] != ele[17][16];
    ele[17][13] != ele[17][17];
    ele[17][13] != ele[17][18];
    ele[17][13] != ele[17][19];
    ele[17][13] != ele[17][20];
    ele[17][13] != ele[17][21];
    ele[17][13] != ele[17][22];
    ele[17][13] != ele[17][23];
    ele[17][13] != ele[17][24];
    ele[17][13] != ele[17][25];
    ele[17][13] != ele[17][26];
    ele[17][13] != ele[17][27];
    ele[17][13] != ele[17][28];
    ele[17][13] != ele[17][29];
    ele[17][13] != ele[17][30];
    ele[17][13] != ele[17][31];
    ele[17][13] != ele[17][32];
    ele[17][13] != ele[17][33];
    ele[17][13] != ele[17][34];
    ele[17][13] != ele[17][35];
    ele[17][13] != ele[18][13];
    ele[17][13] != ele[19][13];
    ele[17][13] != ele[20][13];
    ele[17][13] != ele[21][13];
    ele[17][13] != ele[22][13];
    ele[17][13] != ele[23][13];
    ele[17][13] != ele[24][13];
    ele[17][13] != ele[25][13];
    ele[17][13] != ele[26][13];
    ele[17][13] != ele[27][13];
    ele[17][13] != ele[28][13];
    ele[17][13] != ele[29][13];
    ele[17][13] != ele[30][13];
    ele[17][13] != ele[31][13];
    ele[17][13] != ele[32][13];
    ele[17][13] != ele[33][13];
    ele[17][13] != ele[34][13];
    ele[17][13] != ele[35][13];
    ele[17][14] != ele[17][15];
    ele[17][14] != ele[17][16];
    ele[17][14] != ele[17][17];
    ele[17][14] != ele[17][18];
    ele[17][14] != ele[17][19];
    ele[17][14] != ele[17][20];
    ele[17][14] != ele[17][21];
    ele[17][14] != ele[17][22];
    ele[17][14] != ele[17][23];
    ele[17][14] != ele[17][24];
    ele[17][14] != ele[17][25];
    ele[17][14] != ele[17][26];
    ele[17][14] != ele[17][27];
    ele[17][14] != ele[17][28];
    ele[17][14] != ele[17][29];
    ele[17][14] != ele[17][30];
    ele[17][14] != ele[17][31];
    ele[17][14] != ele[17][32];
    ele[17][14] != ele[17][33];
    ele[17][14] != ele[17][34];
    ele[17][14] != ele[17][35];
    ele[17][14] != ele[18][14];
    ele[17][14] != ele[19][14];
    ele[17][14] != ele[20][14];
    ele[17][14] != ele[21][14];
    ele[17][14] != ele[22][14];
    ele[17][14] != ele[23][14];
    ele[17][14] != ele[24][14];
    ele[17][14] != ele[25][14];
    ele[17][14] != ele[26][14];
    ele[17][14] != ele[27][14];
    ele[17][14] != ele[28][14];
    ele[17][14] != ele[29][14];
    ele[17][14] != ele[30][14];
    ele[17][14] != ele[31][14];
    ele[17][14] != ele[32][14];
    ele[17][14] != ele[33][14];
    ele[17][14] != ele[34][14];
    ele[17][14] != ele[35][14];
    ele[17][15] != ele[17][16];
    ele[17][15] != ele[17][17];
    ele[17][15] != ele[17][18];
    ele[17][15] != ele[17][19];
    ele[17][15] != ele[17][20];
    ele[17][15] != ele[17][21];
    ele[17][15] != ele[17][22];
    ele[17][15] != ele[17][23];
    ele[17][15] != ele[17][24];
    ele[17][15] != ele[17][25];
    ele[17][15] != ele[17][26];
    ele[17][15] != ele[17][27];
    ele[17][15] != ele[17][28];
    ele[17][15] != ele[17][29];
    ele[17][15] != ele[17][30];
    ele[17][15] != ele[17][31];
    ele[17][15] != ele[17][32];
    ele[17][15] != ele[17][33];
    ele[17][15] != ele[17][34];
    ele[17][15] != ele[17][35];
    ele[17][15] != ele[18][15];
    ele[17][15] != ele[19][15];
    ele[17][15] != ele[20][15];
    ele[17][15] != ele[21][15];
    ele[17][15] != ele[22][15];
    ele[17][15] != ele[23][15];
    ele[17][15] != ele[24][15];
    ele[17][15] != ele[25][15];
    ele[17][15] != ele[26][15];
    ele[17][15] != ele[27][15];
    ele[17][15] != ele[28][15];
    ele[17][15] != ele[29][15];
    ele[17][15] != ele[30][15];
    ele[17][15] != ele[31][15];
    ele[17][15] != ele[32][15];
    ele[17][15] != ele[33][15];
    ele[17][15] != ele[34][15];
    ele[17][15] != ele[35][15];
    ele[17][16] != ele[17][17];
    ele[17][16] != ele[17][18];
    ele[17][16] != ele[17][19];
    ele[17][16] != ele[17][20];
    ele[17][16] != ele[17][21];
    ele[17][16] != ele[17][22];
    ele[17][16] != ele[17][23];
    ele[17][16] != ele[17][24];
    ele[17][16] != ele[17][25];
    ele[17][16] != ele[17][26];
    ele[17][16] != ele[17][27];
    ele[17][16] != ele[17][28];
    ele[17][16] != ele[17][29];
    ele[17][16] != ele[17][30];
    ele[17][16] != ele[17][31];
    ele[17][16] != ele[17][32];
    ele[17][16] != ele[17][33];
    ele[17][16] != ele[17][34];
    ele[17][16] != ele[17][35];
    ele[17][16] != ele[18][16];
    ele[17][16] != ele[19][16];
    ele[17][16] != ele[20][16];
    ele[17][16] != ele[21][16];
    ele[17][16] != ele[22][16];
    ele[17][16] != ele[23][16];
    ele[17][16] != ele[24][16];
    ele[17][16] != ele[25][16];
    ele[17][16] != ele[26][16];
    ele[17][16] != ele[27][16];
    ele[17][16] != ele[28][16];
    ele[17][16] != ele[29][16];
    ele[17][16] != ele[30][16];
    ele[17][16] != ele[31][16];
    ele[17][16] != ele[32][16];
    ele[17][16] != ele[33][16];
    ele[17][16] != ele[34][16];
    ele[17][16] != ele[35][16];
    ele[17][17] != ele[17][18];
    ele[17][17] != ele[17][19];
    ele[17][17] != ele[17][20];
    ele[17][17] != ele[17][21];
    ele[17][17] != ele[17][22];
    ele[17][17] != ele[17][23];
    ele[17][17] != ele[17][24];
    ele[17][17] != ele[17][25];
    ele[17][17] != ele[17][26];
    ele[17][17] != ele[17][27];
    ele[17][17] != ele[17][28];
    ele[17][17] != ele[17][29];
    ele[17][17] != ele[17][30];
    ele[17][17] != ele[17][31];
    ele[17][17] != ele[17][32];
    ele[17][17] != ele[17][33];
    ele[17][17] != ele[17][34];
    ele[17][17] != ele[17][35];
    ele[17][17] != ele[18][17];
    ele[17][17] != ele[19][17];
    ele[17][17] != ele[20][17];
    ele[17][17] != ele[21][17];
    ele[17][17] != ele[22][17];
    ele[17][17] != ele[23][17];
    ele[17][17] != ele[24][17];
    ele[17][17] != ele[25][17];
    ele[17][17] != ele[26][17];
    ele[17][17] != ele[27][17];
    ele[17][17] != ele[28][17];
    ele[17][17] != ele[29][17];
    ele[17][17] != ele[30][17];
    ele[17][17] != ele[31][17];
    ele[17][17] != ele[32][17];
    ele[17][17] != ele[33][17];
    ele[17][17] != ele[34][17];
    ele[17][17] != ele[35][17];
    ele[17][18] != ele[17][19];
    ele[17][18] != ele[17][20];
    ele[17][18] != ele[17][21];
    ele[17][18] != ele[17][22];
    ele[17][18] != ele[17][23];
    ele[17][18] != ele[17][24];
    ele[17][18] != ele[17][25];
    ele[17][18] != ele[17][26];
    ele[17][18] != ele[17][27];
    ele[17][18] != ele[17][28];
    ele[17][18] != ele[17][29];
    ele[17][18] != ele[17][30];
    ele[17][18] != ele[17][31];
    ele[17][18] != ele[17][32];
    ele[17][18] != ele[17][33];
    ele[17][18] != ele[17][34];
    ele[17][18] != ele[17][35];
    ele[17][18] != ele[18][18];
    ele[17][18] != ele[19][18];
    ele[17][18] != ele[20][18];
    ele[17][18] != ele[21][18];
    ele[17][18] != ele[22][18];
    ele[17][18] != ele[23][18];
    ele[17][18] != ele[24][18];
    ele[17][18] != ele[25][18];
    ele[17][18] != ele[26][18];
    ele[17][18] != ele[27][18];
    ele[17][18] != ele[28][18];
    ele[17][18] != ele[29][18];
    ele[17][18] != ele[30][18];
    ele[17][18] != ele[31][18];
    ele[17][18] != ele[32][18];
    ele[17][18] != ele[33][18];
    ele[17][18] != ele[34][18];
    ele[17][18] != ele[35][18];
    ele[17][19] != ele[17][20];
    ele[17][19] != ele[17][21];
    ele[17][19] != ele[17][22];
    ele[17][19] != ele[17][23];
    ele[17][19] != ele[17][24];
    ele[17][19] != ele[17][25];
    ele[17][19] != ele[17][26];
    ele[17][19] != ele[17][27];
    ele[17][19] != ele[17][28];
    ele[17][19] != ele[17][29];
    ele[17][19] != ele[17][30];
    ele[17][19] != ele[17][31];
    ele[17][19] != ele[17][32];
    ele[17][19] != ele[17][33];
    ele[17][19] != ele[17][34];
    ele[17][19] != ele[17][35];
    ele[17][19] != ele[18][19];
    ele[17][19] != ele[19][19];
    ele[17][19] != ele[20][19];
    ele[17][19] != ele[21][19];
    ele[17][19] != ele[22][19];
    ele[17][19] != ele[23][19];
    ele[17][19] != ele[24][19];
    ele[17][19] != ele[25][19];
    ele[17][19] != ele[26][19];
    ele[17][19] != ele[27][19];
    ele[17][19] != ele[28][19];
    ele[17][19] != ele[29][19];
    ele[17][19] != ele[30][19];
    ele[17][19] != ele[31][19];
    ele[17][19] != ele[32][19];
    ele[17][19] != ele[33][19];
    ele[17][19] != ele[34][19];
    ele[17][19] != ele[35][19];
    ele[17][2] != ele[17][10];
    ele[17][2] != ele[17][11];
    ele[17][2] != ele[17][12];
    ele[17][2] != ele[17][13];
    ele[17][2] != ele[17][14];
    ele[17][2] != ele[17][15];
    ele[17][2] != ele[17][16];
    ele[17][2] != ele[17][17];
    ele[17][2] != ele[17][18];
    ele[17][2] != ele[17][19];
    ele[17][2] != ele[17][20];
    ele[17][2] != ele[17][21];
    ele[17][2] != ele[17][22];
    ele[17][2] != ele[17][23];
    ele[17][2] != ele[17][24];
    ele[17][2] != ele[17][25];
    ele[17][2] != ele[17][26];
    ele[17][2] != ele[17][27];
    ele[17][2] != ele[17][28];
    ele[17][2] != ele[17][29];
    ele[17][2] != ele[17][3];
    ele[17][2] != ele[17][30];
    ele[17][2] != ele[17][31];
    ele[17][2] != ele[17][32];
    ele[17][2] != ele[17][33];
    ele[17][2] != ele[17][34];
    ele[17][2] != ele[17][35];
    ele[17][2] != ele[17][4];
    ele[17][2] != ele[17][5];
    ele[17][2] != ele[17][6];
    ele[17][2] != ele[17][7];
    ele[17][2] != ele[17][8];
    ele[17][2] != ele[17][9];
    ele[17][2] != ele[18][2];
    ele[17][2] != ele[19][2];
    ele[17][2] != ele[20][2];
    ele[17][2] != ele[21][2];
    ele[17][2] != ele[22][2];
    ele[17][2] != ele[23][2];
    ele[17][2] != ele[24][2];
    ele[17][2] != ele[25][2];
    ele[17][2] != ele[26][2];
    ele[17][2] != ele[27][2];
    ele[17][2] != ele[28][2];
    ele[17][2] != ele[29][2];
    ele[17][2] != ele[30][2];
    ele[17][2] != ele[31][2];
    ele[17][2] != ele[32][2];
    ele[17][2] != ele[33][2];
    ele[17][2] != ele[34][2];
    ele[17][2] != ele[35][2];
    ele[17][20] != ele[17][21];
    ele[17][20] != ele[17][22];
    ele[17][20] != ele[17][23];
    ele[17][20] != ele[17][24];
    ele[17][20] != ele[17][25];
    ele[17][20] != ele[17][26];
    ele[17][20] != ele[17][27];
    ele[17][20] != ele[17][28];
    ele[17][20] != ele[17][29];
    ele[17][20] != ele[17][30];
    ele[17][20] != ele[17][31];
    ele[17][20] != ele[17][32];
    ele[17][20] != ele[17][33];
    ele[17][20] != ele[17][34];
    ele[17][20] != ele[17][35];
    ele[17][20] != ele[18][20];
    ele[17][20] != ele[19][20];
    ele[17][20] != ele[20][20];
    ele[17][20] != ele[21][20];
    ele[17][20] != ele[22][20];
    ele[17][20] != ele[23][20];
    ele[17][20] != ele[24][20];
    ele[17][20] != ele[25][20];
    ele[17][20] != ele[26][20];
    ele[17][20] != ele[27][20];
    ele[17][20] != ele[28][20];
    ele[17][20] != ele[29][20];
    ele[17][20] != ele[30][20];
    ele[17][20] != ele[31][20];
    ele[17][20] != ele[32][20];
    ele[17][20] != ele[33][20];
    ele[17][20] != ele[34][20];
    ele[17][20] != ele[35][20];
    ele[17][21] != ele[17][22];
    ele[17][21] != ele[17][23];
    ele[17][21] != ele[17][24];
    ele[17][21] != ele[17][25];
    ele[17][21] != ele[17][26];
    ele[17][21] != ele[17][27];
    ele[17][21] != ele[17][28];
    ele[17][21] != ele[17][29];
    ele[17][21] != ele[17][30];
    ele[17][21] != ele[17][31];
    ele[17][21] != ele[17][32];
    ele[17][21] != ele[17][33];
    ele[17][21] != ele[17][34];
    ele[17][21] != ele[17][35];
    ele[17][21] != ele[18][21];
    ele[17][21] != ele[19][21];
    ele[17][21] != ele[20][21];
    ele[17][21] != ele[21][21];
    ele[17][21] != ele[22][21];
    ele[17][21] != ele[23][21];
    ele[17][21] != ele[24][21];
    ele[17][21] != ele[25][21];
    ele[17][21] != ele[26][21];
    ele[17][21] != ele[27][21];
    ele[17][21] != ele[28][21];
    ele[17][21] != ele[29][21];
    ele[17][21] != ele[30][21];
    ele[17][21] != ele[31][21];
    ele[17][21] != ele[32][21];
    ele[17][21] != ele[33][21];
    ele[17][21] != ele[34][21];
    ele[17][21] != ele[35][21];
    ele[17][22] != ele[17][23];
    ele[17][22] != ele[17][24];
    ele[17][22] != ele[17][25];
    ele[17][22] != ele[17][26];
    ele[17][22] != ele[17][27];
    ele[17][22] != ele[17][28];
    ele[17][22] != ele[17][29];
    ele[17][22] != ele[17][30];
    ele[17][22] != ele[17][31];
    ele[17][22] != ele[17][32];
    ele[17][22] != ele[17][33];
    ele[17][22] != ele[17][34];
    ele[17][22] != ele[17][35];
    ele[17][22] != ele[18][22];
    ele[17][22] != ele[19][22];
    ele[17][22] != ele[20][22];
    ele[17][22] != ele[21][22];
    ele[17][22] != ele[22][22];
    ele[17][22] != ele[23][22];
    ele[17][22] != ele[24][22];
    ele[17][22] != ele[25][22];
    ele[17][22] != ele[26][22];
    ele[17][22] != ele[27][22];
    ele[17][22] != ele[28][22];
    ele[17][22] != ele[29][22];
    ele[17][22] != ele[30][22];
    ele[17][22] != ele[31][22];
    ele[17][22] != ele[32][22];
    ele[17][22] != ele[33][22];
    ele[17][22] != ele[34][22];
    ele[17][22] != ele[35][22];
    ele[17][23] != ele[17][24];
    ele[17][23] != ele[17][25];
    ele[17][23] != ele[17][26];
    ele[17][23] != ele[17][27];
    ele[17][23] != ele[17][28];
    ele[17][23] != ele[17][29];
    ele[17][23] != ele[17][30];
    ele[17][23] != ele[17][31];
    ele[17][23] != ele[17][32];
    ele[17][23] != ele[17][33];
    ele[17][23] != ele[17][34];
    ele[17][23] != ele[17][35];
    ele[17][23] != ele[18][23];
    ele[17][23] != ele[19][23];
    ele[17][23] != ele[20][23];
    ele[17][23] != ele[21][23];
    ele[17][23] != ele[22][23];
    ele[17][23] != ele[23][23];
    ele[17][23] != ele[24][23];
    ele[17][23] != ele[25][23];
    ele[17][23] != ele[26][23];
    ele[17][23] != ele[27][23];
    ele[17][23] != ele[28][23];
    ele[17][23] != ele[29][23];
    ele[17][23] != ele[30][23];
    ele[17][23] != ele[31][23];
    ele[17][23] != ele[32][23];
    ele[17][23] != ele[33][23];
    ele[17][23] != ele[34][23];
    ele[17][23] != ele[35][23];
    ele[17][24] != ele[17][25];
    ele[17][24] != ele[17][26];
    ele[17][24] != ele[17][27];
    ele[17][24] != ele[17][28];
    ele[17][24] != ele[17][29];
    ele[17][24] != ele[17][30];
    ele[17][24] != ele[17][31];
    ele[17][24] != ele[17][32];
    ele[17][24] != ele[17][33];
    ele[17][24] != ele[17][34];
    ele[17][24] != ele[17][35];
    ele[17][24] != ele[18][24];
    ele[17][24] != ele[19][24];
    ele[17][24] != ele[20][24];
    ele[17][24] != ele[21][24];
    ele[17][24] != ele[22][24];
    ele[17][24] != ele[23][24];
    ele[17][24] != ele[24][24];
    ele[17][24] != ele[25][24];
    ele[17][24] != ele[26][24];
    ele[17][24] != ele[27][24];
    ele[17][24] != ele[28][24];
    ele[17][24] != ele[29][24];
    ele[17][24] != ele[30][24];
    ele[17][24] != ele[31][24];
    ele[17][24] != ele[32][24];
    ele[17][24] != ele[33][24];
    ele[17][24] != ele[34][24];
    ele[17][24] != ele[35][24];
    ele[17][25] != ele[17][26];
    ele[17][25] != ele[17][27];
    ele[17][25] != ele[17][28];
    ele[17][25] != ele[17][29];
    ele[17][25] != ele[17][30];
    ele[17][25] != ele[17][31];
    ele[17][25] != ele[17][32];
    ele[17][25] != ele[17][33];
    ele[17][25] != ele[17][34];
    ele[17][25] != ele[17][35];
    ele[17][25] != ele[18][25];
    ele[17][25] != ele[19][25];
    ele[17][25] != ele[20][25];
    ele[17][25] != ele[21][25];
    ele[17][25] != ele[22][25];
    ele[17][25] != ele[23][25];
    ele[17][25] != ele[24][25];
    ele[17][25] != ele[25][25];
    ele[17][25] != ele[26][25];
    ele[17][25] != ele[27][25];
    ele[17][25] != ele[28][25];
    ele[17][25] != ele[29][25];
    ele[17][25] != ele[30][25];
    ele[17][25] != ele[31][25];
    ele[17][25] != ele[32][25];
    ele[17][25] != ele[33][25];
    ele[17][25] != ele[34][25];
    ele[17][25] != ele[35][25];
    ele[17][26] != ele[17][27];
    ele[17][26] != ele[17][28];
    ele[17][26] != ele[17][29];
    ele[17][26] != ele[17][30];
    ele[17][26] != ele[17][31];
    ele[17][26] != ele[17][32];
    ele[17][26] != ele[17][33];
    ele[17][26] != ele[17][34];
    ele[17][26] != ele[17][35];
    ele[17][26] != ele[18][26];
    ele[17][26] != ele[19][26];
    ele[17][26] != ele[20][26];
    ele[17][26] != ele[21][26];
    ele[17][26] != ele[22][26];
    ele[17][26] != ele[23][26];
    ele[17][26] != ele[24][26];
    ele[17][26] != ele[25][26];
    ele[17][26] != ele[26][26];
    ele[17][26] != ele[27][26];
    ele[17][26] != ele[28][26];
    ele[17][26] != ele[29][26];
    ele[17][26] != ele[30][26];
    ele[17][26] != ele[31][26];
    ele[17][26] != ele[32][26];
    ele[17][26] != ele[33][26];
    ele[17][26] != ele[34][26];
    ele[17][26] != ele[35][26];
    ele[17][27] != ele[17][28];
    ele[17][27] != ele[17][29];
    ele[17][27] != ele[17][30];
    ele[17][27] != ele[17][31];
    ele[17][27] != ele[17][32];
    ele[17][27] != ele[17][33];
    ele[17][27] != ele[17][34];
    ele[17][27] != ele[17][35];
    ele[17][27] != ele[18][27];
    ele[17][27] != ele[19][27];
    ele[17][27] != ele[20][27];
    ele[17][27] != ele[21][27];
    ele[17][27] != ele[22][27];
    ele[17][27] != ele[23][27];
    ele[17][27] != ele[24][27];
    ele[17][27] != ele[25][27];
    ele[17][27] != ele[26][27];
    ele[17][27] != ele[27][27];
    ele[17][27] != ele[28][27];
    ele[17][27] != ele[29][27];
    ele[17][27] != ele[30][27];
    ele[17][27] != ele[31][27];
    ele[17][27] != ele[32][27];
    ele[17][27] != ele[33][27];
    ele[17][27] != ele[34][27];
    ele[17][27] != ele[35][27];
    ele[17][28] != ele[17][29];
    ele[17][28] != ele[17][30];
    ele[17][28] != ele[17][31];
    ele[17][28] != ele[17][32];
    ele[17][28] != ele[17][33];
    ele[17][28] != ele[17][34];
    ele[17][28] != ele[17][35];
    ele[17][28] != ele[18][28];
    ele[17][28] != ele[19][28];
    ele[17][28] != ele[20][28];
    ele[17][28] != ele[21][28];
    ele[17][28] != ele[22][28];
    ele[17][28] != ele[23][28];
    ele[17][28] != ele[24][28];
    ele[17][28] != ele[25][28];
    ele[17][28] != ele[26][28];
    ele[17][28] != ele[27][28];
    ele[17][28] != ele[28][28];
    ele[17][28] != ele[29][28];
    ele[17][28] != ele[30][28];
    ele[17][28] != ele[31][28];
    ele[17][28] != ele[32][28];
    ele[17][28] != ele[33][28];
    ele[17][28] != ele[34][28];
    ele[17][28] != ele[35][28];
    ele[17][29] != ele[17][30];
    ele[17][29] != ele[17][31];
    ele[17][29] != ele[17][32];
    ele[17][29] != ele[17][33];
    ele[17][29] != ele[17][34];
    ele[17][29] != ele[17][35];
    ele[17][29] != ele[18][29];
    ele[17][29] != ele[19][29];
    ele[17][29] != ele[20][29];
    ele[17][29] != ele[21][29];
    ele[17][29] != ele[22][29];
    ele[17][29] != ele[23][29];
    ele[17][29] != ele[24][29];
    ele[17][29] != ele[25][29];
    ele[17][29] != ele[26][29];
    ele[17][29] != ele[27][29];
    ele[17][29] != ele[28][29];
    ele[17][29] != ele[29][29];
    ele[17][29] != ele[30][29];
    ele[17][29] != ele[31][29];
    ele[17][29] != ele[32][29];
    ele[17][29] != ele[33][29];
    ele[17][29] != ele[34][29];
    ele[17][29] != ele[35][29];
    ele[17][3] != ele[17][10];
    ele[17][3] != ele[17][11];
    ele[17][3] != ele[17][12];
    ele[17][3] != ele[17][13];
    ele[17][3] != ele[17][14];
    ele[17][3] != ele[17][15];
    ele[17][3] != ele[17][16];
    ele[17][3] != ele[17][17];
    ele[17][3] != ele[17][18];
    ele[17][3] != ele[17][19];
    ele[17][3] != ele[17][20];
    ele[17][3] != ele[17][21];
    ele[17][3] != ele[17][22];
    ele[17][3] != ele[17][23];
    ele[17][3] != ele[17][24];
    ele[17][3] != ele[17][25];
    ele[17][3] != ele[17][26];
    ele[17][3] != ele[17][27];
    ele[17][3] != ele[17][28];
    ele[17][3] != ele[17][29];
    ele[17][3] != ele[17][30];
    ele[17][3] != ele[17][31];
    ele[17][3] != ele[17][32];
    ele[17][3] != ele[17][33];
    ele[17][3] != ele[17][34];
    ele[17][3] != ele[17][35];
    ele[17][3] != ele[17][4];
    ele[17][3] != ele[17][5];
    ele[17][3] != ele[17][6];
    ele[17][3] != ele[17][7];
    ele[17][3] != ele[17][8];
    ele[17][3] != ele[17][9];
    ele[17][3] != ele[18][3];
    ele[17][3] != ele[19][3];
    ele[17][3] != ele[20][3];
    ele[17][3] != ele[21][3];
    ele[17][3] != ele[22][3];
    ele[17][3] != ele[23][3];
    ele[17][3] != ele[24][3];
    ele[17][3] != ele[25][3];
    ele[17][3] != ele[26][3];
    ele[17][3] != ele[27][3];
    ele[17][3] != ele[28][3];
    ele[17][3] != ele[29][3];
    ele[17][3] != ele[30][3];
    ele[17][3] != ele[31][3];
    ele[17][3] != ele[32][3];
    ele[17][3] != ele[33][3];
    ele[17][3] != ele[34][3];
    ele[17][3] != ele[35][3];
    ele[17][30] != ele[17][31];
    ele[17][30] != ele[17][32];
    ele[17][30] != ele[17][33];
    ele[17][30] != ele[17][34];
    ele[17][30] != ele[17][35];
    ele[17][30] != ele[18][30];
    ele[17][30] != ele[19][30];
    ele[17][30] != ele[20][30];
    ele[17][30] != ele[21][30];
    ele[17][30] != ele[22][30];
    ele[17][30] != ele[23][30];
    ele[17][30] != ele[24][30];
    ele[17][30] != ele[25][30];
    ele[17][30] != ele[26][30];
    ele[17][30] != ele[27][30];
    ele[17][30] != ele[28][30];
    ele[17][30] != ele[29][30];
    ele[17][30] != ele[30][30];
    ele[17][30] != ele[31][30];
    ele[17][30] != ele[32][30];
    ele[17][30] != ele[33][30];
    ele[17][30] != ele[34][30];
    ele[17][30] != ele[35][30];
    ele[17][31] != ele[17][32];
    ele[17][31] != ele[17][33];
    ele[17][31] != ele[17][34];
    ele[17][31] != ele[17][35];
    ele[17][31] != ele[18][31];
    ele[17][31] != ele[19][31];
    ele[17][31] != ele[20][31];
    ele[17][31] != ele[21][31];
    ele[17][31] != ele[22][31];
    ele[17][31] != ele[23][31];
    ele[17][31] != ele[24][31];
    ele[17][31] != ele[25][31];
    ele[17][31] != ele[26][31];
    ele[17][31] != ele[27][31];
    ele[17][31] != ele[28][31];
    ele[17][31] != ele[29][31];
    ele[17][31] != ele[30][31];
    ele[17][31] != ele[31][31];
    ele[17][31] != ele[32][31];
    ele[17][31] != ele[33][31];
    ele[17][31] != ele[34][31];
    ele[17][31] != ele[35][31];
    ele[17][32] != ele[17][33];
    ele[17][32] != ele[17][34];
    ele[17][32] != ele[17][35];
    ele[17][32] != ele[18][32];
    ele[17][32] != ele[19][32];
    ele[17][32] != ele[20][32];
    ele[17][32] != ele[21][32];
    ele[17][32] != ele[22][32];
    ele[17][32] != ele[23][32];
    ele[17][32] != ele[24][32];
    ele[17][32] != ele[25][32];
    ele[17][32] != ele[26][32];
    ele[17][32] != ele[27][32];
    ele[17][32] != ele[28][32];
    ele[17][32] != ele[29][32];
    ele[17][32] != ele[30][32];
    ele[17][32] != ele[31][32];
    ele[17][32] != ele[32][32];
    ele[17][32] != ele[33][32];
    ele[17][32] != ele[34][32];
    ele[17][32] != ele[35][32];
    ele[17][33] != ele[17][34];
    ele[17][33] != ele[17][35];
    ele[17][33] != ele[18][33];
    ele[17][33] != ele[19][33];
    ele[17][33] != ele[20][33];
    ele[17][33] != ele[21][33];
    ele[17][33] != ele[22][33];
    ele[17][33] != ele[23][33];
    ele[17][33] != ele[24][33];
    ele[17][33] != ele[25][33];
    ele[17][33] != ele[26][33];
    ele[17][33] != ele[27][33];
    ele[17][33] != ele[28][33];
    ele[17][33] != ele[29][33];
    ele[17][33] != ele[30][33];
    ele[17][33] != ele[31][33];
    ele[17][33] != ele[32][33];
    ele[17][33] != ele[33][33];
    ele[17][33] != ele[34][33];
    ele[17][33] != ele[35][33];
    ele[17][34] != ele[17][35];
    ele[17][34] != ele[18][34];
    ele[17][34] != ele[19][34];
    ele[17][34] != ele[20][34];
    ele[17][34] != ele[21][34];
    ele[17][34] != ele[22][34];
    ele[17][34] != ele[23][34];
    ele[17][34] != ele[24][34];
    ele[17][34] != ele[25][34];
    ele[17][34] != ele[26][34];
    ele[17][34] != ele[27][34];
    ele[17][34] != ele[28][34];
    ele[17][34] != ele[29][34];
    ele[17][34] != ele[30][34];
    ele[17][34] != ele[31][34];
    ele[17][34] != ele[32][34];
    ele[17][34] != ele[33][34];
    ele[17][34] != ele[34][34];
    ele[17][34] != ele[35][34];
    ele[17][35] != ele[18][35];
    ele[17][35] != ele[19][35];
    ele[17][35] != ele[20][35];
    ele[17][35] != ele[21][35];
    ele[17][35] != ele[22][35];
    ele[17][35] != ele[23][35];
    ele[17][35] != ele[24][35];
    ele[17][35] != ele[25][35];
    ele[17][35] != ele[26][35];
    ele[17][35] != ele[27][35];
    ele[17][35] != ele[28][35];
    ele[17][35] != ele[29][35];
    ele[17][35] != ele[30][35];
    ele[17][35] != ele[31][35];
    ele[17][35] != ele[32][35];
    ele[17][35] != ele[33][35];
    ele[17][35] != ele[34][35];
    ele[17][35] != ele[35][35];
    ele[17][4] != ele[17][10];
    ele[17][4] != ele[17][11];
    ele[17][4] != ele[17][12];
    ele[17][4] != ele[17][13];
    ele[17][4] != ele[17][14];
    ele[17][4] != ele[17][15];
    ele[17][4] != ele[17][16];
    ele[17][4] != ele[17][17];
    ele[17][4] != ele[17][18];
    ele[17][4] != ele[17][19];
    ele[17][4] != ele[17][20];
    ele[17][4] != ele[17][21];
    ele[17][4] != ele[17][22];
    ele[17][4] != ele[17][23];
    ele[17][4] != ele[17][24];
    ele[17][4] != ele[17][25];
    ele[17][4] != ele[17][26];
    ele[17][4] != ele[17][27];
    ele[17][4] != ele[17][28];
    ele[17][4] != ele[17][29];
    ele[17][4] != ele[17][30];
    ele[17][4] != ele[17][31];
    ele[17][4] != ele[17][32];
    ele[17][4] != ele[17][33];
    ele[17][4] != ele[17][34];
    ele[17][4] != ele[17][35];
    ele[17][4] != ele[17][5];
    ele[17][4] != ele[17][6];
    ele[17][4] != ele[17][7];
    ele[17][4] != ele[17][8];
    ele[17][4] != ele[17][9];
    ele[17][4] != ele[18][4];
    ele[17][4] != ele[19][4];
    ele[17][4] != ele[20][4];
    ele[17][4] != ele[21][4];
    ele[17][4] != ele[22][4];
    ele[17][4] != ele[23][4];
    ele[17][4] != ele[24][4];
    ele[17][4] != ele[25][4];
    ele[17][4] != ele[26][4];
    ele[17][4] != ele[27][4];
    ele[17][4] != ele[28][4];
    ele[17][4] != ele[29][4];
    ele[17][4] != ele[30][4];
    ele[17][4] != ele[31][4];
    ele[17][4] != ele[32][4];
    ele[17][4] != ele[33][4];
    ele[17][4] != ele[34][4];
    ele[17][4] != ele[35][4];
    ele[17][5] != ele[17][10];
    ele[17][5] != ele[17][11];
    ele[17][5] != ele[17][12];
    ele[17][5] != ele[17][13];
    ele[17][5] != ele[17][14];
    ele[17][5] != ele[17][15];
    ele[17][5] != ele[17][16];
    ele[17][5] != ele[17][17];
    ele[17][5] != ele[17][18];
    ele[17][5] != ele[17][19];
    ele[17][5] != ele[17][20];
    ele[17][5] != ele[17][21];
    ele[17][5] != ele[17][22];
    ele[17][5] != ele[17][23];
    ele[17][5] != ele[17][24];
    ele[17][5] != ele[17][25];
    ele[17][5] != ele[17][26];
    ele[17][5] != ele[17][27];
    ele[17][5] != ele[17][28];
    ele[17][5] != ele[17][29];
    ele[17][5] != ele[17][30];
    ele[17][5] != ele[17][31];
    ele[17][5] != ele[17][32];
    ele[17][5] != ele[17][33];
    ele[17][5] != ele[17][34];
    ele[17][5] != ele[17][35];
    ele[17][5] != ele[17][6];
    ele[17][5] != ele[17][7];
    ele[17][5] != ele[17][8];
    ele[17][5] != ele[17][9];
    ele[17][5] != ele[18][5];
    ele[17][5] != ele[19][5];
    ele[17][5] != ele[20][5];
    ele[17][5] != ele[21][5];
    ele[17][5] != ele[22][5];
    ele[17][5] != ele[23][5];
    ele[17][5] != ele[24][5];
    ele[17][5] != ele[25][5];
    ele[17][5] != ele[26][5];
    ele[17][5] != ele[27][5];
    ele[17][5] != ele[28][5];
    ele[17][5] != ele[29][5];
    ele[17][5] != ele[30][5];
    ele[17][5] != ele[31][5];
    ele[17][5] != ele[32][5];
    ele[17][5] != ele[33][5];
    ele[17][5] != ele[34][5];
    ele[17][5] != ele[35][5];
    ele[17][6] != ele[17][10];
    ele[17][6] != ele[17][11];
    ele[17][6] != ele[17][12];
    ele[17][6] != ele[17][13];
    ele[17][6] != ele[17][14];
    ele[17][6] != ele[17][15];
    ele[17][6] != ele[17][16];
    ele[17][6] != ele[17][17];
    ele[17][6] != ele[17][18];
    ele[17][6] != ele[17][19];
    ele[17][6] != ele[17][20];
    ele[17][6] != ele[17][21];
    ele[17][6] != ele[17][22];
    ele[17][6] != ele[17][23];
    ele[17][6] != ele[17][24];
    ele[17][6] != ele[17][25];
    ele[17][6] != ele[17][26];
    ele[17][6] != ele[17][27];
    ele[17][6] != ele[17][28];
    ele[17][6] != ele[17][29];
    ele[17][6] != ele[17][30];
    ele[17][6] != ele[17][31];
    ele[17][6] != ele[17][32];
    ele[17][6] != ele[17][33];
    ele[17][6] != ele[17][34];
    ele[17][6] != ele[17][35];
    ele[17][6] != ele[17][7];
    ele[17][6] != ele[17][8];
    ele[17][6] != ele[17][9];
    ele[17][6] != ele[18][6];
    ele[17][6] != ele[19][6];
    ele[17][6] != ele[20][6];
    ele[17][6] != ele[21][6];
    ele[17][6] != ele[22][6];
    ele[17][6] != ele[23][6];
    ele[17][6] != ele[24][6];
    ele[17][6] != ele[25][6];
    ele[17][6] != ele[26][6];
    ele[17][6] != ele[27][6];
    ele[17][6] != ele[28][6];
    ele[17][6] != ele[29][6];
    ele[17][6] != ele[30][6];
    ele[17][6] != ele[31][6];
    ele[17][6] != ele[32][6];
    ele[17][6] != ele[33][6];
    ele[17][6] != ele[34][6];
    ele[17][6] != ele[35][6];
    ele[17][7] != ele[17][10];
    ele[17][7] != ele[17][11];
    ele[17][7] != ele[17][12];
    ele[17][7] != ele[17][13];
    ele[17][7] != ele[17][14];
    ele[17][7] != ele[17][15];
    ele[17][7] != ele[17][16];
    ele[17][7] != ele[17][17];
    ele[17][7] != ele[17][18];
    ele[17][7] != ele[17][19];
    ele[17][7] != ele[17][20];
    ele[17][7] != ele[17][21];
    ele[17][7] != ele[17][22];
    ele[17][7] != ele[17][23];
    ele[17][7] != ele[17][24];
    ele[17][7] != ele[17][25];
    ele[17][7] != ele[17][26];
    ele[17][7] != ele[17][27];
    ele[17][7] != ele[17][28];
    ele[17][7] != ele[17][29];
    ele[17][7] != ele[17][30];
    ele[17][7] != ele[17][31];
    ele[17][7] != ele[17][32];
    ele[17][7] != ele[17][33];
    ele[17][7] != ele[17][34];
    ele[17][7] != ele[17][35];
    ele[17][7] != ele[17][8];
    ele[17][7] != ele[17][9];
    ele[17][7] != ele[18][7];
    ele[17][7] != ele[19][7];
    ele[17][7] != ele[20][7];
    ele[17][7] != ele[21][7];
    ele[17][7] != ele[22][7];
    ele[17][7] != ele[23][7];
    ele[17][7] != ele[24][7];
    ele[17][7] != ele[25][7];
    ele[17][7] != ele[26][7];
    ele[17][7] != ele[27][7];
    ele[17][7] != ele[28][7];
    ele[17][7] != ele[29][7];
    ele[17][7] != ele[30][7];
    ele[17][7] != ele[31][7];
    ele[17][7] != ele[32][7];
    ele[17][7] != ele[33][7];
    ele[17][7] != ele[34][7];
    ele[17][7] != ele[35][7];
    ele[17][8] != ele[17][10];
    ele[17][8] != ele[17][11];
    ele[17][8] != ele[17][12];
    ele[17][8] != ele[17][13];
    ele[17][8] != ele[17][14];
    ele[17][8] != ele[17][15];
    ele[17][8] != ele[17][16];
    ele[17][8] != ele[17][17];
    ele[17][8] != ele[17][18];
    ele[17][8] != ele[17][19];
    ele[17][8] != ele[17][20];
    ele[17][8] != ele[17][21];
    ele[17][8] != ele[17][22];
    ele[17][8] != ele[17][23];
    ele[17][8] != ele[17][24];
    ele[17][8] != ele[17][25];
    ele[17][8] != ele[17][26];
    ele[17][8] != ele[17][27];
    ele[17][8] != ele[17][28];
    ele[17][8] != ele[17][29];
    ele[17][8] != ele[17][30];
    ele[17][8] != ele[17][31];
    ele[17][8] != ele[17][32];
    ele[17][8] != ele[17][33];
    ele[17][8] != ele[17][34];
    ele[17][8] != ele[17][35];
    ele[17][8] != ele[17][9];
    ele[17][8] != ele[18][8];
    ele[17][8] != ele[19][8];
    ele[17][8] != ele[20][8];
    ele[17][8] != ele[21][8];
    ele[17][8] != ele[22][8];
    ele[17][8] != ele[23][8];
    ele[17][8] != ele[24][8];
    ele[17][8] != ele[25][8];
    ele[17][8] != ele[26][8];
    ele[17][8] != ele[27][8];
    ele[17][8] != ele[28][8];
    ele[17][8] != ele[29][8];
    ele[17][8] != ele[30][8];
    ele[17][8] != ele[31][8];
    ele[17][8] != ele[32][8];
    ele[17][8] != ele[33][8];
    ele[17][8] != ele[34][8];
    ele[17][8] != ele[35][8];
    ele[17][9] != ele[17][10];
    ele[17][9] != ele[17][11];
    ele[17][9] != ele[17][12];
    ele[17][9] != ele[17][13];
    ele[17][9] != ele[17][14];
    ele[17][9] != ele[17][15];
    ele[17][9] != ele[17][16];
    ele[17][9] != ele[17][17];
    ele[17][9] != ele[17][18];
    ele[17][9] != ele[17][19];
    ele[17][9] != ele[17][20];
    ele[17][9] != ele[17][21];
    ele[17][9] != ele[17][22];
    ele[17][9] != ele[17][23];
    ele[17][9] != ele[17][24];
    ele[17][9] != ele[17][25];
    ele[17][9] != ele[17][26];
    ele[17][9] != ele[17][27];
    ele[17][9] != ele[17][28];
    ele[17][9] != ele[17][29];
    ele[17][9] != ele[17][30];
    ele[17][9] != ele[17][31];
    ele[17][9] != ele[17][32];
    ele[17][9] != ele[17][33];
    ele[17][9] != ele[17][34];
    ele[17][9] != ele[17][35];
    ele[17][9] != ele[18][9];
    ele[17][9] != ele[19][9];
    ele[17][9] != ele[20][9];
    ele[17][9] != ele[21][9];
    ele[17][9] != ele[22][9];
    ele[17][9] != ele[23][9];
    ele[17][9] != ele[24][9];
    ele[17][9] != ele[25][9];
    ele[17][9] != ele[26][9];
    ele[17][9] != ele[27][9];
    ele[17][9] != ele[28][9];
    ele[17][9] != ele[29][9];
    ele[17][9] != ele[30][9];
    ele[17][9] != ele[31][9];
    ele[17][9] != ele[32][9];
    ele[17][9] != ele[33][9];
    ele[17][9] != ele[34][9];
    ele[17][9] != ele[35][9];
    ele[18][0] != ele[18][1];
    ele[18][0] != ele[18][10];
    ele[18][0] != ele[18][11];
    ele[18][0] != ele[18][12];
    ele[18][0] != ele[18][13];
    ele[18][0] != ele[18][14];
    ele[18][0] != ele[18][15];
    ele[18][0] != ele[18][16];
    ele[18][0] != ele[18][17];
    ele[18][0] != ele[18][18];
    ele[18][0] != ele[18][19];
    ele[18][0] != ele[18][2];
    ele[18][0] != ele[18][20];
    ele[18][0] != ele[18][21];
    ele[18][0] != ele[18][22];
    ele[18][0] != ele[18][23];
    ele[18][0] != ele[18][24];
    ele[18][0] != ele[18][25];
    ele[18][0] != ele[18][26];
    ele[18][0] != ele[18][27];
    ele[18][0] != ele[18][28];
    ele[18][0] != ele[18][29];
    ele[18][0] != ele[18][3];
    ele[18][0] != ele[18][30];
    ele[18][0] != ele[18][31];
    ele[18][0] != ele[18][32];
    ele[18][0] != ele[18][33];
    ele[18][0] != ele[18][34];
    ele[18][0] != ele[18][35];
    ele[18][0] != ele[18][4];
    ele[18][0] != ele[18][5];
    ele[18][0] != ele[18][6];
    ele[18][0] != ele[18][7];
    ele[18][0] != ele[18][8];
    ele[18][0] != ele[18][9];
    ele[18][0] != ele[19][0];
    ele[18][0] != ele[19][1];
    ele[18][0] != ele[19][2];
    ele[18][0] != ele[19][3];
    ele[18][0] != ele[19][4];
    ele[18][0] != ele[19][5];
    ele[18][0] != ele[20][0];
    ele[18][0] != ele[20][1];
    ele[18][0] != ele[20][2];
    ele[18][0] != ele[20][3];
    ele[18][0] != ele[20][4];
    ele[18][0] != ele[20][5];
    ele[18][0] != ele[21][0];
    ele[18][0] != ele[21][1];
    ele[18][0] != ele[21][2];
    ele[18][0] != ele[21][3];
    ele[18][0] != ele[21][4];
    ele[18][0] != ele[21][5];
    ele[18][0] != ele[22][0];
    ele[18][0] != ele[22][1];
    ele[18][0] != ele[22][2];
    ele[18][0] != ele[22][3];
    ele[18][0] != ele[22][4];
    ele[18][0] != ele[22][5];
    ele[18][0] != ele[23][0];
    ele[18][0] != ele[23][1];
    ele[18][0] != ele[23][2];
    ele[18][0] != ele[23][3];
    ele[18][0] != ele[23][4];
    ele[18][0] != ele[23][5];
    ele[18][0] != ele[24][0];
    ele[18][0] != ele[25][0];
    ele[18][0] != ele[26][0];
    ele[18][0] != ele[27][0];
    ele[18][0] != ele[28][0];
    ele[18][0] != ele[29][0];
    ele[18][0] != ele[30][0];
    ele[18][0] != ele[31][0];
    ele[18][0] != ele[32][0];
    ele[18][0] != ele[33][0];
    ele[18][0] != ele[34][0];
    ele[18][0] != ele[35][0];
    ele[18][1] != ele[18][10];
    ele[18][1] != ele[18][11];
    ele[18][1] != ele[18][12];
    ele[18][1] != ele[18][13];
    ele[18][1] != ele[18][14];
    ele[18][1] != ele[18][15];
    ele[18][1] != ele[18][16];
    ele[18][1] != ele[18][17];
    ele[18][1] != ele[18][18];
    ele[18][1] != ele[18][19];
    ele[18][1] != ele[18][2];
    ele[18][1] != ele[18][20];
    ele[18][1] != ele[18][21];
    ele[18][1] != ele[18][22];
    ele[18][1] != ele[18][23];
    ele[18][1] != ele[18][24];
    ele[18][1] != ele[18][25];
    ele[18][1] != ele[18][26];
    ele[18][1] != ele[18][27];
    ele[18][1] != ele[18][28];
    ele[18][1] != ele[18][29];
    ele[18][1] != ele[18][3];
    ele[18][1] != ele[18][30];
    ele[18][1] != ele[18][31];
    ele[18][1] != ele[18][32];
    ele[18][1] != ele[18][33];
    ele[18][1] != ele[18][34];
    ele[18][1] != ele[18][35];
    ele[18][1] != ele[18][4];
    ele[18][1] != ele[18][5];
    ele[18][1] != ele[18][6];
    ele[18][1] != ele[18][7];
    ele[18][1] != ele[18][8];
    ele[18][1] != ele[18][9];
    ele[18][1] != ele[19][0];
    ele[18][1] != ele[19][1];
    ele[18][1] != ele[19][2];
    ele[18][1] != ele[19][3];
    ele[18][1] != ele[19][4];
    ele[18][1] != ele[19][5];
    ele[18][1] != ele[20][0];
    ele[18][1] != ele[20][1];
    ele[18][1] != ele[20][2];
    ele[18][1] != ele[20][3];
    ele[18][1] != ele[20][4];
    ele[18][1] != ele[20][5];
    ele[18][1] != ele[21][0];
    ele[18][1] != ele[21][1];
    ele[18][1] != ele[21][2];
    ele[18][1] != ele[21][3];
    ele[18][1] != ele[21][4];
    ele[18][1] != ele[21][5];
    ele[18][1] != ele[22][0];
    ele[18][1] != ele[22][1];
    ele[18][1] != ele[22][2];
    ele[18][1] != ele[22][3];
    ele[18][1] != ele[22][4];
    ele[18][1] != ele[22][5];
    ele[18][1] != ele[23][0];
    ele[18][1] != ele[23][1];
    ele[18][1] != ele[23][2];
    ele[18][1] != ele[23][3];
    ele[18][1] != ele[23][4];
    ele[18][1] != ele[23][5];
    ele[18][1] != ele[24][1];
    ele[18][1] != ele[25][1];
    ele[18][1] != ele[26][1];
    ele[18][1] != ele[27][1];
    ele[18][1] != ele[28][1];
    ele[18][1] != ele[29][1];
    ele[18][1] != ele[30][1];
    ele[18][1] != ele[31][1];
    ele[18][1] != ele[32][1];
    ele[18][1] != ele[33][1];
    ele[18][1] != ele[34][1];
    ele[18][1] != ele[35][1];
    ele[18][10] != ele[18][11];
    ele[18][10] != ele[18][12];
    ele[18][10] != ele[18][13];
    ele[18][10] != ele[18][14];
    ele[18][10] != ele[18][15];
    ele[18][10] != ele[18][16];
    ele[18][10] != ele[18][17];
    ele[18][10] != ele[18][18];
    ele[18][10] != ele[18][19];
    ele[18][10] != ele[18][20];
    ele[18][10] != ele[18][21];
    ele[18][10] != ele[18][22];
    ele[18][10] != ele[18][23];
    ele[18][10] != ele[18][24];
    ele[18][10] != ele[18][25];
    ele[18][10] != ele[18][26];
    ele[18][10] != ele[18][27];
    ele[18][10] != ele[18][28];
    ele[18][10] != ele[18][29];
    ele[18][10] != ele[18][30];
    ele[18][10] != ele[18][31];
    ele[18][10] != ele[18][32];
    ele[18][10] != ele[18][33];
    ele[18][10] != ele[18][34];
    ele[18][10] != ele[18][35];
    ele[18][10] != ele[19][10];
    ele[18][10] != ele[19][11];
    ele[18][10] != ele[19][6];
    ele[18][10] != ele[19][7];
    ele[18][10] != ele[19][8];
    ele[18][10] != ele[19][9];
    ele[18][10] != ele[20][10];
    ele[18][10] != ele[20][11];
    ele[18][10] != ele[20][6];
    ele[18][10] != ele[20][7];
    ele[18][10] != ele[20][8];
    ele[18][10] != ele[20][9];
    ele[18][10] != ele[21][10];
    ele[18][10] != ele[21][11];
    ele[18][10] != ele[21][6];
    ele[18][10] != ele[21][7];
    ele[18][10] != ele[21][8];
    ele[18][10] != ele[21][9];
    ele[18][10] != ele[22][10];
    ele[18][10] != ele[22][11];
    ele[18][10] != ele[22][6];
    ele[18][10] != ele[22][7];
    ele[18][10] != ele[22][8];
    ele[18][10] != ele[22][9];
    ele[18][10] != ele[23][10];
    ele[18][10] != ele[23][11];
    ele[18][10] != ele[23][6];
    ele[18][10] != ele[23][7];
    ele[18][10] != ele[23][8];
    ele[18][10] != ele[23][9];
    ele[18][10] != ele[24][10];
    ele[18][10] != ele[25][10];
    ele[18][10] != ele[26][10];
    ele[18][10] != ele[27][10];
    ele[18][10] != ele[28][10];
    ele[18][10] != ele[29][10];
    ele[18][10] != ele[30][10];
    ele[18][10] != ele[31][10];
    ele[18][10] != ele[32][10];
    ele[18][10] != ele[33][10];
    ele[18][10] != ele[34][10];
    ele[18][10] != ele[35][10];
    ele[18][11] != ele[18][12];
    ele[18][11] != ele[18][13];
    ele[18][11] != ele[18][14];
    ele[18][11] != ele[18][15];
    ele[18][11] != ele[18][16];
    ele[18][11] != ele[18][17];
    ele[18][11] != ele[18][18];
    ele[18][11] != ele[18][19];
    ele[18][11] != ele[18][20];
    ele[18][11] != ele[18][21];
    ele[18][11] != ele[18][22];
    ele[18][11] != ele[18][23];
    ele[18][11] != ele[18][24];
    ele[18][11] != ele[18][25];
    ele[18][11] != ele[18][26];
    ele[18][11] != ele[18][27];
    ele[18][11] != ele[18][28];
    ele[18][11] != ele[18][29];
    ele[18][11] != ele[18][30];
    ele[18][11] != ele[18][31];
    ele[18][11] != ele[18][32];
    ele[18][11] != ele[18][33];
    ele[18][11] != ele[18][34];
    ele[18][11] != ele[18][35];
    ele[18][11] != ele[19][10];
    ele[18][11] != ele[19][11];
    ele[18][11] != ele[19][6];
    ele[18][11] != ele[19][7];
    ele[18][11] != ele[19][8];
    ele[18][11] != ele[19][9];
    ele[18][11] != ele[20][10];
    ele[18][11] != ele[20][11];
    ele[18][11] != ele[20][6];
    ele[18][11] != ele[20][7];
    ele[18][11] != ele[20][8];
    ele[18][11] != ele[20][9];
    ele[18][11] != ele[21][10];
    ele[18][11] != ele[21][11];
    ele[18][11] != ele[21][6];
    ele[18][11] != ele[21][7];
    ele[18][11] != ele[21][8];
    ele[18][11] != ele[21][9];
    ele[18][11] != ele[22][10];
    ele[18][11] != ele[22][11];
    ele[18][11] != ele[22][6];
    ele[18][11] != ele[22][7];
    ele[18][11] != ele[22][8];
    ele[18][11] != ele[22][9];
    ele[18][11] != ele[23][10];
    ele[18][11] != ele[23][11];
    ele[18][11] != ele[23][6];
    ele[18][11] != ele[23][7];
    ele[18][11] != ele[23][8];
    ele[18][11] != ele[23][9];
    ele[18][11] != ele[24][11];
    ele[18][11] != ele[25][11];
    ele[18][11] != ele[26][11];
    ele[18][11] != ele[27][11];
    ele[18][11] != ele[28][11];
    ele[18][11] != ele[29][11];
    ele[18][11] != ele[30][11];
    ele[18][11] != ele[31][11];
    ele[18][11] != ele[32][11];
    ele[18][11] != ele[33][11];
    ele[18][11] != ele[34][11];
    ele[18][11] != ele[35][11];
    ele[18][12] != ele[18][13];
    ele[18][12] != ele[18][14];
    ele[18][12] != ele[18][15];
    ele[18][12] != ele[18][16];
    ele[18][12] != ele[18][17];
    ele[18][12] != ele[18][18];
    ele[18][12] != ele[18][19];
    ele[18][12] != ele[18][20];
    ele[18][12] != ele[18][21];
    ele[18][12] != ele[18][22];
    ele[18][12] != ele[18][23];
    ele[18][12] != ele[18][24];
    ele[18][12] != ele[18][25];
    ele[18][12] != ele[18][26];
    ele[18][12] != ele[18][27];
    ele[18][12] != ele[18][28];
    ele[18][12] != ele[18][29];
    ele[18][12] != ele[18][30];
    ele[18][12] != ele[18][31];
    ele[18][12] != ele[18][32];
    ele[18][12] != ele[18][33];
    ele[18][12] != ele[18][34];
    ele[18][12] != ele[18][35];
    ele[18][12] != ele[19][12];
    ele[18][12] != ele[19][13];
    ele[18][12] != ele[19][14];
    ele[18][12] != ele[19][15];
    ele[18][12] != ele[19][16];
    ele[18][12] != ele[19][17];
    ele[18][12] != ele[20][12];
    ele[18][12] != ele[20][13];
    ele[18][12] != ele[20][14];
    ele[18][12] != ele[20][15];
    ele[18][12] != ele[20][16];
    ele[18][12] != ele[20][17];
    ele[18][12] != ele[21][12];
    ele[18][12] != ele[21][13];
    ele[18][12] != ele[21][14];
    ele[18][12] != ele[21][15];
    ele[18][12] != ele[21][16];
    ele[18][12] != ele[21][17];
    ele[18][12] != ele[22][12];
    ele[18][12] != ele[22][13];
    ele[18][12] != ele[22][14];
    ele[18][12] != ele[22][15];
    ele[18][12] != ele[22][16];
    ele[18][12] != ele[22][17];
    ele[18][12] != ele[23][12];
    ele[18][12] != ele[23][13];
    ele[18][12] != ele[23][14];
    ele[18][12] != ele[23][15];
    ele[18][12] != ele[23][16];
    ele[18][12] != ele[23][17];
    ele[18][12] != ele[24][12];
    ele[18][12] != ele[25][12];
    ele[18][12] != ele[26][12];
    ele[18][12] != ele[27][12];
    ele[18][12] != ele[28][12];
    ele[18][12] != ele[29][12];
    ele[18][12] != ele[30][12];
    ele[18][12] != ele[31][12];
    ele[18][12] != ele[32][12];
    ele[18][12] != ele[33][12];
    ele[18][12] != ele[34][12];
    ele[18][12] != ele[35][12];
    ele[18][13] != ele[18][14];
    ele[18][13] != ele[18][15];
    ele[18][13] != ele[18][16];
    ele[18][13] != ele[18][17];
    ele[18][13] != ele[18][18];
    ele[18][13] != ele[18][19];
    ele[18][13] != ele[18][20];
    ele[18][13] != ele[18][21];
    ele[18][13] != ele[18][22];
    ele[18][13] != ele[18][23];
    ele[18][13] != ele[18][24];
    ele[18][13] != ele[18][25];
    ele[18][13] != ele[18][26];
    ele[18][13] != ele[18][27];
    ele[18][13] != ele[18][28];
    ele[18][13] != ele[18][29];
    ele[18][13] != ele[18][30];
    ele[18][13] != ele[18][31];
    ele[18][13] != ele[18][32];
    ele[18][13] != ele[18][33];
    ele[18][13] != ele[18][34];
    ele[18][13] != ele[18][35];
    ele[18][13] != ele[19][12];
    ele[18][13] != ele[19][13];
    ele[18][13] != ele[19][14];
    ele[18][13] != ele[19][15];
    ele[18][13] != ele[19][16];
    ele[18][13] != ele[19][17];
    ele[18][13] != ele[20][12];
    ele[18][13] != ele[20][13];
    ele[18][13] != ele[20][14];
    ele[18][13] != ele[20][15];
    ele[18][13] != ele[20][16];
    ele[18][13] != ele[20][17];
    ele[18][13] != ele[21][12];
    ele[18][13] != ele[21][13];
    ele[18][13] != ele[21][14];
    ele[18][13] != ele[21][15];
    ele[18][13] != ele[21][16];
    ele[18][13] != ele[21][17];
    ele[18][13] != ele[22][12];
    ele[18][13] != ele[22][13];
    ele[18][13] != ele[22][14];
    ele[18][13] != ele[22][15];
    ele[18][13] != ele[22][16];
    ele[18][13] != ele[22][17];
    ele[18][13] != ele[23][12];
    ele[18][13] != ele[23][13];
    ele[18][13] != ele[23][14];
    ele[18][13] != ele[23][15];
    ele[18][13] != ele[23][16];
    ele[18][13] != ele[23][17];
    ele[18][13] != ele[24][13];
    ele[18][13] != ele[25][13];
    ele[18][13] != ele[26][13];
    ele[18][13] != ele[27][13];
    ele[18][13] != ele[28][13];
    ele[18][13] != ele[29][13];
    ele[18][13] != ele[30][13];
    ele[18][13] != ele[31][13];
    ele[18][13] != ele[32][13];
    ele[18][13] != ele[33][13];
    ele[18][13] != ele[34][13];
    ele[18][13] != ele[35][13];
    ele[18][14] != ele[18][15];
    ele[18][14] != ele[18][16];
    ele[18][14] != ele[18][17];
    ele[18][14] != ele[18][18];
    ele[18][14] != ele[18][19];
    ele[18][14] != ele[18][20];
    ele[18][14] != ele[18][21];
    ele[18][14] != ele[18][22];
    ele[18][14] != ele[18][23];
    ele[18][14] != ele[18][24];
    ele[18][14] != ele[18][25];
    ele[18][14] != ele[18][26];
    ele[18][14] != ele[18][27];
    ele[18][14] != ele[18][28];
    ele[18][14] != ele[18][29];
    ele[18][14] != ele[18][30];
    ele[18][14] != ele[18][31];
    ele[18][14] != ele[18][32];
    ele[18][14] != ele[18][33];
    ele[18][14] != ele[18][34];
    ele[18][14] != ele[18][35];
    ele[18][14] != ele[19][12];
    ele[18][14] != ele[19][13];
    ele[18][14] != ele[19][14];
    ele[18][14] != ele[19][15];
    ele[18][14] != ele[19][16];
    ele[18][14] != ele[19][17];
    ele[18][14] != ele[20][12];
    ele[18][14] != ele[20][13];
    ele[18][14] != ele[20][14];
    ele[18][14] != ele[20][15];
    ele[18][14] != ele[20][16];
    ele[18][14] != ele[20][17];
    ele[18][14] != ele[21][12];
    ele[18][14] != ele[21][13];
    ele[18][14] != ele[21][14];
    ele[18][14] != ele[21][15];
    ele[18][14] != ele[21][16];
    ele[18][14] != ele[21][17];
    ele[18][14] != ele[22][12];
    ele[18][14] != ele[22][13];
    ele[18][14] != ele[22][14];
    ele[18][14] != ele[22][15];
    ele[18][14] != ele[22][16];
    ele[18][14] != ele[22][17];
    ele[18][14] != ele[23][12];
    ele[18][14] != ele[23][13];
    ele[18][14] != ele[23][14];
    ele[18][14] != ele[23][15];
    ele[18][14] != ele[23][16];
    ele[18][14] != ele[23][17];
    ele[18][14] != ele[24][14];
    ele[18][14] != ele[25][14];
    ele[18][14] != ele[26][14];
    ele[18][14] != ele[27][14];
    ele[18][14] != ele[28][14];
    ele[18][14] != ele[29][14];
    ele[18][14] != ele[30][14];
    ele[18][14] != ele[31][14];
    ele[18][14] != ele[32][14];
    ele[18][14] != ele[33][14];
    ele[18][14] != ele[34][14];
    ele[18][14] != ele[35][14];
    ele[18][15] != ele[18][16];
    ele[18][15] != ele[18][17];
    ele[18][15] != ele[18][18];
    ele[18][15] != ele[18][19];
    ele[18][15] != ele[18][20];
    ele[18][15] != ele[18][21];
    ele[18][15] != ele[18][22];
    ele[18][15] != ele[18][23];
    ele[18][15] != ele[18][24];
    ele[18][15] != ele[18][25];
    ele[18][15] != ele[18][26];
    ele[18][15] != ele[18][27];
    ele[18][15] != ele[18][28];
    ele[18][15] != ele[18][29];
    ele[18][15] != ele[18][30];
    ele[18][15] != ele[18][31];
    ele[18][15] != ele[18][32];
    ele[18][15] != ele[18][33];
    ele[18][15] != ele[18][34];
    ele[18][15] != ele[18][35];
    ele[18][15] != ele[19][12];
    ele[18][15] != ele[19][13];
    ele[18][15] != ele[19][14];
    ele[18][15] != ele[19][15];
    ele[18][15] != ele[19][16];
    ele[18][15] != ele[19][17];
    ele[18][15] != ele[20][12];
    ele[18][15] != ele[20][13];
    ele[18][15] != ele[20][14];
    ele[18][15] != ele[20][15];
    ele[18][15] != ele[20][16];
    ele[18][15] != ele[20][17];
    ele[18][15] != ele[21][12];
    ele[18][15] != ele[21][13];
    ele[18][15] != ele[21][14];
    ele[18][15] != ele[21][15];
    ele[18][15] != ele[21][16];
    ele[18][15] != ele[21][17];
    ele[18][15] != ele[22][12];
    ele[18][15] != ele[22][13];
    ele[18][15] != ele[22][14];
    ele[18][15] != ele[22][15];
    ele[18][15] != ele[22][16];
    ele[18][15] != ele[22][17];
    ele[18][15] != ele[23][12];
    ele[18][15] != ele[23][13];
    ele[18][15] != ele[23][14];
    ele[18][15] != ele[23][15];
    ele[18][15] != ele[23][16];
    ele[18][15] != ele[23][17];
    ele[18][15] != ele[24][15];
    ele[18][15] != ele[25][15];
    ele[18][15] != ele[26][15];
    ele[18][15] != ele[27][15];
    ele[18][15] != ele[28][15];
    ele[18][15] != ele[29][15];
    ele[18][15] != ele[30][15];
    ele[18][15] != ele[31][15];
    ele[18][15] != ele[32][15];
    ele[18][15] != ele[33][15];
    ele[18][15] != ele[34][15];
    ele[18][15] != ele[35][15];
    ele[18][16] != ele[18][17];
    ele[18][16] != ele[18][18];
    ele[18][16] != ele[18][19];
    ele[18][16] != ele[18][20];
    ele[18][16] != ele[18][21];
    ele[18][16] != ele[18][22];
    ele[18][16] != ele[18][23];
    ele[18][16] != ele[18][24];
    ele[18][16] != ele[18][25];
    ele[18][16] != ele[18][26];
    ele[18][16] != ele[18][27];
    ele[18][16] != ele[18][28];
    ele[18][16] != ele[18][29];
    ele[18][16] != ele[18][30];
    ele[18][16] != ele[18][31];
    ele[18][16] != ele[18][32];
    ele[18][16] != ele[18][33];
    ele[18][16] != ele[18][34];
    ele[18][16] != ele[18][35];
    ele[18][16] != ele[19][12];
    ele[18][16] != ele[19][13];
    ele[18][16] != ele[19][14];
    ele[18][16] != ele[19][15];
    ele[18][16] != ele[19][16];
    ele[18][16] != ele[19][17];
    ele[18][16] != ele[20][12];
    ele[18][16] != ele[20][13];
    ele[18][16] != ele[20][14];
    ele[18][16] != ele[20][15];
    ele[18][16] != ele[20][16];
    ele[18][16] != ele[20][17];
    ele[18][16] != ele[21][12];
    ele[18][16] != ele[21][13];
    ele[18][16] != ele[21][14];
    ele[18][16] != ele[21][15];
    ele[18][16] != ele[21][16];
    ele[18][16] != ele[21][17];
    ele[18][16] != ele[22][12];
    ele[18][16] != ele[22][13];
    ele[18][16] != ele[22][14];
    ele[18][16] != ele[22][15];
    ele[18][16] != ele[22][16];
    ele[18][16] != ele[22][17];
    ele[18][16] != ele[23][12];
    ele[18][16] != ele[23][13];
    ele[18][16] != ele[23][14];
    ele[18][16] != ele[23][15];
    ele[18][16] != ele[23][16];
    ele[18][16] != ele[23][17];
    ele[18][16] != ele[24][16];
    ele[18][16] != ele[25][16];
    ele[18][16] != ele[26][16];
    ele[18][16] != ele[27][16];
    ele[18][16] != ele[28][16];
    ele[18][16] != ele[29][16];
    ele[18][16] != ele[30][16];
    ele[18][16] != ele[31][16];
    ele[18][16] != ele[32][16];
    ele[18][16] != ele[33][16];
    ele[18][16] != ele[34][16];
    ele[18][16] != ele[35][16];
    ele[18][17] != ele[18][18];
    ele[18][17] != ele[18][19];
    ele[18][17] != ele[18][20];
    ele[18][17] != ele[18][21];
    ele[18][17] != ele[18][22];
    ele[18][17] != ele[18][23];
    ele[18][17] != ele[18][24];
    ele[18][17] != ele[18][25];
    ele[18][17] != ele[18][26];
    ele[18][17] != ele[18][27];
    ele[18][17] != ele[18][28];
    ele[18][17] != ele[18][29];
    ele[18][17] != ele[18][30];
    ele[18][17] != ele[18][31];
    ele[18][17] != ele[18][32];
    ele[18][17] != ele[18][33];
    ele[18][17] != ele[18][34];
    ele[18][17] != ele[18][35];
    ele[18][17] != ele[19][12];
    ele[18][17] != ele[19][13];
    ele[18][17] != ele[19][14];
    ele[18][17] != ele[19][15];
    ele[18][17] != ele[19][16];
    ele[18][17] != ele[19][17];
    ele[18][17] != ele[20][12];
    ele[18][17] != ele[20][13];
    ele[18][17] != ele[20][14];
    ele[18][17] != ele[20][15];
    ele[18][17] != ele[20][16];
    ele[18][17] != ele[20][17];
    ele[18][17] != ele[21][12];
    ele[18][17] != ele[21][13];
    ele[18][17] != ele[21][14];
    ele[18][17] != ele[21][15];
    ele[18][17] != ele[21][16];
    ele[18][17] != ele[21][17];
    ele[18][17] != ele[22][12];
    ele[18][17] != ele[22][13];
    ele[18][17] != ele[22][14];
    ele[18][17] != ele[22][15];
    ele[18][17] != ele[22][16];
    ele[18][17] != ele[22][17];
    ele[18][17] != ele[23][12];
    ele[18][17] != ele[23][13];
    ele[18][17] != ele[23][14];
    ele[18][17] != ele[23][15];
    ele[18][17] != ele[23][16];
    ele[18][17] != ele[23][17];
    ele[18][17] != ele[24][17];
    ele[18][17] != ele[25][17];
    ele[18][17] != ele[26][17];
    ele[18][17] != ele[27][17];
    ele[18][17] != ele[28][17];
    ele[18][17] != ele[29][17];
    ele[18][17] != ele[30][17];
    ele[18][17] != ele[31][17];
    ele[18][17] != ele[32][17];
    ele[18][17] != ele[33][17];
    ele[18][17] != ele[34][17];
    ele[18][17] != ele[35][17];
    ele[18][18] != ele[18][19];
    ele[18][18] != ele[18][20];
    ele[18][18] != ele[18][21];
    ele[18][18] != ele[18][22];
    ele[18][18] != ele[18][23];
    ele[18][18] != ele[18][24];
    ele[18][18] != ele[18][25];
    ele[18][18] != ele[18][26];
    ele[18][18] != ele[18][27];
    ele[18][18] != ele[18][28];
    ele[18][18] != ele[18][29];
    ele[18][18] != ele[18][30];
    ele[18][18] != ele[18][31];
    ele[18][18] != ele[18][32];
    ele[18][18] != ele[18][33];
    ele[18][18] != ele[18][34];
    ele[18][18] != ele[18][35];
    ele[18][18] != ele[19][18];
    ele[18][18] != ele[19][19];
    ele[18][18] != ele[19][20];
    ele[18][18] != ele[19][21];
    ele[18][18] != ele[19][22];
    ele[18][18] != ele[19][23];
    ele[18][18] != ele[20][18];
    ele[18][18] != ele[20][19];
    ele[18][18] != ele[20][20];
    ele[18][18] != ele[20][21];
    ele[18][18] != ele[20][22];
    ele[18][18] != ele[20][23];
    ele[18][18] != ele[21][18];
    ele[18][18] != ele[21][19];
    ele[18][18] != ele[21][20];
    ele[18][18] != ele[21][21];
    ele[18][18] != ele[21][22];
    ele[18][18] != ele[21][23];
    ele[18][18] != ele[22][18];
    ele[18][18] != ele[22][19];
    ele[18][18] != ele[22][20];
    ele[18][18] != ele[22][21];
    ele[18][18] != ele[22][22];
    ele[18][18] != ele[22][23];
    ele[18][18] != ele[23][18];
    ele[18][18] != ele[23][19];
    ele[18][18] != ele[23][20];
    ele[18][18] != ele[23][21];
    ele[18][18] != ele[23][22];
    ele[18][18] != ele[23][23];
    ele[18][18] != ele[24][18];
    ele[18][18] != ele[25][18];
    ele[18][18] != ele[26][18];
    ele[18][18] != ele[27][18];
    ele[18][18] != ele[28][18];
    ele[18][18] != ele[29][18];
    ele[18][18] != ele[30][18];
    ele[18][18] != ele[31][18];
    ele[18][18] != ele[32][18];
    ele[18][18] != ele[33][18];
    ele[18][18] != ele[34][18];
    ele[18][18] != ele[35][18];
    ele[18][19] != ele[18][20];
    ele[18][19] != ele[18][21];
    ele[18][19] != ele[18][22];
    ele[18][19] != ele[18][23];
    ele[18][19] != ele[18][24];
    ele[18][19] != ele[18][25];
    ele[18][19] != ele[18][26];
    ele[18][19] != ele[18][27];
    ele[18][19] != ele[18][28];
    ele[18][19] != ele[18][29];
    ele[18][19] != ele[18][30];
    ele[18][19] != ele[18][31];
    ele[18][19] != ele[18][32];
    ele[18][19] != ele[18][33];
    ele[18][19] != ele[18][34];
    ele[18][19] != ele[18][35];
    ele[18][19] != ele[19][18];
    ele[18][19] != ele[19][19];
    ele[18][19] != ele[19][20];
    ele[18][19] != ele[19][21];
    ele[18][19] != ele[19][22];
    ele[18][19] != ele[19][23];
    ele[18][19] != ele[20][18];
    ele[18][19] != ele[20][19];
    ele[18][19] != ele[20][20];
    ele[18][19] != ele[20][21];
    ele[18][19] != ele[20][22];
    ele[18][19] != ele[20][23];
    ele[18][19] != ele[21][18];
    ele[18][19] != ele[21][19];
    ele[18][19] != ele[21][20];
    ele[18][19] != ele[21][21];
    ele[18][19] != ele[21][22];
    ele[18][19] != ele[21][23];
    ele[18][19] != ele[22][18];
    ele[18][19] != ele[22][19];
    ele[18][19] != ele[22][20];
    ele[18][19] != ele[22][21];
    ele[18][19] != ele[22][22];
    ele[18][19] != ele[22][23];
    ele[18][19] != ele[23][18];
    ele[18][19] != ele[23][19];
    ele[18][19] != ele[23][20];
    ele[18][19] != ele[23][21];
    ele[18][19] != ele[23][22];
    ele[18][19] != ele[23][23];
    ele[18][19] != ele[24][19];
    ele[18][19] != ele[25][19];
    ele[18][19] != ele[26][19];
    ele[18][19] != ele[27][19];
    ele[18][19] != ele[28][19];
    ele[18][19] != ele[29][19];
    ele[18][19] != ele[30][19];
    ele[18][19] != ele[31][19];
    ele[18][19] != ele[32][19];
    ele[18][19] != ele[33][19];
    ele[18][19] != ele[34][19];
    ele[18][19] != ele[35][19];
    ele[18][2] != ele[18][10];
    ele[18][2] != ele[18][11];
    ele[18][2] != ele[18][12];
    ele[18][2] != ele[18][13];
    ele[18][2] != ele[18][14];
    ele[18][2] != ele[18][15];
    ele[18][2] != ele[18][16];
    ele[18][2] != ele[18][17];
    ele[18][2] != ele[18][18];
    ele[18][2] != ele[18][19];
    ele[18][2] != ele[18][20];
    ele[18][2] != ele[18][21];
    ele[18][2] != ele[18][22];
    ele[18][2] != ele[18][23];
    ele[18][2] != ele[18][24];
    ele[18][2] != ele[18][25];
    ele[18][2] != ele[18][26];
    ele[18][2] != ele[18][27];
    ele[18][2] != ele[18][28];
    ele[18][2] != ele[18][29];
    ele[18][2] != ele[18][3];
    ele[18][2] != ele[18][30];
    ele[18][2] != ele[18][31];
    ele[18][2] != ele[18][32];
    ele[18][2] != ele[18][33];
    ele[18][2] != ele[18][34];
    ele[18][2] != ele[18][35];
    ele[18][2] != ele[18][4];
    ele[18][2] != ele[18][5];
    ele[18][2] != ele[18][6];
    ele[18][2] != ele[18][7];
    ele[18][2] != ele[18][8];
    ele[18][2] != ele[18][9];
    ele[18][2] != ele[19][0];
    ele[18][2] != ele[19][1];
    ele[18][2] != ele[19][2];
    ele[18][2] != ele[19][3];
    ele[18][2] != ele[19][4];
    ele[18][2] != ele[19][5];
    ele[18][2] != ele[20][0];
    ele[18][2] != ele[20][1];
    ele[18][2] != ele[20][2];
    ele[18][2] != ele[20][3];
    ele[18][2] != ele[20][4];
    ele[18][2] != ele[20][5];
    ele[18][2] != ele[21][0];
    ele[18][2] != ele[21][1];
    ele[18][2] != ele[21][2];
    ele[18][2] != ele[21][3];
    ele[18][2] != ele[21][4];
    ele[18][2] != ele[21][5];
    ele[18][2] != ele[22][0];
    ele[18][2] != ele[22][1];
    ele[18][2] != ele[22][2];
    ele[18][2] != ele[22][3];
    ele[18][2] != ele[22][4];
    ele[18][2] != ele[22][5];
    ele[18][2] != ele[23][0];
    ele[18][2] != ele[23][1];
    ele[18][2] != ele[23][2];
    ele[18][2] != ele[23][3];
    ele[18][2] != ele[23][4];
    ele[18][2] != ele[23][5];
    ele[18][2] != ele[24][2];
    ele[18][2] != ele[25][2];
    ele[18][2] != ele[26][2];
    ele[18][2] != ele[27][2];
    ele[18][2] != ele[28][2];
    ele[18][2] != ele[29][2];
    ele[18][2] != ele[30][2];
    ele[18][2] != ele[31][2];
    ele[18][2] != ele[32][2];
    ele[18][2] != ele[33][2];
    ele[18][2] != ele[34][2];
    ele[18][2] != ele[35][2];
    ele[18][20] != ele[18][21];
    ele[18][20] != ele[18][22];
    ele[18][20] != ele[18][23];
    ele[18][20] != ele[18][24];
    ele[18][20] != ele[18][25];
    ele[18][20] != ele[18][26];
    ele[18][20] != ele[18][27];
    ele[18][20] != ele[18][28];
    ele[18][20] != ele[18][29];
    ele[18][20] != ele[18][30];
    ele[18][20] != ele[18][31];
    ele[18][20] != ele[18][32];
    ele[18][20] != ele[18][33];
    ele[18][20] != ele[18][34];
    ele[18][20] != ele[18][35];
    ele[18][20] != ele[19][18];
    ele[18][20] != ele[19][19];
    ele[18][20] != ele[19][20];
    ele[18][20] != ele[19][21];
    ele[18][20] != ele[19][22];
    ele[18][20] != ele[19][23];
    ele[18][20] != ele[20][18];
    ele[18][20] != ele[20][19];
    ele[18][20] != ele[20][20];
    ele[18][20] != ele[20][21];
    ele[18][20] != ele[20][22];
    ele[18][20] != ele[20][23];
    ele[18][20] != ele[21][18];
    ele[18][20] != ele[21][19];
    ele[18][20] != ele[21][20];
    ele[18][20] != ele[21][21];
    ele[18][20] != ele[21][22];
    ele[18][20] != ele[21][23];
    ele[18][20] != ele[22][18];
    ele[18][20] != ele[22][19];
    ele[18][20] != ele[22][20];
    ele[18][20] != ele[22][21];
    ele[18][20] != ele[22][22];
    ele[18][20] != ele[22][23];
    ele[18][20] != ele[23][18];
    ele[18][20] != ele[23][19];
    ele[18][20] != ele[23][20];
    ele[18][20] != ele[23][21];
    ele[18][20] != ele[23][22];
    ele[18][20] != ele[23][23];
    ele[18][20] != ele[24][20];
    ele[18][20] != ele[25][20];
    ele[18][20] != ele[26][20];
    ele[18][20] != ele[27][20];
    ele[18][20] != ele[28][20];
    ele[18][20] != ele[29][20];
    ele[18][20] != ele[30][20];
    ele[18][20] != ele[31][20];
    ele[18][20] != ele[32][20];
    ele[18][20] != ele[33][20];
    ele[18][20] != ele[34][20];
    ele[18][20] != ele[35][20];
    ele[18][21] != ele[18][22];
    ele[18][21] != ele[18][23];
    ele[18][21] != ele[18][24];
    ele[18][21] != ele[18][25];
    ele[18][21] != ele[18][26];
    ele[18][21] != ele[18][27];
    ele[18][21] != ele[18][28];
    ele[18][21] != ele[18][29];
    ele[18][21] != ele[18][30];
    ele[18][21] != ele[18][31];
    ele[18][21] != ele[18][32];
    ele[18][21] != ele[18][33];
    ele[18][21] != ele[18][34];
    ele[18][21] != ele[18][35];
    ele[18][21] != ele[19][18];
    ele[18][21] != ele[19][19];
    ele[18][21] != ele[19][20];
    ele[18][21] != ele[19][21];
    ele[18][21] != ele[19][22];
    ele[18][21] != ele[19][23];
    ele[18][21] != ele[20][18];
    ele[18][21] != ele[20][19];
    ele[18][21] != ele[20][20];
    ele[18][21] != ele[20][21];
    ele[18][21] != ele[20][22];
    ele[18][21] != ele[20][23];
    ele[18][21] != ele[21][18];
    ele[18][21] != ele[21][19];
    ele[18][21] != ele[21][20];
    ele[18][21] != ele[21][21];
    ele[18][21] != ele[21][22];
    ele[18][21] != ele[21][23];
    ele[18][21] != ele[22][18];
    ele[18][21] != ele[22][19];
    ele[18][21] != ele[22][20];
    ele[18][21] != ele[22][21];
    ele[18][21] != ele[22][22];
    ele[18][21] != ele[22][23];
    ele[18][21] != ele[23][18];
    ele[18][21] != ele[23][19];
    ele[18][21] != ele[23][20];
    ele[18][21] != ele[23][21];
    ele[18][21] != ele[23][22];
    ele[18][21] != ele[23][23];
    ele[18][21] != ele[24][21];
    ele[18][21] != ele[25][21];
    ele[18][21] != ele[26][21];
    ele[18][21] != ele[27][21];
    ele[18][21] != ele[28][21];
    ele[18][21] != ele[29][21];
    ele[18][21] != ele[30][21];
    ele[18][21] != ele[31][21];
    ele[18][21] != ele[32][21];
    ele[18][21] != ele[33][21];
    ele[18][21] != ele[34][21];
    ele[18][21] != ele[35][21];
    ele[18][22] != ele[18][23];
    ele[18][22] != ele[18][24];
    ele[18][22] != ele[18][25];
    ele[18][22] != ele[18][26];
    ele[18][22] != ele[18][27];
    ele[18][22] != ele[18][28];
    ele[18][22] != ele[18][29];
    ele[18][22] != ele[18][30];
    ele[18][22] != ele[18][31];
    ele[18][22] != ele[18][32];
    ele[18][22] != ele[18][33];
    ele[18][22] != ele[18][34];
    ele[18][22] != ele[18][35];
    ele[18][22] != ele[19][18];
    ele[18][22] != ele[19][19];
    ele[18][22] != ele[19][20];
    ele[18][22] != ele[19][21];
    ele[18][22] != ele[19][22];
    ele[18][22] != ele[19][23];
    ele[18][22] != ele[20][18];
    ele[18][22] != ele[20][19];
    ele[18][22] != ele[20][20];
    ele[18][22] != ele[20][21];
    ele[18][22] != ele[20][22];
    ele[18][22] != ele[20][23];
    ele[18][22] != ele[21][18];
    ele[18][22] != ele[21][19];
    ele[18][22] != ele[21][20];
    ele[18][22] != ele[21][21];
    ele[18][22] != ele[21][22];
    ele[18][22] != ele[21][23];
    ele[18][22] != ele[22][18];
    ele[18][22] != ele[22][19];
    ele[18][22] != ele[22][20];
    ele[18][22] != ele[22][21];
    ele[18][22] != ele[22][22];
    ele[18][22] != ele[22][23];
    ele[18][22] != ele[23][18];
    ele[18][22] != ele[23][19];
    ele[18][22] != ele[23][20];
    ele[18][22] != ele[23][21];
    ele[18][22] != ele[23][22];
    ele[18][22] != ele[23][23];
    ele[18][22] != ele[24][22];
    ele[18][22] != ele[25][22];
    ele[18][22] != ele[26][22];
    ele[18][22] != ele[27][22];
    ele[18][22] != ele[28][22];
    ele[18][22] != ele[29][22];
    ele[18][22] != ele[30][22];
    ele[18][22] != ele[31][22];
    ele[18][22] != ele[32][22];
    ele[18][22] != ele[33][22];
    ele[18][22] != ele[34][22];
    ele[18][22] != ele[35][22];
    ele[18][23] != ele[18][24];
    ele[18][23] != ele[18][25];
    ele[18][23] != ele[18][26];
    ele[18][23] != ele[18][27];
    ele[18][23] != ele[18][28];
    ele[18][23] != ele[18][29];
    ele[18][23] != ele[18][30];
    ele[18][23] != ele[18][31];
    ele[18][23] != ele[18][32];
    ele[18][23] != ele[18][33];
    ele[18][23] != ele[18][34];
    ele[18][23] != ele[18][35];
    ele[18][23] != ele[19][18];
    ele[18][23] != ele[19][19];
    ele[18][23] != ele[19][20];
    ele[18][23] != ele[19][21];
    ele[18][23] != ele[19][22];
    ele[18][23] != ele[19][23];
    ele[18][23] != ele[20][18];
    ele[18][23] != ele[20][19];
    ele[18][23] != ele[20][20];
    ele[18][23] != ele[20][21];
    ele[18][23] != ele[20][22];
    ele[18][23] != ele[20][23];
    ele[18][23] != ele[21][18];
    ele[18][23] != ele[21][19];
    ele[18][23] != ele[21][20];
    ele[18][23] != ele[21][21];
    ele[18][23] != ele[21][22];
    ele[18][23] != ele[21][23];
    ele[18][23] != ele[22][18];
    ele[18][23] != ele[22][19];
    ele[18][23] != ele[22][20];
    ele[18][23] != ele[22][21];
    ele[18][23] != ele[22][22];
    ele[18][23] != ele[22][23];
    ele[18][23] != ele[23][18];
    ele[18][23] != ele[23][19];
    ele[18][23] != ele[23][20];
    ele[18][23] != ele[23][21];
    ele[18][23] != ele[23][22];
    ele[18][23] != ele[23][23];
    ele[18][23] != ele[24][23];
    ele[18][23] != ele[25][23];
    ele[18][23] != ele[26][23];
    ele[18][23] != ele[27][23];
    ele[18][23] != ele[28][23];
    ele[18][23] != ele[29][23];
    ele[18][23] != ele[30][23];
    ele[18][23] != ele[31][23];
    ele[18][23] != ele[32][23];
    ele[18][23] != ele[33][23];
    ele[18][23] != ele[34][23];
    ele[18][23] != ele[35][23];
    ele[18][24] != ele[18][25];
    ele[18][24] != ele[18][26];
    ele[18][24] != ele[18][27];
    ele[18][24] != ele[18][28];
    ele[18][24] != ele[18][29];
    ele[18][24] != ele[18][30];
    ele[18][24] != ele[18][31];
    ele[18][24] != ele[18][32];
    ele[18][24] != ele[18][33];
    ele[18][24] != ele[18][34];
    ele[18][24] != ele[18][35];
    ele[18][24] != ele[19][24];
    ele[18][24] != ele[19][25];
    ele[18][24] != ele[19][26];
    ele[18][24] != ele[19][27];
    ele[18][24] != ele[19][28];
    ele[18][24] != ele[19][29];
    ele[18][24] != ele[20][24];
    ele[18][24] != ele[20][25];
    ele[18][24] != ele[20][26];
    ele[18][24] != ele[20][27];
    ele[18][24] != ele[20][28];
    ele[18][24] != ele[20][29];
    ele[18][24] != ele[21][24];
    ele[18][24] != ele[21][25];
    ele[18][24] != ele[21][26];
    ele[18][24] != ele[21][27];
    ele[18][24] != ele[21][28];
    ele[18][24] != ele[21][29];
    ele[18][24] != ele[22][24];
    ele[18][24] != ele[22][25];
    ele[18][24] != ele[22][26];
    ele[18][24] != ele[22][27];
    ele[18][24] != ele[22][28];
    ele[18][24] != ele[22][29];
    ele[18][24] != ele[23][24];
    ele[18][24] != ele[23][25];
    ele[18][24] != ele[23][26];
    ele[18][24] != ele[23][27];
    ele[18][24] != ele[23][28];
    ele[18][24] != ele[23][29];
    ele[18][24] != ele[24][24];
    ele[18][24] != ele[25][24];
    ele[18][24] != ele[26][24];
    ele[18][24] != ele[27][24];
    ele[18][24] != ele[28][24];
    ele[18][24] != ele[29][24];
    ele[18][24] != ele[30][24];
    ele[18][24] != ele[31][24];
    ele[18][24] != ele[32][24];
    ele[18][24] != ele[33][24];
    ele[18][24] != ele[34][24];
    ele[18][24] != ele[35][24];
    ele[18][25] != ele[18][26];
    ele[18][25] != ele[18][27];
    ele[18][25] != ele[18][28];
    ele[18][25] != ele[18][29];
    ele[18][25] != ele[18][30];
    ele[18][25] != ele[18][31];
    ele[18][25] != ele[18][32];
    ele[18][25] != ele[18][33];
    ele[18][25] != ele[18][34];
    ele[18][25] != ele[18][35];
    ele[18][25] != ele[19][24];
    ele[18][25] != ele[19][25];
    ele[18][25] != ele[19][26];
    ele[18][25] != ele[19][27];
    ele[18][25] != ele[19][28];
    ele[18][25] != ele[19][29];
    ele[18][25] != ele[20][24];
    ele[18][25] != ele[20][25];
    ele[18][25] != ele[20][26];
    ele[18][25] != ele[20][27];
    ele[18][25] != ele[20][28];
    ele[18][25] != ele[20][29];
    ele[18][25] != ele[21][24];
    ele[18][25] != ele[21][25];
    ele[18][25] != ele[21][26];
    ele[18][25] != ele[21][27];
    ele[18][25] != ele[21][28];
    ele[18][25] != ele[21][29];
    ele[18][25] != ele[22][24];
    ele[18][25] != ele[22][25];
    ele[18][25] != ele[22][26];
    ele[18][25] != ele[22][27];
    ele[18][25] != ele[22][28];
    ele[18][25] != ele[22][29];
    ele[18][25] != ele[23][24];
    ele[18][25] != ele[23][25];
    ele[18][25] != ele[23][26];
    ele[18][25] != ele[23][27];
    ele[18][25] != ele[23][28];
    ele[18][25] != ele[23][29];
    ele[18][25] != ele[24][25];
    ele[18][25] != ele[25][25];
    ele[18][25] != ele[26][25];
    ele[18][25] != ele[27][25];
    ele[18][25] != ele[28][25];
    ele[18][25] != ele[29][25];
    ele[18][25] != ele[30][25];
    ele[18][25] != ele[31][25];
    ele[18][25] != ele[32][25];
    ele[18][25] != ele[33][25];
    ele[18][25] != ele[34][25];
    ele[18][25] != ele[35][25];
    ele[18][26] != ele[18][27];
    ele[18][26] != ele[18][28];
    ele[18][26] != ele[18][29];
    ele[18][26] != ele[18][30];
    ele[18][26] != ele[18][31];
    ele[18][26] != ele[18][32];
    ele[18][26] != ele[18][33];
    ele[18][26] != ele[18][34];
    ele[18][26] != ele[18][35];
    ele[18][26] != ele[19][24];
    ele[18][26] != ele[19][25];
    ele[18][26] != ele[19][26];
    ele[18][26] != ele[19][27];
    ele[18][26] != ele[19][28];
    ele[18][26] != ele[19][29];
    ele[18][26] != ele[20][24];
    ele[18][26] != ele[20][25];
    ele[18][26] != ele[20][26];
    ele[18][26] != ele[20][27];
    ele[18][26] != ele[20][28];
    ele[18][26] != ele[20][29];
    ele[18][26] != ele[21][24];
    ele[18][26] != ele[21][25];
    ele[18][26] != ele[21][26];
    ele[18][26] != ele[21][27];
    ele[18][26] != ele[21][28];
    ele[18][26] != ele[21][29];
    ele[18][26] != ele[22][24];
    ele[18][26] != ele[22][25];
    ele[18][26] != ele[22][26];
    ele[18][26] != ele[22][27];
    ele[18][26] != ele[22][28];
    ele[18][26] != ele[22][29];
    ele[18][26] != ele[23][24];
    ele[18][26] != ele[23][25];
    ele[18][26] != ele[23][26];
    ele[18][26] != ele[23][27];
    ele[18][26] != ele[23][28];
    ele[18][26] != ele[23][29];
    ele[18][26] != ele[24][26];
    ele[18][26] != ele[25][26];
    ele[18][26] != ele[26][26];
    ele[18][26] != ele[27][26];
    ele[18][26] != ele[28][26];
    ele[18][26] != ele[29][26];
    ele[18][26] != ele[30][26];
    ele[18][26] != ele[31][26];
    ele[18][26] != ele[32][26];
    ele[18][26] != ele[33][26];
    ele[18][26] != ele[34][26];
    ele[18][26] != ele[35][26];
    ele[18][27] != ele[18][28];
    ele[18][27] != ele[18][29];
    ele[18][27] != ele[18][30];
    ele[18][27] != ele[18][31];
    ele[18][27] != ele[18][32];
    ele[18][27] != ele[18][33];
    ele[18][27] != ele[18][34];
    ele[18][27] != ele[18][35];
    ele[18][27] != ele[19][24];
    ele[18][27] != ele[19][25];
    ele[18][27] != ele[19][26];
    ele[18][27] != ele[19][27];
    ele[18][27] != ele[19][28];
    ele[18][27] != ele[19][29];
    ele[18][27] != ele[20][24];
    ele[18][27] != ele[20][25];
    ele[18][27] != ele[20][26];
    ele[18][27] != ele[20][27];
    ele[18][27] != ele[20][28];
    ele[18][27] != ele[20][29];
    ele[18][27] != ele[21][24];
    ele[18][27] != ele[21][25];
    ele[18][27] != ele[21][26];
    ele[18][27] != ele[21][27];
    ele[18][27] != ele[21][28];
    ele[18][27] != ele[21][29];
    ele[18][27] != ele[22][24];
    ele[18][27] != ele[22][25];
    ele[18][27] != ele[22][26];
    ele[18][27] != ele[22][27];
    ele[18][27] != ele[22][28];
    ele[18][27] != ele[22][29];
    ele[18][27] != ele[23][24];
    ele[18][27] != ele[23][25];
    ele[18][27] != ele[23][26];
    ele[18][27] != ele[23][27];
    ele[18][27] != ele[23][28];
    ele[18][27] != ele[23][29];
    ele[18][27] != ele[24][27];
    ele[18][27] != ele[25][27];
    ele[18][27] != ele[26][27];
    ele[18][27] != ele[27][27];
    ele[18][27] != ele[28][27];
    ele[18][27] != ele[29][27];
    ele[18][27] != ele[30][27];
    ele[18][27] != ele[31][27];
    ele[18][27] != ele[32][27];
    ele[18][27] != ele[33][27];
    ele[18][27] != ele[34][27];
    ele[18][27] != ele[35][27];
    ele[18][28] != ele[18][29];
    ele[18][28] != ele[18][30];
    ele[18][28] != ele[18][31];
    ele[18][28] != ele[18][32];
    ele[18][28] != ele[18][33];
    ele[18][28] != ele[18][34];
    ele[18][28] != ele[18][35];
    ele[18][28] != ele[19][24];
    ele[18][28] != ele[19][25];
    ele[18][28] != ele[19][26];
    ele[18][28] != ele[19][27];
    ele[18][28] != ele[19][28];
    ele[18][28] != ele[19][29];
    ele[18][28] != ele[20][24];
    ele[18][28] != ele[20][25];
    ele[18][28] != ele[20][26];
    ele[18][28] != ele[20][27];
    ele[18][28] != ele[20][28];
    ele[18][28] != ele[20][29];
    ele[18][28] != ele[21][24];
    ele[18][28] != ele[21][25];
    ele[18][28] != ele[21][26];
    ele[18][28] != ele[21][27];
    ele[18][28] != ele[21][28];
    ele[18][28] != ele[21][29];
    ele[18][28] != ele[22][24];
    ele[18][28] != ele[22][25];
    ele[18][28] != ele[22][26];
    ele[18][28] != ele[22][27];
    ele[18][28] != ele[22][28];
    ele[18][28] != ele[22][29];
    ele[18][28] != ele[23][24];
    ele[18][28] != ele[23][25];
    ele[18][28] != ele[23][26];
    ele[18][28] != ele[23][27];
    ele[18][28] != ele[23][28];
    ele[18][28] != ele[23][29];
    ele[18][28] != ele[24][28];
    ele[18][28] != ele[25][28];
    ele[18][28] != ele[26][28];
    ele[18][28] != ele[27][28];
    ele[18][28] != ele[28][28];
    ele[18][28] != ele[29][28];
    ele[18][28] != ele[30][28];
    ele[18][28] != ele[31][28];
    ele[18][28] != ele[32][28];
    ele[18][28] != ele[33][28];
    ele[18][28] != ele[34][28];
    ele[18][28] != ele[35][28];
    ele[18][29] != ele[18][30];
    ele[18][29] != ele[18][31];
    ele[18][29] != ele[18][32];
    ele[18][29] != ele[18][33];
    ele[18][29] != ele[18][34];
    ele[18][29] != ele[18][35];
    ele[18][29] != ele[19][24];
    ele[18][29] != ele[19][25];
    ele[18][29] != ele[19][26];
    ele[18][29] != ele[19][27];
    ele[18][29] != ele[19][28];
    ele[18][29] != ele[19][29];
    ele[18][29] != ele[20][24];
    ele[18][29] != ele[20][25];
    ele[18][29] != ele[20][26];
    ele[18][29] != ele[20][27];
    ele[18][29] != ele[20][28];
    ele[18][29] != ele[20][29];
    ele[18][29] != ele[21][24];
    ele[18][29] != ele[21][25];
    ele[18][29] != ele[21][26];
    ele[18][29] != ele[21][27];
    ele[18][29] != ele[21][28];
    ele[18][29] != ele[21][29];
    ele[18][29] != ele[22][24];
    ele[18][29] != ele[22][25];
    ele[18][29] != ele[22][26];
    ele[18][29] != ele[22][27];
    ele[18][29] != ele[22][28];
    ele[18][29] != ele[22][29];
    ele[18][29] != ele[23][24];
    ele[18][29] != ele[23][25];
    ele[18][29] != ele[23][26];
    ele[18][29] != ele[23][27];
    ele[18][29] != ele[23][28];
    ele[18][29] != ele[23][29];
    ele[18][29] != ele[24][29];
    ele[18][29] != ele[25][29];
    ele[18][29] != ele[26][29];
    ele[18][29] != ele[27][29];
    ele[18][29] != ele[28][29];
    ele[18][29] != ele[29][29];
    ele[18][29] != ele[30][29];
    ele[18][29] != ele[31][29];
    ele[18][29] != ele[32][29];
    ele[18][29] != ele[33][29];
    ele[18][29] != ele[34][29];
    ele[18][29] != ele[35][29];
    ele[18][3] != ele[18][10];
    ele[18][3] != ele[18][11];
    ele[18][3] != ele[18][12];
    ele[18][3] != ele[18][13];
    ele[18][3] != ele[18][14];
    ele[18][3] != ele[18][15];
    ele[18][3] != ele[18][16];
    ele[18][3] != ele[18][17];
    ele[18][3] != ele[18][18];
    ele[18][3] != ele[18][19];
    ele[18][3] != ele[18][20];
    ele[18][3] != ele[18][21];
    ele[18][3] != ele[18][22];
    ele[18][3] != ele[18][23];
    ele[18][3] != ele[18][24];
    ele[18][3] != ele[18][25];
    ele[18][3] != ele[18][26];
    ele[18][3] != ele[18][27];
    ele[18][3] != ele[18][28];
    ele[18][3] != ele[18][29];
    ele[18][3] != ele[18][30];
    ele[18][3] != ele[18][31];
    ele[18][3] != ele[18][32];
    ele[18][3] != ele[18][33];
    ele[18][3] != ele[18][34];
    ele[18][3] != ele[18][35];
    ele[18][3] != ele[18][4];
    ele[18][3] != ele[18][5];
    ele[18][3] != ele[18][6];
    ele[18][3] != ele[18][7];
    ele[18][3] != ele[18][8];
    ele[18][3] != ele[18][9];
    ele[18][3] != ele[19][0];
    ele[18][3] != ele[19][1];
    ele[18][3] != ele[19][2];
    ele[18][3] != ele[19][3];
    ele[18][3] != ele[19][4];
    ele[18][3] != ele[19][5];
    ele[18][3] != ele[20][0];
    ele[18][3] != ele[20][1];
    ele[18][3] != ele[20][2];
    ele[18][3] != ele[20][3];
    ele[18][3] != ele[20][4];
    ele[18][3] != ele[20][5];
    ele[18][3] != ele[21][0];
    ele[18][3] != ele[21][1];
    ele[18][3] != ele[21][2];
    ele[18][3] != ele[21][3];
    ele[18][3] != ele[21][4];
    ele[18][3] != ele[21][5];
    ele[18][3] != ele[22][0];
    ele[18][3] != ele[22][1];
    ele[18][3] != ele[22][2];
    ele[18][3] != ele[22][3];
    ele[18][3] != ele[22][4];
    ele[18][3] != ele[22][5];
    ele[18][3] != ele[23][0];
    ele[18][3] != ele[23][1];
    ele[18][3] != ele[23][2];
    ele[18][3] != ele[23][3];
    ele[18][3] != ele[23][4];
    ele[18][3] != ele[23][5];
    ele[18][3] != ele[24][3];
    ele[18][3] != ele[25][3];
    ele[18][3] != ele[26][3];
    ele[18][3] != ele[27][3];
    ele[18][3] != ele[28][3];
    ele[18][3] != ele[29][3];
    ele[18][3] != ele[30][3];
    ele[18][3] != ele[31][3];
    ele[18][3] != ele[32][3];
    ele[18][3] != ele[33][3];
    ele[18][3] != ele[34][3];
    ele[18][3] != ele[35][3];
    ele[18][30] != ele[18][31];
    ele[18][30] != ele[18][32];
    ele[18][30] != ele[18][33];
    ele[18][30] != ele[18][34];
    ele[18][30] != ele[18][35];
    ele[18][30] != ele[19][30];
    ele[18][30] != ele[19][31];
    ele[18][30] != ele[19][32];
    ele[18][30] != ele[19][33];
    ele[18][30] != ele[19][34];
    ele[18][30] != ele[19][35];
    ele[18][30] != ele[20][30];
    ele[18][30] != ele[20][31];
    ele[18][30] != ele[20][32];
    ele[18][30] != ele[20][33];
    ele[18][30] != ele[20][34];
    ele[18][30] != ele[20][35];
    ele[18][30] != ele[21][30];
    ele[18][30] != ele[21][31];
    ele[18][30] != ele[21][32];
    ele[18][30] != ele[21][33];
    ele[18][30] != ele[21][34];
    ele[18][30] != ele[21][35];
    ele[18][30] != ele[22][30];
    ele[18][30] != ele[22][31];
    ele[18][30] != ele[22][32];
    ele[18][30] != ele[22][33];
    ele[18][30] != ele[22][34];
    ele[18][30] != ele[22][35];
    ele[18][30] != ele[23][30];
    ele[18][30] != ele[23][31];
    ele[18][30] != ele[23][32];
    ele[18][30] != ele[23][33];
    ele[18][30] != ele[23][34];
    ele[18][30] != ele[23][35];
    ele[18][30] != ele[24][30];
    ele[18][30] != ele[25][30];
    ele[18][30] != ele[26][30];
    ele[18][30] != ele[27][30];
    ele[18][30] != ele[28][30];
    ele[18][30] != ele[29][30];
    ele[18][30] != ele[30][30];
    ele[18][30] != ele[31][30];
    ele[18][30] != ele[32][30];
    ele[18][30] != ele[33][30];
    ele[18][30] != ele[34][30];
    ele[18][30] != ele[35][30];
    ele[18][31] != ele[18][32];
    ele[18][31] != ele[18][33];
    ele[18][31] != ele[18][34];
    ele[18][31] != ele[18][35];
    ele[18][31] != ele[19][30];
    ele[18][31] != ele[19][31];
    ele[18][31] != ele[19][32];
    ele[18][31] != ele[19][33];
    ele[18][31] != ele[19][34];
    ele[18][31] != ele[19][35];
    ele[18][31] != ele[20][30];
    ele[18][31] != ele[20][31];
    ele[18][31] != ele[20][32];
    ele[18][31] != ele[20][33];
    ele[18][31] != ele[20][34];
    ele[18][31] != ele[20][35];
    ele[18][31] != ele[21][30];
    ele[18][31] != ele[21][31];
    ele[18][31] != ele[21][32];
    ele[18][31] != ele[21][33];
    ele[18][31] != ele[21][34];
    ele[18][31] != ele[21][35];
    ele[18][31] != ele[22][30];
    ele[18][31] != ele[22][31];
    ele[18][31] != ele[22][32];
    ele[18][31] != ele[22][33];
    ele[18][31] != ele[22][34];
    ele[18][31] != ele[22][35];
    ele[18][31] != ele[23][30];
    ele[18][31] != ele[23][31];
    ele[18][31] != ele[23][32];
    ele[18][31] != ele[23][33];
    ele[18][31] != ele[23][34];
    ele[18][31] != ele[23][35];
    ele[18][31] != ele[24][31];
    ele[18][31] != ele[25][31];
    ele[18][31] != ele[26][31];
    ele[18][31] != ele[27][31];
    ele[18][31] != ele[28][31];
    ele[18][31] != ele[29][31];
    ele[18][31] != ele[30][31];
    ele[18][31] != ele[31][31];
    ele[18][31] != ele[32][31];
    ele[18][31] != ele[33][31];
    ele[18][31] != ele[34][31];
    ele[18][31] != ele[35][31];
    ele[18][32] != ele[18][33];
    ele[18][32] != ele[18][34];
    ele[18][32] != ele[18][35];
    ele[18][32] != ele[19][30];
    ele[18][32] != ele[19][31];
    ele[18][32] != ele[19][32];
    ele[18][32] != ele[19][33];
    ele[18][32] != ele[19][34];
    ele[18][32] != ele[19][35];
    ele[18][32] != ele[20][30];
    ele[18][32] != ele[20][31];
    ele[18][32] != ele[20][32];
    ele[18][32] != ele[20][33];
    ele[18][32] != ele[20][34];
    ele[18][32] != ele[20][35];
    ele[18][32] != ele[21][30];
    ele[18][32] != ele[21][31];
    ele[18][32] != ele[21][32];
    ele[18][32] != ele[21][33];
    ele[18][32] != ele[21][34];
    ele[18][32] != ele[21][35];
    ele[18][32] != ele[22][30];
    ele[18][32] != ele[22][31];
    ele[18][32] != ele[22][32];
    ele[18][32] != ele[22][33];
    ele[18][32] != ele[22][34];
    ele[18][32] != ele[22][35];
    ele[18][32] != ele[23][30];
    ele[18][32] != ele[23][31];
    ele[18][32] != ele[23][32];
    ele[18][32] != ele[23][33];
    ele[18][32] != ele[23][34];
    ele[18][32] != ele[23][35];
    ele[18][32] != ele[24][32];
    ele[18][32] != ele[25][32];
    ele[18][32] != ele[26][32];
    ele[18][32] != ele[27][32];
    ele[18][32] != ele[28][32];
    ele[18][32] != ele[29][32];
    ele[18][32] != ele[30][32];
    ele[18][32] != ele[31][32];
    ele[18][32] != ele[32][32];
    ele[18][32] != ele[33][32];
    ele[18][32] != ele[34][32];
    ele[18][32] != ele[35][32];
    ele[18][33] != ele[18][34];
    ele[18][33] != ele[18][35];
    ele[18][33] != ele[19][30];
    ele[18][33] != ele[19][31];
    ele[18][33] != ele[19][32];
    ele[18][33] != ele[19][33];
    ele[18][33] != ele[19][34];
    ele[18][33] != ele[19][35];
    ele[18][33] != ele[20][30];
    ele[18][33] != ele[20][31];
    ele[18][33] != ele[20][32];
    ele[18][33] != ele[20][33];
    ele[18][33] != ele[20][34];
    ele[18][33] != ele[20][35];
    ele[18][33] != ele[21][30];
    ele[18][33] != ele[21][31];
    ele[18][33] != ele[21][32];
    ele[18][33] != ele[21][33];
    ele[18][33] != ele[21][34];
    ele[18][33] != ele[21][35];
    ele[18][33] != ele[22][30];
    ele[18][33] != ele[22][31];
    ele[18][33] != ele[22][32];
    ele[18][33] != ele[22][33];
    ele[18][33] != ele[22][34];
    ele[18][33] != ele[22][35];
    ele[18][33] != ele[23][30];
    ele[18][33] != ele[23][31];
    ele[18][33] != ele[23][32];
    ele[18][33] != ele[23][33];
    ele[18][33] != ele[23][34];
    ele[18][33] != ele[23][35];
    ele[18][33] != ele[24][33];
    ele[18][33] != ele[25][33];
    ele[18][33] != ele[26][33];
    ele[18][33] != ele[27][33];
    ele[18][33] != ele[28][33];
    ele[18][33] != ele[29][33];
    ele[18][33] != ele[30][33];
    ele[18][33] != ele[31][33];
    ele[18][33] != ele[32][33];
    ele[18][33] != ele[33][33];
    ele[18][33] != ele[34][33];
    ele[18][33] != ele[35][33];
    ele[18][34] != ele[18][35];
    ele[18][34] != ele[19][30];
    ele[18][34] != ele[19][31];
    ele[18][34] != ele[19][32];
    ele[18][34] != ele[19][33];
    ele[18][34] != ele[19][34];
    ele[18][34] != ele[19][35];
    ele[18][34] != ele[20][30];
    ele[18][34] != ele[20][31];
    ele[18][34] != ele[20][32];
    ele[18][34] != ele[20][33];
    ele[18][34] != ele[20][34];
    ele[18][34] != ele[20][35];
    ele[18][34] != ele[21][30];
    ele[18][34] != ele[21][31];
    ele[18][34] != ele[21][32];
    ele[18][34] != ele[21][33];
    ele[18][34] != ele[21][34];
    ele[18][34] != ele[21][35];
    ele[18][34] != ele[22][30];
    ele[18][34] != ele[22][31];
    ele[18][34] != ele[22][32];
    ele[18][34] != ele[22][33];
    ele[18][34] != ele[22][34];
    ele[18][34] != ele[22][35];
    ele[18][34] != ele[23][30];
    ele[18][34] != ele[23][31];
    ele[18][34] != ele[23][32];
    ele[18][34] != ele[23][33];
    ele[18][34] != ele[23][34];
    ele[18][34] != ele[23][35];
    ele[18][34] != ele[24][34];
    ele[18][34] != ele[25][34];
    ele[18][34] != ele[26][34];
    ele[18][34] != ele[27][34];
    ele[18][34] != ele[28][34];
    ele[18][34] != ele[29][34];
    ele[18][34] != ele[30][34];
    ele[18][34] != ele[31][34];
    ele[18][34] != ele[32][34];
    ele[18][34] != ele[33][34];
    ele[18][34] != ele[34][34];
    ele[18][34] != ele[35][34];
    ele[18][35] != ele[19][30];
    ele[18][35] != ele[19][31];
    ele[18][35] != ele[19][32];
    ele[18][35] != ele[19][33];
    ele[18][35] != ele[19][34];
    ele[18][35] != ele[19][35];
    ele[18][35] != ele[20][30];
    ele[18][35] != ele[20][31];
    ele[18][35] != ele[20][32];
    ele[18][35] != ele[20][33];
    ele[18][35] != ele[20][34];
    ele[18][35] != ele[20][35];
    ele[18][35] != ele[21][30];
    ele[18][35] != ele[21][31];
    ele[18][35] != ele[21][32];
    ele[18][35] != ele[21][33];
    ele[18][35] != ele[21][34];
    ele[18][35] != ele[21][35];
    ele[18][35] != ele[22][30];
    ele[18][35] != ele[22][31];
    ele[18][35] != ele[22][32];
    ele[18][35] != ele[22][33];
    ele[18][35] != ele[22][34];
    ele[18][35] != ele[22][35];
    ele[18][35] != ele[23][30];
    ele[18][35] != ele[23][31];
    ele[18][35] != ele[23][32];
    ele[18][35] != ele[23][33];
    ele[18][35] != ele[23][34];
    ele[18][35] != ele[23][35];
    ele[18][35] != ele[24][35];
    ele[18][35] != ele[25][35];
    ele[18][35] != ele[26][35];
    ele[18][35] != ele[27][35];
    ele[18][35] != ele[28][35];
    ele[18][35] != ele[29][35];
    ele[18][35] != ele[30][35];
    ele[18][35] != ele[31][35];
    ele[18][35] != ele[32][35];
    ele[18][35] != ele[33][35];
    ele[18][35] != ele[34][35];
    ele[18][35] != ele[35][35];
    ele[18][4] != ele[18][10];
    ele[18][4] != ele[18][11];
    ele[18][4] != ele[18][12];
    ele[18][4] != ele[18][13];
    ele[18][4] != ele[18][14];
    ele[18][4] != ele[18][15];
    ele[18][4] != ele[18][16];
    ele[18][4] != ele[18][17];
    ele[18][4] != ele[18][18];
    ele[18][4] != ele[18][19];
    ele[18][4] != ele[18][20];
    ele[18][4] != ele[18][21];
    ele[18][4] != ele[18][22];
    ele[18][4] != ele[18][23];
    ele[18][4] != ele[18][24];
    ele[18][4] != ele[18][25];
    ele[18][4] != ele[18][26];
    ele[18][4] != ele[18][27];
    ele[18][4] != ele[18][28];
    ele[18][4] != ele[18][29];
    ele[18][4] != ele[18][30];
    ele[18][4] != ele[18][31];
    ele[18][4] != ele[18][32];
    ele[18][4] != ele[18][33];
    ele[18][4] != ele[18][34];
    ele[18][4] != ele[18][35];
    ele[18][4] != ele[18][5];
    ele[18][4] != ele[18][6];
    ele[18][4] != ele[18][7];
    ele[18][4] != ele[18][8];
    ele[18][4] != ele[18][9];
    ele[18][4] != ele[19][0];
    ele[18][4] != ele[19][1];
    ele[18][4] != ele[19][2];
    ele[18][4] != ele[19][3];
    ele[18][4] != ele[19][4];
    ele[18][4] != ele[19][5];
    ele[18][4] != ele[20][0];
    ele[18][4] != ele[20][1];
    ele[18][4] != ele[20][2];
    ele[18][4] != ele[20][3];
    ele[18][4] != ele[20][4];
    ele[18][4] != ele[20][5];
    ele[18][4] != ele[21][0];
    ele[18][4] != ele[21][1];
    ele[18][4] != ele[21][2];
    ele[18][4] != ele[21][3];
    ele[18][4] != ele[21][4];
    ele[18][4] != ele[21][5];
    ele[18][4] != ele[22][0];
    ele[18][4] != ele[22][1];
    ele[18][4] != ele[22][2];
    ele[18][4] != ele[22][3];
    ele[18][4] != ele[22][4];
    ele[18][4] != ele[22][5];
    ele[18][4] != ele[23][0];
    ele[18][4] != ele[23][1];
    ele[18][4] != ele[23][2];
    ele[18][4] != ele[23][3];
    ele[18][4] != ele[23][4];
    ele[18][4] != ele[23][5];
    ele[18][4] != ele[24][4];
    ele[18][4] != ele[25][4];
    ele[18][4] != ele[26][4];
    ele[18][4] != ele[27][4];
    ele[18][4] != ele[28][4];
    ele[18][4] != ele[29][4];
    ele[18][4] != ele[30][4];
    ele[18][4] != ele[31][4];
    ele[18][4] != ele[32][4];
    ele[18][4] != ele[33][4];
    ele[18][4] != ele[34][4];
    ele[18][4] != ele[35][4];
    ele[18][5] != ele[18][10];
    ele[18][5] != ele[18][11];
    ele[18][5] != ele[18][12];
    ele[18][5] != ele[18][13];
    ele[18][5] != ele[18][14];
    ele[18][5] != ele[18][15];
    ele[18][5] != ele[18][16];
    ele[18][5] != ele[18][17];
    ele[18][5] != ele[18][18];
    ele[18][5] != ele[18][19];
    ele[18][5] != ele[18][20];
    ele[18][5] != ele[18][21];
    ele[18][5] != ele[18][22];
    ele[18][5] != ele[18][23];
    ele[18][5] != ele[18][24];
    ele[18][5] != ele[18][25];
    ele[18][5] != ele[18][26];
    ele[18][5] != ele[18][27];
    ele[18][5] != ele[18][28];
    ele[18][5] != ele[18][29];
    ele[18][5] != ele[18][30];
    ele[18][5] != ele[18][31];
    ele[18][5] != ele[18][32];
    ele[18][5] != ele[18][33];
    ele[18][5] != ele[18][34];
    ele[18][5] != ele[18][35];
    ele[18][5] != ele[18][6];
    ele[18][5] != ele[18][7];
    ele[18][5] != ele[18][8];
    ele[18][5] != ele[18][9];
    ele[18][5] != ele[19][0];
    ele[18][5] != ele[19][1];
    ele[18][5] != ele[19][2];
    ele[18][5] != ele[19][3];
    ele[18][5] != ele[19][4];
    ele[18][5] != ele[19][5];
    ele[18][5] != ele[20][0];
    ele[18][5] != ele[20][1];
    ele[18][5] != ele[20][2];
    ele[18][5] != ele[20][3];
    ele[18][5] != ele[20][4];
    ele[18][5] != ele[20][5];
    ele[18][5] != ele[21][0];
    ele[18][5] != ele[21][1];
    ele[18][5] != ele[21][2];
    ele[18][5] != ele[21][3];
    ele[18][5] != ele[21][4];
    ele[18][5] != ele[21][5];
    ele[18][5] != ele[22][0];
    ele[18][5] != ele[22][1];
    ele[18][5] != ele[22][2];
    ele[18][5] != ele[22][3];
    ele[18][5] != ele[22][4];
    ele[18][5] != ele[22][5];
    ele[18][5] != ele[23][0];
    ele[18][5] != ele[23][1];
    ele[18][5] != ele[23][2];
    ele[18][5] != ele[23][3];
    ele[18][5] != ele[23][4];
    ele[18][5] != ele[23][5];
    ele[18][5] != ele[24][5];
    ele[18][5] != ele[25][5];
    ele[18][5] != ele[26][5];
    ele[18][5] != ele[27][5];
    ele[18][5] != ele[28][5];
    ele[18][5] != ele[29][5];
    ele[18][5] != ele[30][5];
    ele[18][5] != ele[31][5];
    ele[18][5] != ele[32][5];
    ele[18][5] != ele[33][5];
    ele[18][5] != ele[34][5];
    ele[18][5] != ele[35][5];
    ele[18][6] != ele[18][10];
    ele[18][6] != ele[18][11];
    ele[18][6] != ele[18][12];
    ele[18][6] != ele[18][13];
    ele[18][6] != ele[18][14];
    ele[18][6] != ele[18][15];
    ele[18][6] != ele[18][16];
    ele[18][6] != ele[18][17];
    ele[18][6] != ele[18][18];
    ele[18][6] != ele[18][19];
    ele[18][6] != ele[18][20];
    ele[18][6] != ele[18][21];
    ele[18][6] != ele[18][22];
    ele[18][6] != ele[18][23];
    ele[18][6] != ele[18][24];
    ele[18][6] != ele[18][25];
    ele[18][6] != ele[18][26];
    ele[18][6] != ele[18][27];
    ele[18][6] != ele[18][28];
    ele[18][6] != ele[18][29];
    ele[18][6] != ele[18][30];
    ele[18][6] != ele[18][31];
    ele[18][6] != ele[18][32];
    ele[18][6] != ele[18][33];
    ele[18][6] != ele[18][34];
    ele[18][6] != ele[18][35];
    ele[18][6] != ele[18][7];
    ele[18][6] != ele[18][8];
    ele[18][6] != ele[18][9];
    ele[18][6] != ele[19][10];
    ele[18][6] != ele[19][11];
    ele[18][6] != ele[19][6];
    ele[18][6] != ele[19][7];
    ele[18][6] != ele[19][8];
    ele[18][6] != ele[19][9];
    ele[18][6] != ele[20][10];
    ele[18][6] != ele[20][11];
    ele[18][6] != ele[20][6];
    ele[18][6] != ele[20][7];
    ele[18][6] != ele[20][8];
    ele[18][6] != ele[20][9];
    ele[18][6] != ele[21][10];
    ele[18][6] != ele[21][11];
    ele[18][6] != ele[21][6];
    ele[18][6] != ele[21][7];
    ele[18][6] != ele[21][8];
    ele[18][6] != ele[21][9];
    ele[18][6] != ele[22][10];
    ele[18][6] != ele[22][11];
    ele[18][6] != ele[22][6];
    ele[18][6] != ele[22][7];
    ele[18][6] != ele[22][8];
    ele[18][6] != ele[22][9];
    ele[18][6] != ele[23][10];
    ele[18][6] != ele[23][11];
    ele[18][6] != ele[23][6];
    ele[18][6] != ele[23][7];
    ele[18][6] != ele[23][8];
    ele[18][6] != ele[23][9];
    ele[18][6] != ele[24][6];
    ele[18][6] != ele[25][6];
    ele[18][6] != ele[26][6];
    ele[18][6] != ele[27][6];
    ele[18][6] != ele[28][6];
    ele[18][6] != ele[29][6];
    ele[18][6] != ele[30][6];
    ele[18][6] != ele[31][6];
    ele[18][6] != ele[32][6];
    ele[18][6] != ele[33][6];
    ele[18][6] != ele[34][6];
    ele[18][6] != ele[35][6];
    ele[18][7] != ele[18][10];
    ele[18][7] != ele[18][11];
    ele[18][7] != ele[18][12];
    ele[18][7] != ele[18][13];
    ele[18][7] != ele[18][14];
    ele[18][7] != ele[18][15];
    ele[18][7] != ele[18][16];
    ele[18][7] != ele[18][17];
    ele[18][7] != ele[18][18];
    ele[18][7] != ele[18][19];
    ele[18][7] != ele[18][20];
    ele[18][7] != ele[18][21];
    ele[18][7] != ele[18][22];
    ele[18][7] != ele[18][23];
    ele[18][7] != ele[18][24];
    ele[18][7] != ele[18][25];
    ele[18][7] != ele[18][26];
    ele[18][7] != ele[18][27];
    ele[18][7] != ele[18][28];
    ele[18][7] != ele[18][29];
    ele[18][7] != ele[18][30];
    ele[18][7] != ele[18][31];
    ele[18][7] != ele[18][32];
    ele[18][7] != ele[18][33];
    ele[18][7] != ele[18][34];
    ele[18][7] != ele[18][35];
    ele[18][7] != ele[18][8];
    ele[18][7] != ele[18][9];
    ele[18][7] != ele[19][10];
    ele[18][7] != ele[19][11];
    ele[18][7] != ele[19][6];
    ele[18][7] != ele[19][7];
    ele[18][7] != ele[19][8];
    ele[18][7] != ele[19][9];
    ele[18][7] != ele[20][10];
    ele[18][7] != ele[20][11];
    ele[18][7] != ele[20][6];
    ele[18][7] != ele[20][7];
    ele[18][7] != ele[20][8];
    ele[18][7] != ele[20][9];
    ele[18][7] != ele[21][10];
    ele[18][7] != ele[21][11];
    ele[18][7] != ele[21][6];
    ele[18][7] != ele[21][7];
    ele[18][7] != ele[21][8];
    ele[18][7] != ele[21][9];
    ele[18][7] != ele[22][10];
    ele[18][7] != ele[22][11];
    ele[18][7] != ele[22][6];
    ele[18][7] != ele[22][7];
    ele[18][7] != ele[22][8];
    ele[18][7] != ele[22][9];
    ele[18][7] != ele[23][10];
    ele[18][7] != ele[23][11];
    ele[18][7] != ele[23][6];
    ele[18][7] != ele[23][7];
    ele[18][7] != ele[23][8];
    ele[18][7] != ele[23][9];
    ele[18][7] != ele[24][7];
    ele[18][7] != ele[25][7];
    ele[18][7] != ele[26][7];
    ele[18][7] != ele[27][7];
    ele[18][7] != ele[28][7];
    ele[18][7] != ele[29][7];
    ele[18][7] != ele[30][7];
    ele[18][7] != ele[31][7];
    ele[18][7] != ele[32][7];
    ele[18][7] != ele[33][7];
    ele[18][7] != ele[34][7];
    ele[18][7] != ele[35][7];
    ele[18][8] != ele[18][10];
    ele[18][8] != ele[18][11];
    ele[18][8] != ele[18][12];
    ele[18][8] != ele[18][13];
    ele[18][8] != ele[18][14];
    ele[18][8] != ele[18][15];
    ele[18][8] != ele[18][16];
    ele[18][8] != ele[18][17];
    ele[18][8] != ele[18][18];
    ele[18][8] != ele[18][19];
    ele[18][8] != ele[18][20];
    ele[18][8] != ele[18][21];
    ele[18][8] != ele[18][22];
    ele[18][8] != ele[18][23];
    ele[18][8] != ele[18][24];
    ele[18][8] != ele[18][25];
    ele[18][8] != ele[18][26];
    ele[18][8] != ele[18][27];
    ele[18][8] != ele[18][28];
    ele[18][8] != ele[18][29];
    ele[18][8] != ele[18][30];
    ele[18][8] != ele[18][31];
    ele[18][8] != ele[18][32];
    ele[18][8] != ele[18][33];
    ele[18][8] != ele[18][34];
    ele[18][8] != ele[18][35];
    ele[18][8] != ele[18][9];
    ele[18][8] != ele[19][10];
    ele[18][8] != ele[19][11];
    ele[18][8] != ele[19][6];
    ele[18][8] != ele[19][7];
    ele[18][8] != ele[19][8];
    ele[18][8] != ele[19][9];
    ele[18][8] != ele[20][10];
    ele[18][8] != ele[20][11];
    ele[18][8] != ele[20][6];
    ele[18][8] != ele[20][7];
    ele[18][8] != ele[20][8];
    ele[18][8] != ele[20][9];
    ele[18][8] != ele[21][10];
    ele[18][8] != ele[21][11];
    ele[18][8] != ele[21][6];
    ele[18][8] != ele[21][7];
    ele[18][8] != ele[21][8];
    ele[18][8] != ele[21][9];
    ele[18][8] != ele[22][10];
    ele[18][8] != ele[22][11];
    ele[18][8] != ele[22][6];
    ele[18][8] != ele[22][7];
    ele[18][8] != ele[22][8];
    ele[18][8] != ele[22][9];
    ele[18][8] != ele[23][10];
    ele[18][8] != ele[23][11];
    ele[18][8] != ele[23][6];
    ele[18][8] != ele[23][7];
    ele[18][8] != ele[23][8];
    ele[18][8] != ele[23][9];
    ele[18][8] != ele[24][8];
    ele[18][8] != ele[25][8];
    ele[18][8] != ele[26][8];
    ele[18][8] != ele[27][8];
    ele[18][8] != ele[28][8];
    ele[18][8] != ele[29][8];
    ele[18][8] != ele[30][8];
    ele[18][8] != ele[31][8];
    ele[18][8] != ele[32][8];
    ele[18][8] != ele[33][8];
    ele[18][8] != ele[34][8];
    ele[18][8] != ele[35][8];
    ele[18][9] != ele[18][10];
    ele[18][9] != ele[18][11];
    ele[18][9] != ele[18][12];
    ele[18][9] != ele[18][13];
    ele[18][9] != ele[18][14];
    ele[18][9] != ele[18][15];
    ele[18][9] != ele[18][16];
    ele[18][9] != ele[18][17];
    ele[18][9] != ele[18][18];
    ele[18][9] != ele[18][19];
    ele[18][9] != ele[18][20];
    ele[18][9] != ele[18][21];
    ele[18][9] != ele[18][22];
    ele[18][9] != ele[18][23];
    ele[18][9] != ele[18][24];
    ele[18][9] != ele[18][25];
    ele[18][9] != ele[18][26];
    ele[18][9] != ele[18][27];
    ele[18][9] != ele[18][28];
    ele[18][9] != ele[18][29];
    ele[18][9] != ele[18][30];
    ele[18][9] != ele[18][31];
    ele[18][9] != ele[18][32];
    ele[18][9] != ele[18][33];
    ele[18][9] != ele[18][34];
    ele[18][9] != ele[18][35];
    ele[18][9] != ele[19][10];
    ele[18][9] != ele[19][11];
    ele[18][9] != ele[19][6];
    ele[18][9] != ele[19][7];
    ele[18][9] != ele[19][8];
    ele[18][9] != ele[19][9];
    ele[18][9] != ele[20][10];
    ele[18][9] != ele[20][11];
    ele[18][9] != ele[20][6];
    ele[18][9] != ele[20][7];
    ele[18][9] != ele[20][8];
    ele[18][9] != ele[20][9];
    ele[18][9] != ele[21][10];
    ele[18][9] != ele[21][11];
    ele[18][9] != ele[21][6];
    ele[18][9] != ele[21][7];
    ele[18][9] != ele[21][8];
    ele[18][9] != ele[21][9];
    ele[18][9] != ele[22][10];
    ele[18][9] != ele[22][11];
    ele[18][9] != ele[22][6];
    ele[18][9] != ele[22][7];
    ele[18][9] != ele[22][8];
    ele[18][9] != ele[22][9];
    ele[18][9] != ele[23][10];
    ele[18][9] != ele[23][11];
    ele[18][9] != ele[23][6];
    ele[18][9] != ele[23][7];
    ele[18][9] != ele[23][8];
    ele[18][9] != ele[23][9];
    ele[18][9] != ele[24][9];
    ele[18][9] != ele[25][9];
    ele[18][9] != ele[26][9];
    ele[18][9] != ele[27][9];
    ele[18][9] != ele[28][9];
    ele[18][9] != ele[29][9];
    ele[18][9] != ele[30][9];
    ele[18][9] != ele[31][9];
    ele[18][9] != ele[32][9];
    ele[18][9] != ele[33][9];
    ele[18][9] != ele[34][9];
    ele[18][9] != ele[35][9];
    ele[19][0] != ele[19][1];
    ele[19][0] != ele[19][10];
    ele[19][0] != ele[19][11];
    ele[19][0] != ele[19][12];
    ele[19][0] != ele[19][13];
    ele[19][0] != ele[19][14];
    ele[19][0] != ele[19][15];
    ele[19][0] != ele[19][16];
    ele[19][0] != ele[19][17];
    ele[19][0] != ele[19][18];
    ele[19][0] != ele[19][19];
    ele[19][0] != ele[19][2];
    ele[19][0] != ele[19][20];
    ele[19][0] != ele[19][21];
    ele[19][0] != ele[19][22];
    ele[19][0] != ele[19][23];
    ele[19][0] != ele[19][24];
    ele[19][0] != ele[19][25];
    ele[19][0] != ele[19][26];
    ele[19][0] != ele[19][27];
    ele[19][0] != ele[19][28];
    ele[19][0] != ele[19][29];
    ele[19][0] != ele[19][3];
    ele[19][0] != ele[19][30];
    ele[19][0] != ele[19][31];
    ele[19][0] != ele[19][32];
    ele[19][0] != ele[19][33];
    ele[19][0] != ele[19][34];
    ele[19][0] != ele[19][35];
    ele[19][0] != ele[19][4];
    ele[19][0] != ele[19][5];
    ele[19][0] != ele[19][6];
    ele[19][0] != ele[19][7];
    ele[19][0] != ele[19][8];
    ele[19][0] != ele[19][9];
    ele[19][0] != ele[20][0];
    ele[19][0] != ele[20][1];
    ele[19][0] != ele[20][2];
    ele[19][0] != ele[20][3];
    ele[19][0] != ele[20][4];
    ele[19][0] != ele[20][5];
    ele[19][0] != ele[21][0];
    ele[19][0] != ele[21][1];
    ele[19][0] != ele[21][2];
    ele[19][0] != ele[21][3];
    ele[19][0] != ele[21][4];
    ele[19][0] != ele[21][5];
    ele[19][0] != ele[22][0];
    ele[19][0] != ele[22][1];
    ele[19][0] != ele[22][2];
    ele[19][0] != ele[22][3];
    ele[19][0] != ele[22][4];
    ele[19][0] != ele[22][5];
    ele[19][0] != ele[23][0];
    ele[19][0] != ele[23][1];
    ele[19][0] != ele[23][2];
    ele[19][0] != ele[23][3];
    ele[19][0] != ele[23][4];
    ele[19][0] != ele[23][5];
    ele[19][0] != ele[24][0];
    ele[19][0] != ele[25][0];
    ele[19][0] != ele[26][0];
    ele[19][0] != ele[27][0];
    ele[19][0] != ele[28][0];
    ele[19][0] != ele[29][0];
    ele[19][0] != ele[30][0];
    ele[19][0] != ele[31][0];
    ele[19][0] != ele[32][0];
    ele[19][0] != ele[33][0];
    ele[19][0] != ele[34][0];
    ele[19][0] != ele[35][0];
    ele[19][1] != ele[19][10];
    ele[19][1] != ele[19][11];
    ele[19][1] != ele[19][12];
    ele[19][1] != ele[19][13];
    ele[19][1] != ele[19][14];
    ele[19][1] != ele[19][15];
    ele[19][1] != ele[19][16];
    ele[19][1] != ele[19][17];
    ele[19][1] != ele[19][18];
    ele[19][1] != ele[19][19];
    ele[19][1] != ele[19][2];
    ele[19][1] != ele[19][20];
    ele[19][1] != ele[19][21];
    ele[19][1] != ele[19][22];
    ele[19][1] != ele[19][23];
    ele[19][1] != ele[19][24];
    ele[19][1] != ele[19][25];
    ele[19][1] != ele[19][26];
    ele[19][1] != ele[19][27];
    ele[19][1] != ele[19][28];
    ele[19][1] != ele[19][29];
    ele[19][1] != ele[19][3];
    ele[19][1] != ele[19][30];
    ele[19][1] != ele[19][31];
    ele[19][1] != ele[19][32];
    ele[19][1] != ele[19][33];
    ele[19][1] != ele[19][34];
    ele[19][1] != ele[19][35];
    ele[19][1] != ele[19][4];
    ele[19][1] != ele[19][5];
    ele[19][1] != ele[19][6];
    ele[19][1] != ele[19][7];
    ele[19][1] != ele[19][8];
    ele[19][1] != ele[19][9];
    ele[19][1] != ele[20][0];
    ele[19][1] != ele[20][1];
    ele[19][1] != ele[20][2];
    ele[19][1] != ele[20][3];
    ele[19][1] != ele[20][4];
    ele[19][1] != ele[20][5];
    ele[19][1] != ele[21][0];
    ele[19][1] != ele[21][1];
    ele[19][1] != ele[21][2];
    ele[19][1] != ele[21][3];
    ele[19][1] != ele[21][4];
    ele[19][1] != ele[21][5];
    ele[19][1] != ele[22][0];
    ele[19][1] != ele[22][1];
    ele[19][1] != ele[22][2];
    ele[19][1] != ele[22][3];
    ele[19][1] != ele[22][4];
    ele[19][1] != ele[22][5];
    ele[19][1] != ele[23][0];
    ele[19][1] != ele[23][1];
    ele[19][1] != ele[23][2];
    ele[19][1] != ele[23][3];
    ele[19][1] != ele[23][4];
    ele[19][1] != ele[23][5];
    ele[19][1] != ele[24][1];
    ele[19][1] != ele[25][1];
    ele[19][1] != ele[26][1];
    ele[19][1] != ele[27][1];
    ele[19][1] != ele[28][1];
    ele[19][1] != ele[29][1];
    ele[19][1] != ele[30][1];
    ele[19][1] != ele[31][1];
    ele[19][1] != ele[32][1];
    ele[19][1] != ele[33][1];
    ele[19][1] != ele[34][1];
    ele[19][1] != ele[35][1];
    ele[19][10] != ele[19][11];
    ele[19][10] != ele[19][12];
    ele[19][10] != ele[19][13];
    ele[19][10] != ele[19][14];
    ele[19][10] != ele[19][15];
    ele[19][10] != ele[19][16];
    ele[19][10] != ele[19][17];
    ele[19][10] != ele[19][18];
    ele[19][10] != ele[19][19];
    ele[19][10] != ele[19][20];
    ele[19][10] != ele[19][21];
    ele[19][10] != ele[19][22];
    ele[19][10] != ele[19][23];
    ele[19][10] != ele[19][24];
    ele[19][10] != ele[19][25];
    ele[19][10] != ele[19][26];
    ele[19][10] != ele[19][27];
    ele[19][10] != ele[19][28];
    ele[19][10] != ele[19][29];
    ele[19][10] != ele[19][30];
    ele[19][10] != ele[19][31];
    ele[19][10] != ele[19][32];
    ele[19][10] != ele[19][33];
    ele[19][10] != ele[19][34];
    ele[19][10] != ele[19][35];
    ele[19][10] != ele[20][10];
    ele[19][10] != ele[20][11];
    ele[19][10] != ele[20][6];
    ele[19][10] != ele[20][7];
    ele[19][10] != ele[20][8];
    ele[19][10] != ele[20][9];
    ele[19][10] != ele[21][10];
    ele[19][10] != ele[21][11];
    ele[19][10] != ele[21][6];
    ele[19][10] != ele[21][7];
    ele[19][10] != ele[21][8];
    ele[19][10] != ele[21][9];
    ele[19][10] != ele[22][10];
    ele[19][10] != ele[22][11];
    ele[19][10] != ele[22][6];
    ele[19][10] != ele[22][7];
    ele[19][10] != ele[22][8];
    ele[19][10] != ele[22][9];
    ele[19][10] != ele[23][10];
    ele[19][10] != ele[23][11];
    ele[19][10] != ele[23][6];
    ele[19][10] != ele[23][7];
    ele[19][10] != ele[23][8];
    ele[19][10] != ele[23][9];
    ele[19][10] != ele[24][10];
    ele[19][10] != ele[25][10];
    ele[19][10] != ele[26][10];
    ele[19][10] != ele[27][10];
    ele[19][10] != ele[28][10];
    ele[19][10] != ele[29][10];
    ele[19][10] != ele[30][10];
    ele[19][10] != ele[31][10];
    ele[19][10] != ele[32][10];
    ele[19][10] != ele[33][10];
    ele[19][10] != ele[34][10];
    ele[19][10] != ele[35][10];
    ele[19][11] != ele[19][12];
    ele[19][11] != ele[19][13];
    ele[19][11] != ele[19][14];
    ele[19][11] != ele[19][15];
    ele[19][11] != ele[19][16];
    ele[19][11] != ele[19][17];
    ele[19][11] != ele[19][18];
    ele[19][11] != ele[19][19];
    ele[19][11] != ele[19][20];
    ele[19][11] != ele[19][21];
    ele[19][11] != ele[19][22];
    ele[19][11] != ele[19][23];
    ele[19][11] != ele[19][24];
    ele[19][11] != ele[19][25];
    ele[19][11] != ele[19][26];
    ele[19][11] != ele[19][27];
    ele[19][11] != ele[19][28];
    ele[19][11] != ele[19][29];
    ele[19][11] != ele[19][30];
    ele[19][11] != ele[19][31];
    ele[19][11] != ele[19][32];
    ele[19][11] != ele[19][33];
    ele[19][11] != ele[19][34];
    ele[19][11] != ele[19][35];
    ele[19][11] != ele[20][10];
    ele[19][11] != ele[20][11];
    ele[19][11] != ele[20][6];
    ele[19][11] != ele[20][7];
    ele[19][11] != ele[20][8];
    ele[19][11] != ele[20][9];
    ele[19][11] != ele[21][10];
    ele[19][11] != ele[21][11];
    ele[19][11] != ele[21][6];
    ele[19][11] != ele[21][7];
    ele[19][11] != ele[21][8];
    ele[19][11] != ele[21][9];
    ele[19][11] != ele[22][10];
    ele[19][11] != ele[22][11];
    ele[19][11] != ele[22][6];
    ele[19][11] != ele[22][7];
    ele[19][11] != ele[22][8];
    ele[19][11] != ele[22][9];
    ele[19][11] != ele[23][10];
    ele[19][11] != ele[23][11];
    ele[19][11] != ele[23][6];
    ele[19][11] != ele[23][7];
    ele[19][11] != ele[23][8];
    ele[19][11] != ele[23][9];
    ele[19][11] != ele[24][11];
    ele[19][11] != ele[25][11];
    ele[19][11] != ele[26][11];
    ele[19][11] != ele[27][11];
    ele[19][11] != ele[28][11];
    ele[19][11] != ele[29][11];
    ele[19][11] != ele[30][11];
    ele[19][11] != ele[31][11];
    ele[19][11] != ele[32][11];
    ele[19][11] != ele[33][11];
    ele[19][11] != ele[34][11];
    ele[19][11] != ele[35][11];
    ele[19][12] != ele[19][13];
    ele[19][12] != ele[19][14];
    ele[19][12] != ele[19][15];
    ele[19][12] != ele[19][16];
    ele[19][12] != ele[19][17];
    ele[19][12] != ele[19][18];
    ele[19][12] != ele[19][19];
    ele[19][12] != ele[19][20];
    ele[19][12] != ele[19][21];
    ele[19][12] != ele[19][22];
    ele[19][12] != ele[19][23];
    ele[19][12] != ele[19][24];
    ele[19][12] != ele[19][25];
    ele[19][12] != ele[19][26];
    ele[19][12] != ele[19][27];
    ele[19][12] != ele[19][28];
    ele[19][12] != ele[19][29];
    ele[19][12] != ele[19][30];
    ele[19][12] != ele[19][31];
    ele[19][12] != ele[19][32];
    ele[19][12] != ele[19][33];
    ele[19][12] != ele[19][34];
    ele[19][12] != ele[19][35];
    ele[19][12] != ele[20][12];
    ele[19][12] != ele[20][13];
    ele[19][12] != ele[20][14];
    ele[19][12] != ele[20][15];
    ele[19][12] != ele[20][16];
    ele[19][12] != ele[20][17];
    ele[19][12] != ele[21][12];
    ele[19][12] != ele[21][13];
    ele[19][12] != ele[21][14];
    ele[19][12] != ele[21][15];
    ele[19][12] != ele[21][16];
    ele[19][12] != ele[21][17];
    ele[19][12] != ele[22][12];
    ele[19][12] != ele[22][13];
    ele[19][12] != ele[22][14];
    ele[19][12] != ele[22][15];
    ele[19][12] != ele[22][16];
    ele[19][12] != ele[22][17];
    ele[19][12] != ele[23][12];
    ele[19][12] != ele[23][13];
    ele[19][12] != ele[23][14];
    ele[19][12] != ele[23][15];
    ele[19][12] != ele[23][16];
    ele[19][12] != ele[23][17];
    ele[19][12] != ele[24][12];
    ele[19][12] != ele[25][12];
    ele[19][12] != ele[26][12];
    ele[19][12] != ele[27][12];
    ele[19][12] != ele[28][12];
    ele[19][12] != ele[29][12];
    ele[19][12] != ele[30][12];
    ele[19][12] != ele[31][12];
    ele[19][12] != ele[32][12];
    ele[19][12] != ele[33][12];
    ele[19][12] != ele[34][12];
    ele[19][12] != ele[35][12];
    ele[19][13] != ele[19][14];
    ele[19][13] != ele[19][15];
    ele[19][13] != ele[19][16];
    ele[19][13] != ele[19][17];
    ele[19][13] != ele[19][18];
    ele[19][13] != ele[19][19];
    ele[19][13] != ele[19][20];
    ele[19][13] != ele[19][21];
    ele[19][13] != ele[19][22];
    ele[19][13] != ele[19][23];
    ele[19][13] != ele[19][24];
    ele[19][13] != ele[19][25];
    ele[19][13] != ele[19][26];
    ele[19][13] != ele[19][27];
    ele[19][13] != ele[19][28];
    ele[19][13] != ele[19][29];
    ele[19][13] != ele[19][30];
    ele[19][13] != ele[19][31];
    ele[19][13] != ele[19][32];
    ele[19][13] != ele[19][33];
    ele[19][13] != ele[19][34];
    ele[19][13] != ele[19][35];
    ele[19][13] != ele[20][12];
    ele[19][13] != ele[20][13];
    ele[19][13] != ele[20][14];
    ele[19][13] != ele[20][15];
    ele[19][13] != ele[20][16];
    ele[19][13] != ele[20][17];
    ele[19][13] != ele[21][12];
    ele[19][13] != ele[21][13];
    ele[19][13] != ele[21][14];
    ele[19][13] != ele[21][15];
    ele[19][13] != ele[21][16];
    ele[19][13] != ele[21][17];
    ele[19][13] != ele[22][12];
    ele[19][13] != ele[22][13];
    ele[19][13] != ele[22][14];
    ele[19][13] != ele[22][15];
    ele[19][13] != ele[22][16];
    ele[19][13] != ele[22][17];
    ele[19][13] != ele[23][12];
    ele[19][13] != ele[23][13];
    ele[19][13] != ele[23][14];
    ele[19][13] != ele[23][15];
    ele[19][13] != ele[23][16];
    ele[19][13] != ele[23][17];
    ele[19][13] != ele[24][13];
    ele[19][13] != ele[25][13];
    ele[19][13] != ele[26][13];
    ele[19][13] != ele[27][13];
    ele[19][13] != ele[28][13];
    ele[19][13] != ele[29][13];
    ele[19][13] != ele[30][13];
    ele[19][13] != ele[31][13];
    ele[19][13] != ele[32][13];
    ele[19][13] != ele[33][13];
    ele[19][13] != ele[34][13];
    ele[19][13] != ele[35][13];
    ele[19][14] != ele[19][15];
    ele[19][14] != ele[19][16];
    ele[19][14] != ele[19][17];
    ele[19][14] != ele[19][18];
    ele[19][14] != ele[19][19];
    ele[19][14] != ele[19][20];
    ele[19][14] != ele[19][21];
    ele[19][14] != ele[19][22];
    ele[19][14] != ele[19][23];
    ele[19][14] != ele[19][24];
    ele[19][14] != ele[19][25];
    ele[19][14] != ele[19][26];
    ele[19][14] != ele[19][27];
    ele[19][14] != ele[19][28];
    ele[19][14] != ele[19][29];
    ele[19][14] != ele[19][30];
    ele[19][14] != ele[19][31];
    ele[19][14] != ele[19][32];
    ele[19][14] != ele[19][33];
    ele[19][14] != ele[19][34];
    ele[19][14] != ele[19][35];
    ele[19][14] != ele[20][12];
    ele[19][14] != ele[20][13];
    ele[19][14] != ele[20][14];
    ele[19][14] != ele[20][15];
    ele[19][14] != ele[20][16];
    ele[19][14] != ele[20][17];
    ele[19][14] != ele[21][12];
    ele[19][14] != ele[21][13];
    ele[19][14] != ele[21][14];
    ele[19][14] != ele[21][15];
    ele[19][14] != ele[21][16];
    ele[19][14] != ele[21][17];
    ele[19][14] != ele[22][12];
    ele[19][14] != ele[22][13];
    ele[19][14] != ele[22][14];
    ele[19][14] != ele[22][15];
    ele[19][14] != ele[22][16];
    ele[19][14] != ele[22][17];
    ele[19][14] != ele[23][12];
    ele[19][14] != ele[23][13];
    ele[19][14] != ele[23][14];
    ele[19][14] != ele[23][15];
    ele[19][14] != ele[23][16];
    ele[19][14] != ele[23][17];
    ele[19][14] != ele[24][14];
    ele[19][14] != ele[25][14];
    ele[19][14] != ele[26][14];
    ele[19][14] != ele[27][14];
    ele[19][14] != ele[28][14];
    ele[19][14] != ele[29][14];
    ele[19][14] != ele[30][14];
    ele[19][14] != ele[31][14];
    ele[19][14] != ele[32][14];
    ele[19][14] != ele[33][14];
    ele[19][14] != ele[34][14];
    ele[19][14] != ele[35][14];
    ele[19][15] != ele[19][16];
    ele[19][15] != ele[19][17];
    ele[19][15] != ele[19][18];
    ele[19][15] != ele[19][19];
    ele[19][15] != ele[19][20];
    ele[19][15] != ele[19][21];
    ele[19][15] != ele[19][22];
    ele[19][15] != ele[19][23];
    ele[19][15] != ele[19][24];
    ele[19][15] != ele[19][25];
    ele[19][15] != ele[19][26];
    ele[19][15] != ele[19][27];
    ele[19][15] != ele[19][28];
    ele[19][15] != ele[19][29];
    ele[19][15] != ele[19][30];
    ele[19][15] != ele[19][31];
    ele[19][15] != ele[19][32];
    ele[19][15] != ele[19][33];
    ele[19][15] != ele[19][34];
    ele[19][15] != ele[19][35];
    ele[19][15] != ele[20][12];
    ele[19][15] != ele[20][13];
    ele[19][15] != ele[20][14];
    ele[19][15] != ele[20][15];
    ele[19][15] != ele[20][16];
    ele[19][15] != ele[20][17];
    ele[19][15] != ele[21][12];
    ele[19][15] != ele[21][13];
    ele[19][15] != ele[21][14];
    ele[19][15] != ele[21][15];
    ele[19][15] != ele[21][16];
    ele[19][15] != ele[21][17];
    ele[19][15] != ele[22][12];
    ele[19][15] != ele[22][13];
    ele[19][15] != ele[22][14];
    ele[19][15] != ele[22][15];
    ele[19][15] != ele[22][16];
    ele[19][15] != ele[22][17];
    ele[19][15] != ele[23][12];
    ele[19][15] != ele[23][13];
    ele[19][15] != ele[23][14];
    ele[19][15] != ele[23][15];
    ele[19][15] != ele[23][16];
    ele[19][15] != ele[23][17];
    ele[19][15] != ele[24][15];
    ele[19][15] != ele[25][15];
    ele[19][15] != ele[26][15];
    ele[19][15] != ele[27][15];
    ele[19][15] != ele[28][15];
    ele[19][15] != ele[29][15];
    ele[19][15] != ele[30][15];
    ele[19][15] != ele[31][15];
    ele[19][15] != ele[32][15];
    ele[19][15] != ele[33][15];
    ele[19][15] != ele[34][15];
    ele[19][15] != ele[35][15];
    ele[19][16] != ele[19][17];
    ele[19][16] != ele[19][18];
    ele[19][16] != ele[19][19];
    ele[19][16] != ele[19][20];
    ele[19][16] != ele[19][21];
    ele[19][16] != ele[19][22];
    ele[19][16] != ele[19][23];
    ele[19][16] != ele[19][24];
    ele[19][16] != ele[19][25];
    ele[19][16] != ele[19][26];
    ele[19][16] != ele[19][27];
    ele[19][16] != ele[19][28];
    ele[19][16] != ele[19][29];
    ele[19][16] != ele[19][30];
    ele[19][16] != ele[19][31];
    ele[19][16] != ele[19][32];
    ele[19][16] != ele[19][33];
    ele[19][16] != ele[19][34];
    ele[19][16] != ele[19][35];
    ele[19][16] != ele[20][12];
    ele[19][16] != ele[20][13];
    ele[19][16] != ele[20][14];
    ele[19][16] != ele[20][15];
    ele[19][16] != ele[20][16];
    ele[19][16] != ele[20][17];
    ele[19][16] != ele[21][12];
    ele[19][16] != ele[21][13];
    ele[19][16] != ele[21][14];
    ele[19][16] != ele[21][15];
    ele[19][16] != ele[21][16];
    ele[19][16] != ele[21][17];
    ele[19][16] != ele[22][12];
    ele[19][16] != ele[22][13];
    ele[19][16] != ele[22][14];
    ele[19][16] != ele[22][15];
    ele[19][16] != ele[22][16];
    ele[19][16] != ele[22][17];
    ele[19][16] != ele[23][12];
    ele[19][16] != ele[23][13];
    ele[19][16] != ele[23][14];
    ele[19][16] != ele[23][15];
    ele[19][16] != ele[23][16];
    ele[19][16] != ele[23][17];
    ele[19][16] != ele[24][16];
    ele[19][16] != ele[25][16];
    ele[19][16] != ele[26][16];
    ele[19][16] != ele[27][16];
    ele[19][16] != ele[28][16];
    ele[19][16] != ele[29][16];
    ele[19][16] != ele[30][16];
    ele[19][16] != ele[31][16];
    ele[19][16] != ele[32][16];
    ele[19][16] != ele[33][16];
    ele[19][16] != ele[34][16];
    ele[19][16] != ele[35][16];
    ele[19][17] != ele[19][18];
    ele[19][17] != ele[19][19];
    ele[19][17] != ele[19][20];
    ele[19][17] != ele[19][21];
    ele[19][17] != ele[19][22];
    ele[19][17] != ele[19][23];
    ele[19][17] != ele[19][24];
    ele[19][17] != ele[19][25];
    ele[19][17] != ele[19][26];
    ele[19][17] != ele[19][27];
    ele[19][17] != ele[19][28];
    ele[19][17] != ele[19][29];
    ele[19][17] != ele[19][30];
    ele[19][17] != ele[19][31];
    ele[19][17] != ele[19][32];
    ele[19][17] != ele[19][33];
    ele[19][17] != ele[19][34];
    ele[19][17] != ele[19][35];
    ele[19][17] != ele[20][12];
    ele[19][17] != ele[20][13];
    ele[19][17] != ele[20][14];
    ele[19][17] != ele[20][15];
    ele[19][17] != ele[20][16];
    ele[19][17] != ele[20][17];
    ele[19][17] != ele[21][12];
    ele[19][17] != ele[21][13];
    ele[19][17] != ele[21][14];
    ele[19][17] != ele[21][15];
    ele[19][17] != ele[21][16];
    ele[19][17] != ele[21][17];
    ele[19][17] != ele[22][12];
    ele[19][17] != ele[22][13];
    ele[19][17] != ele[22][14];
    ele[19][17] != ele[22][15];
    ele[19][17] != ele[22][16];
    ele[19][17] != ele[22][17];
    ele[19][17] != ele[23][12];
    ele[19][17] != ele[23][13];
    ele[19][17] != ele[23][14];
    ele[19][17] != ele[23][15];
    ele[19][17] != ele[23][16];
    ele[19][17] != ele[23][17];
    ele[19][17] != ele[24][17];
    ele[19][17] != ele[25][17];
    ele[19][17] != ele[26][17];
    ele[19][17] != ele[27][17];
    ele[19][17] != ele[28][17];
    ele[19][17] != ele[29][17];
    ele[19][17] != ele[30][17];
    ele[19][17] != ele[31][17];
    ele[19][17] != ele[32][17];
    ele[19][17] != ele[33][17];
    ele[19][17] != ele[34][17];
    ele[19][17] != ele[35][17];
    ele[19][18] != ele[19][19];
    ele[19][18] != ele[19][20];
    ele[19][18] != ele[19][21];
    ele[19][18] != ele[19][22];
    ele[19][18] != ele[19][23];
    ele[19][18] != ele[19][24];
    ele[19][18] != ele[19][25];
    ele[19][18] != ele[19][26];
    ele[19][18] != ele[19][27];
    ele[19][18] != ele[19][28];
    ele[19][18] != ele[19][29];
    ele[19][18] != ele[19][30];
    ele[19][18] != ele[19][31];
    ele[19][18] != ele[19][32];
    ele[19][18] != ele[19][33];
    ele[19][18] != ele[19][34];
    ele[19][18] != ele[19][35];
    ele[19][18] != ele[20][18];
    ele[19][18] != ele[20][19];
    ele[19][18] != ele[20][20];
    ele[19][18] != ele[20][21];
    ele[19][18] != ele[20][22];
    ele[19][18] != ele[20][23];
    ele[19][18] != ele[21][18];
    ele[19][18] != ele[21][19];
    ele[19][18] != ele[21][20];
    ele[19][18] != ele[21][21];
    ele[19][18] != ele[21][22];
    ele[19][18] != ele[21][23];
    ele[19][18] != ele[22][18];
    ele[19][18] != ele[22][19];
    ele[19][18] != ele[22][20];
    ele[19][18] != ele[22][21];
    ele[19][18] != ele[22][22];
    ele[19][18] != ele[22][23];
    ele[19][18] != ele[23][18];
    ele[19][18] != ele[23][19];
    ele[19][18] != ele[23][20];
    ele[19][18] != ele[23][21];
    ele[19][18] != ele[23][22];
    ele[19][18] != ele[23][23];
    ele[19][18] != ele[24][18];
    ele[19][18] != ele[25][18];
    ele[19][18] != ele[26][18];
    ele[19][18] != ele[27][18];
    ele[19][18] != ele[28][18];
    ele[19][18] != ele[29][18];
    ele[19][18] != ele[30][18];
    ele[19][18] != ele[31][18];
    ele[19][18] != ele[32][18];
    ele[19][18] != ele[33][18];
    ele[19][18] != ele[34][18];
    ele[19][18] != ele[35][18];
    ele[19][19] != ele[19][20];
    ele[19][19] != ele[19][21];
    ele[19][19] != ele[19][22];
    ele[19][19] != ele[19][23];
    ele[19][19] != ele[19][24];
    ele[19][19] != ele[19][25];
    ele[19][19] != ele[19][26];
    ele[19][19] != ele[19][27];
    ele[19][19] != ele[19][28];
    ele[19][19] != ele[19][29];
    ele[19][19] != ele[19][30];
    ele[19][19] != ele[19][31];
    ele[19][19] != ele[19][32];
    ele[19][19] != ele[19][33];
    ele[19][19] != ele[19][34];
    ele[19][19] != ele[19][35];
    ele[19][19] != ele[20][18];
    ele[19][19] != ele[20][19];
    ele[19][19] != ele[20][20];
    ele[19][19] != ele[20][21];
    ele[19][19] != ele[20][22];
    ele[19][19] != ele[20][23];
    ele[19][19] != ele[21][18];
    ele[19][19] != ele[21][19];
    ele[19][19] != ele[21][20];
    ele[19][19] != ele[21][21];
    ele[19][19] != ele[21][22];
    ele[19][19] != ele[21][23];
    ele[19][19] != ele[22][18];
    ele[19][19] != ele[22][19];
    ele[19][19] != ele[22][20];
    ele[19][19] != ele[22][21];
    ele[19][19] != ele[22][22];
    ele[19][19] != ele[22][23];
    ele[19][19] != ele[23][18];
    ele[19][19] != ele[23][19];
    ele[19][19] != ele[23][20];
    ele[19][19] != ele[23][21];
    ele[19][19] != ele[23][22];
    ele[19][19] != ele[23][23];
    ele[19][19] != ele[24][19];
    ele[19][19] != ele[25][19];
    ele[19][19] != ele[26][19];
    ele[19][19] != ele[27][19];
    ele[19][19] != ele[28][19];
    ele[19][19] != ele[29][19];
    ele[19][19] != ele[30][19];
    ele[19][19] != ele[31][19];
    ele[19][19] != ele[32][19];
    ele[19][19] != ele[33][19];
    ele[19][19] != ele[34][19];
    ele[19][19] != ele[35][19];
    ele[19][2] != ele[19][10];
    ele[19][2] != ele[19][11];
    ele[19][2] != ele[19][12];
    ele[19][2] != ele[19][13];
    ele[19][2] != ele[19][14];
    ele[19][2] != ele[19][15];
    ele[19][2] != ele[19][16];
    ele[19][2] != ele[19][17];
    ele[19][2] != ele[19][18];
    ele[19][2] != ele[19][19];
    ele[19][2] != ele[19][20];
    ele[19][2] != ele[19][21];
    ele[19][2] != ele[19][22];
    ele[19][2] != ele[19][23];
    ele[19][2] != ele[19][24];
    ele[19][2] != ele[19][25];
    ele[19][2] != ele[19][26];
    ele[19][2] != ele[19][27];
    ele[19][2] != ele[19][28];
    ele[19][2] != ele[19][29];
    ele[19][2] != ele[19][3];
    ele[19][2] != ele[19][30];
    ele[19][2] != ele[19][31];
    ele[19][2] != ele[19][32];
    ele[19][2] != ele[19][33];
    ele[19][2] != ele[19][34];
    ele[19][2] != ele[19][35];
    ele[19][2] != ele[19][4];
    ele[19][2] != ele[19][5];
    ele[19][2] != ele[19][6];
    ele[19][2] != ele[19][7];
    ele[19][2] != ele[19][8];
    ele[19][2] != ele[19][9];
    ele[19][2] != ele[20][0];
    ele[19][2] != ele[20][1];
    ele[19][2] != ele[20][2];
    ele[19][2] != ele[20][3];
    ele[19][2] != ele[20][4];
    ele[19][2] != ele[20][5];
    ele[19][2] != ele[21][0];
    ele[19][2] != ele[21][1];
    ele[19][2] != ele[21][2];
    ele[19][2] != ele[21][3];
    ele[19][2] != ele[21][4];
    ele[19][2] != ele[21][5];
    ele[19][2] != ele[22][0];
    ele[19][2] != ele[22][1];
    ele[19][2] != ele[22][2];
    ele[19][2] != ele[22][3];
    ele[19][2] != ele[22][4];
    ele[19][2] != ele[22][5];
    ele[19][2] != ele[23][0];
    ele[19][2] != ele[23][1];
    ele[19][2] != ele[23][2];
    ele[19][2] != ele[23][3];
    ele[19][2] != ele[23][4];
    ele[19][2] != ele[23][5];
    ele[19][2] != ele[24][2];
    ele[19][2] != ele[25][2];
    ele[19][2] != ele[26][2];
    ele[19][2] != ele[27][2];
    ele[19][2] != ele[28][2];
    ele[19][2] != ele[29][2];
    ele[19][2] != ele[30][2];
    ele[19][2] != ele[31][2];
    ele[19][2] != ele[32][2];
    ele[19][2] != ele[33][2];
    ele[19][2] != ele[34][2];
    ele[19][2] != ele[35][2];
    ele[19][20] != ele[19][21];
    ele[19][20] != ele[19][22];
    ele[19][20] != ele[19][23];
    ele[19][20] != ele[19][24];
    ele[19][20] != ele[19][25];
    ele[19][20] != ele[19][26];
    ele[19][20] != ele[19][27];
    ele[19][20] != ele[19][28];
    ele[19][20] != ele[19][29];
    ele[19][20] != ele[19][30];
    ele[19][20] != ele[19][31];
    ele[19][20] != ele[19][32];
    ele[19][20] != ele[19][33];
    ele[19][20] != ele[19][34];
    ele[19][20] != ele[19][35];
    ele[19][20] != ele[20][18];
    ele[19][20] != ele[20][19];
    ele[19][20] != ele[20][20];
    ele[19][20] != ele[20][21];
    ele[19][20] != ele[20][22];
    ele[19][20] != ele[20][23];
    ele[19][20] != ele[21][18];
    ele[19][20] != ele[21][19];
    ele[19][20] != ele[21][20];
    ele[19][20] != ele[21][21];
    ele[19][20] != ele[21][22];
    ele[19][20] != ele[21][23];
    ele[19][20] != ele[22][18];
    ele[19][20] != ele[22][19];
    ele[19][20] != ele[22][20];
    ele[19][20] != ele[22][21];
    ele[19][20] != ele[22][22];
    ele[19][20] != ele[22][23];
    ele[19][20] != ele[23][18];
    ele[19][20] != ele[23][19];
    ele[19][20] != ele[23][20];
    ele[19][20] != ele[23][21];
    ele[19][20] != ele[23][22];
    ele[19][20] != ele[23][23];
    ele[19][20] != ele[24][20];
    ele[19][20] != ele[25][20];
    ele[19][20] != ele[26][20];
    ele[19][20] != ele[27][20];
    ele[19][20] != ele[28][20];
    ele[19][20] != ele[29][20];
    ele[19][20] != ele[30][20];
    ele[19][20] != ele[31][20];
    ele[19][20] != ele[32][20];
    ele[19][20] != ele[33][20];
    ele[19][20] != ele[34][20];
    ele[19][20] != ele[35][20];
    ele[19][21] != ele[19][22];
    ele[19][21] != ele[19][23];
    ele[19][21] != ele[19][24];
    ele[19][21] != ele[19][25];
    ele[19][21] != ele[19][26];
    ele[19][21] != ele[19][27];
    ele[19][21] != ele[19][28];
    ele[19][21] != ele[19][29];
    ele[19][21] != ele[19][30];
    ele[19][21] != ele[19][31];
    ele[19][21] != ele[19][32];
    ele[19][21] != ele[19][33];
    ele[19][21] != ele[19][34];
    ele[19][21] != ele[19][35];
    ele[19][21] != ele[20][18];
    ele[19][21] != ele[20][19];
    ele[19][21] != ele[20][20];
    ele[19][21] != ele[20][21];
    ele[19][21] != ele[20][22];
    ele[19][21] != ele[20][23];
    ele[19][21] != ele[21][18];
    ele[19][21] != ele[21][19];
    ele[19][21] != ele[21][20];
    ele[19][21] != ele[21][21];
    ele[19][21] != ele[21][22];
    ele[19][21] != ele[21][23];
    ele[19][21] != ele[22][18];
    ele[19][21] != ele[22][19];
    ele[19][21] != ele[22][20];
    ele[19][21] != ele[22][21];
    ele[19][21] != ele[22][22];
    ele[19][21] != ele[22][23];
    ele[19][21] != ele[23][18];
    ele[19][21] != ele[23][19];
    ele[19][21] != ele[23][20];
    ele[19][21] != ele[23][21];
    ele[19][21] != ele[23][22];
    ele[19][21] != ele[23][23];
    ele[19][21] != ele[24][21];
    ele[19][21] != ele[25][21];
    ele[19][21] != ele[26][21];
    ele[19][21] != ele[27][21];
    ele[19][21] != ele[28][21];
    ele[19][21] != ele[29][21];
    ele[19][21] != ele[30][21];
    ele[19][21] != ele[31][21];
    ele[19][21] != ele[32][21];
    ele[19][21] != ele[33][21];
    ele[19][21] != ele[34][21];
    ele[19][21] != ele[35][21];
    ele[19][22] != ele[19][23];
    ele[19][22] != ele[19][24];
    ele[19][22] != ele[19][25];
    ele[19][22] != ele[19][26];
    ele[19][22] != ele[19][27];
    ele[19][22] != ele[19][28];
    ele[19][22] != ele[19][29];
    ele[19][22] != ele[19][30];
    ele[19][22] != ele[19][31];
    ele[19][22] != ele[19][32];
    ele[19][22] != ele[19][33];
    ele[19][22] != ele[19][34];
    ele[19][22] != ele[19][35];
    ele[19][22] != ele[20][18];
    ele[19][22] != ele[20][19];
    ele[19][22] != ele[20][20];
    ele[19][22] != ele[20][21];
    ele[19][22] != ele[20][22];
    ele[19][22] != ele[20][23];
    ele[19][22] != ele[21][18];
    ele[19][22] != ele[21][19];
    ele[19][22] != ele[21][20];
    ele[19][22] != ele[21][21];
    ele[19][22] != ele[21][22];
    ele[19][22] != ele[21][23];
    ele[19][22] != ele[22][18];
    ele[19][22] != ele[22][19];
    ele[19][22] != ele[22][20];
    ele[19][22] != ele[22][21];
    ele[19][22] != ele[22][22];
    ele[19][22] != ele[22][23];
    ele[19][22] != ele[23][18];
    ele[19][22] != ele[23][19];
    ele[19][22] != ele[23][20];
    ele[19][22] != ele[23][21];
    ele[19][22] != ele[23][22];
    ele[19][22] != ele[23][23];
    ele[19][22] != ele[24][22];
    ele[19][22] != ele[25][22];
    ele[19][22] != ele[26][22];
    ele[19][22] != ele[27][22];
    ele[19][22] != ele[28][22];
    ele[19][22] != ele[29][22];
    ele[19][22] != ele[30][22];
    ele[19][22] != ele[31][22];
    ele[19][22] != ele[32][22];
    ele[19][22] != ele[33][22];
    ele[19][22] != ele[34][22];
    ele[19][22] != ele[35][22];
    ele[19][23] != ele[19][24];
    ele[19][23] != ele[19][25];
    ele[19][23] != ele[19][26];
    ele[19][23] != ele[19][27];
    ele[19][23] != ele[19][28];
    ele[19][23] != ele[19][29];
    ele[19][23] != ele[19][30];
    ele[19][23] != ele[19][31];
    ele[19][23] != ele[19][32];
    ele[19][23] != ele[19][33];
    ele[19][23] != ele[19][34];
    ele[19][23] != ele[19][35];
    ele[19][23] != ele[20][18];
    ele[19][23] != ele[20][19];
    ele[19][23] != ele[20][20];
    ele[19][23] != ele[20][21];
    ele[19][23] != ele[20][22];
    ele[19][23] != ele[20][23];
    ele[19][23] != ele[21][18];
    ele[19][23] != ele[21][19];
    ele[19][23] != ele[21][20];
    ele[19][23] != ele[21][21];
    ele[19][23] != ele[21][22];
    ele[19][23] != ele[21][23];
    ele[19][23] != ele[22][18];
    ele[19][23] != ele[22][19];
    ele[19][23] != ele[22][20];
    ele[19][23] != ele[22][21];
    ele[19][23] != ele[22][22];
    ele[19][23] != ele[22][23];
    ele[19][23] != ele[23][18];
    ele[19][23] != ele[23][19];
    ele[19][23] != ele[23][20];
    ele[19][23] != ele[23][21];
    ele[19][23] != ele[23][22];
    ele[19][23] != ele[23][23];
    ele[19][23] != ele[24][23];
    ele[19][23] != ele[25][23];
    ele[19][23] != ele[26][23];
    ele[19][23] != ele[27][23];
    ele[19][23] != ele[28][23];
    ele[19][23] != ele[29][23];
    ele[19][23] != ele[30][23];
    ele[19][23] != ele[31][23];
    ele[19][23] != ele[32][23];
    ele[19][23] != ele[33][23];
    ele[19][23] != ele[34][23];
    ele[19][23] != ele[35][23];
    ele[19][24] != ele[19][25];
    ele[19][24] != ele[19][26];
    ele[19][24] != ele[19][27];
    ele[19][24] != ele[19][28];
    ele[19][24] != ele[19][29];
    ele[19][24] != ele[19][30];
    ele[19][24] != ele[19][31];
    ele[19][24] != ele[19][32];
    ele[19][24] != ele[19][33];
    ele[19][24] != ele[19][34];
    ele[19][24] != ele[19][35];
    ele[19][24] != ele[20][24];
    ele[19][24] != ele[20][25];
    ele[19][24] != ele[20][26];
    ele[19][24] != ele[20][27];
    ele[19][24] != ele[20][28];
    ele[19][24] != ele[20][29];
    ele[19][24] != ele[21][24];
    ele[19][24] != ele[21][25];
    ele[19][24] != ele[21][26];
    ele[19][24] != ele[21][27];
    ele[19][24] != ele[21][28];
    ele[19][24] != ele[21][29];
    ele[19][24] != ele[22][24];
    ele[19][24] != ele[22][25];
    ele[19][24] != ele[22][26];
    ele[19][24] != ele[22][27];
    ele[19][24] != ele[22][28];
    ele[19][24] != ele[22][29];
    ele[19][24] != ele[23][24];
    ele[19][24] != ele[23][25];
    ele[19][24] != ele[23][26];
    ele[19][24] != ele[23][27];
    ele[19][24] != ele[23][28];
    ele[19][24] != ele[23][29];
    ele[19][24] != ele[24][24];
    ele[19][24] != ele[25][24];
    ele[19][24] != ele[26][24];
    ele[19][24] != ele[27][24];
    ele[19][24] != ele[28][24];
    ele[19][24] != ele[29][24];
    ele[19][24] != ele[30][24];
    ele[19][24] != ele[31][24];
    ele[19][24] != ele[32][24];
    ele[19][24] != ele[33][24];
    ele[19][24] != ele[34][24];
    ele[19][24] != ele[35][24];
    ele[19][25] != ele[19][26];
    ele[19][25] != ele[19][27];
    ele[19][25] != ele[19][28];
    ele[19][25] != ele[19][29];
    ele[19][25] != ele[19][30];
    ele[19][25] != ele[19][31];
    ele[19][25] != ele[19][32];
    ele[19][25] != ele[19][33];
    ele[19][25] != ele[19][34];
    ele[19][25] != ele[19][35];
    ele[19][25] != ele[20][24];
    ele[19][25] != ele[20][25];
    ele[19][25] != ele[20][26];
    ele[19][25] != ele[20][27];
    ele[19][25] != ele[20][28];
    ele[19][25] != ele[20][29];
    ele[19][25] != ele[21][24];
    ele[19][25] != ele[21][25];
    ele[19][25] != ele[21][26];
    ele[19][25] != ele[21][27];
    ele[19][25] != ele[21][28];
    ele[19][25] != ele[21][29];
    ele[19][25] != ele[22][24];
    ele[19][25] != ele[22][25];
    ele[19][25] != ele[22][26];
    ele[19][25] != ele[22][27];
    ele[19][25] != ele[22][28];
    ele[19][25] != ele[22][29];
    ele[19][25] != ele[23][24];
    ele[19][25] != ele[23][25];
    ele[19][25] != ele[23][26];
    ele[19][25] != ele[23][27];
    ele[19][25] != ele[23][28];
    ele[19][25] != ele[23][29];
    ele[19][25] != ele[24][25];
    ele[19][25] != ele[25][25];
    ele[19][25] != ele[26][25];
    ele[19][25] != ele[27][25];
    ele[19][25] != ele[28][25];
    ele[19][25] != ele[29][25];
    ele[19][25] != ele[30][25];
    ele[19][25] != ele[31][25];
    ele[19][25] != ele[32][25];
    ele[19][25] != ele[33][25];
    ele[19][25] != ele[34][25];
    ele[19][25] != ele[35][25];
    ele[19][26] != ele[19][27];
    ele[19][26] != ele[19][28];
    ele[19][26] != ele[19][29];
    ele[19][26] != ele[19][30];
    ele[19][26] != ele[19][31];
    ele[19][26] != ele[19][32];
    ele[19][26] != ele[19][33];
    ele[19][26] != ele[19][34];
    ele[19][26] != ele[19][35];
    ele[19][26] != ele[20][24];
    ele[19][26] != ele[20][25];
    ele[19][26] != ele[20][26];
    ele[19][26] != ele[20][27];
    ele[19][26] != ele[20][28];
    ele[19][26] != ele[20][29];
    ele[19][26] != ele[21][24];
    ele[19][26] != ele[21][25];
    ele[19][26] != ele[21][26];
    ele[19][26] != ele[21][27];
    ele[19][26] != ele[21][28];
    ele[19][26] != ele[21][29];
    ele[19][26] != ele[22][24];
    ele[19][26] != ele[22][25];
    ele[19][26] != ele[22][26];
    ele[19][26] != ele[22][27];
    ele[19][26] != ele[22][28];
    ele[19][26] != ele[22][29];
    ele[19][26] != ele[23][24];
    ele[19][26] != ele[23][25];
    ele[19][26] != ele[23][26];
    ele[19][26] != ele[23][27];
    ele[19][26] != ele[23][28];
    ele[19][26] != ele[23][29];
    ele[19][26] != ele[24][26];
    ele[19][26] != ele[25][26];
    ele[19][26] != ele[26][26];
    ele[19][26] != ele[27][26];
    ele[19][26] != ele[28][26];
    ele[19][26] != ele[29][26];
    ele[19][26] != ele[30][26];
    ele[19][26] != ele[31][26];
    ele[19][26] != ele[32][26];
    ele[19][26] != ele[33][26];
    ele[19][26] != ele[34][26];
    ele[19][26] != ele[35][26];
    ele[19][27] != ele[19][28];
    ele[19][27] != ele[19][29];
    ele[19][27] != ele[19][30];
    ele[19][27] != ele[19][31];
    ele[19][27] != ele[19][32];
    ele[19][27] != ele[19][33];
    ele[19][27] != ele[19][34];
    ele[19][27] != ele[19][35];
    ele[19][27] != ele[20][24];
    ele[19][27] != ele[20][25];
    ele[19][27] != ele[20][26];
    ele[19][27] != ele[20][27];
    ele[19][27] != ele[20][28];
    ele[19][27] != ele[20][29];
    ele[19][27] != ele[21][24];
    ele[19][27] != ele[21][25];
    ele[19][27] != ele[21][26];
    ele[19][27] != ele[21][27];
    ele[19][27] != ele[21][28];
    ele[19][27] != ele[21][29];
    ele[19][27] != ele[22][24];
    ele[19][27] != ele[22][25];
    ele[19][27] != ele[22][26];
    ele[19][27] != ele[22][27];
    ele[19][27] != ele[22][28];
    ele[19][27] != ele[22][29];
    ele[19][27] != ele[23][24];
    ele[19][27] != ele[23][25];
    ele[19][27] != ele[23][26];
    ele[19][27] != ele[23][27];
    ele[19][27] != ele[23][28];
    ele[19][27] != ele[23][29];
    ele[19][27] != ele[24][27];
    ele[19][27] != ele[25][27];
    ele[19][27] != ele[26][27];
    ele[19][27] != ele[27][27];
    ele[19][27] != ele[28][27];
    ele[19][27] != ele[29][27];
    ele[19][27] != ele[30][27];
    ele[19][27] != ele[31][27];
    ele[19][27] != ele[32][27];
    ele[19][27] != ele[33][27];
    ele[19][27] != ele[34][27];
    ele[19][27] != ele[35][27];
    ele[19][28] != ele[19][29];
    ele[19][28] != ele[19][30];
    ele[19][28] != ele[19][31];
    ele[19][28] != ele[19][32];
    ele[19][28] != ele[19][33];
    ele[19][28] != ele[19][34];
    ele[19][28] != ele[19][35];
    ele[19][28] != ele[20][24];
    ele[19][28] != ele[20][25];
    ele[19][28] != ele[20][26];
    ele[19][28] != ele[20][27];
    ele[19][28] != ele[20][28];
    ele[19][28] != ele[20][29];
    ele[19][28] != ele[21][24];
    ele[19][28] != ele[21][25];
    ele[19][28] != ele[21][26];
    ele[19][28] != ele[21][27];
    ele[19][28] != ele[21][28];
    ele[19][28] != ele[21][29];
    ele[19][28] != ele[22][24];
    ele[19][28] != ele[22][25];
    ele[19][28] != ele[22][26];
    ele[19][28] != ele[22][27];
    ele[19][28] != ele[22][28];
    ele[19][28] != ele[22][29];
    ele[19][28] != ele[23][24];
    ele[19][28] != ele[23][25];
    ele[19][28] != ele[23][26];
    ele[19][28] != ele[23][27];
    ele[19][28] != ele[23][28];
    ele[19][28] != ele[23][29];
    ele[19][28] != ele[24][28];
    ele[19][28] != ele[25][28];
    ele[19][28] != ele[26][28];
    ele[19][28] != ele[27][28];
    ele[19][28] != ele[28][28];
    ele[19][28] != ele[29][28];
    ele[19][28] != ele[30][28];
    ele[19][28] != ele[31][28];
    ele[19][28] != ele[32][28];
    ele[19][28] != ele[33][28];
    ele[19][28] != ele[34][28];
    ele[19][28] != ele[35][28];
    ele[19][29] != ele[19][30];
    ele[19][29] != ele[19][31];
    ele[19][29] != ele[19][32];
    ele[19][29] != ele[19][33];
    ele[19][29] != ele[19][34];
    ele[19][29] != ele[19][35];
    ele[19][29] != ele[20][24];
    ele[19][29] != ele[20][25];
    ele[19][29] != ele[20][26];
    ele[19][29] != ele[20][27];
    ele[19][29] != ele[20][28];
    ele[19][29] != ele[20][29];
    ele[19][29] != ele[21][24];
    ele[19][29] != ele[21][25];
    ele[19][29] != ele[21][26];
    ele[19][29] != ele[21][27];
    ele[19][29] != ele[21][28];
    ele[19][29] != ele[21][29];
    ele[19][29] != ele[22][24];
    ele[19][29] != ele[22][25];
    ele[19][29] != ele[22][26];
    ele[19][29] != ele[22][27];
    ele[19][29] != ele[22][28];
    ele[19][29] != ele[22][29];
    ele[19][29] != ele[23][24];
    ele[19][29] != ele[23][25];
    ele[19][29] != ele[23][26];
    ele[19][29] != ele[23][27];
    ele[19][29] != ele[23][28];
    ele[19][29] != ele[23][29];
    ele[19][29] != ele[24][29];
    ele[19][29] != ele[25][29];
    ele[19][29] != ele[26][29];
    ele[19][29] != ele[27][29];
    ele[19][29] != ele[28][29];
    ele[19][29] != ele[29][29];
    ele[19][29] != ele[30][29];
    ele[19][29] != ele[31][29];
    ele[19][29] != ele[32][29];
    ele[19][29] != ele[33][29];
    ele[19][29] != ele[34][29];
    ele[19][29] != ele[35][29];
    ele[19][3] != ele[19][10];
    ele[19][3] != ele[19][11];
    ele[19][3] != ele[19][12];
    ele[19][3] != ele[19][13];
    ele[19][3] != ele[19][14];
    ele[19][3] != ele[19][15];
    ele[19][3] != ele[19][16];
    ele[19][3] != ele[19][17];
    ele[19][3] != ele[19][18];
    ele[19][3] != ele[19][19];
    ele[19][3] != ele[19][20];
    ele[19][3] != ele[19][21];
    ele[19][3] != ele[19][22];
    ele[19][3] != ele[19][23];
    ele[19][3] != ele[19][24];
    ele[19][3] != ele[19][25];
    ele[19][3] != ele[19][26];
    ele[19][3] != ele[19][27];
    ele[19][3] != ele[19][28];
    ele[19][3] != ele[19][29];
    ele[19][3] != ele[19][30];
    ele[19][3] != ele[19][31];
    ele[19][3] != ele[19][32];
    ele[19][3] != ele[19][33];
    ele[19][3] != ele[19][34];
    ele[19][3] != ele[19][35];
    ele[19][3] != ele[19][4];
    ele[19][3] != ele[19][5];
    ele[19][3] != ele[19][6];
    ele[19][3] != ele[19][7];
    ele[19][3] != ele[19][8];
    ele[19][3] != ele[19][9];
    ele[19][3] != ele[20][0];
    ele[19][3] != ele[20][1];
    ele[19][3] != ele[20][2];
    ele[19][3] != ele[20][3];
    ele[19][3] != ele[20][4];
    ele[19][3] != ele[20][5];
    ele[19][3] != ele[21][0];
    ele[19][3] != ele[21][1];
    ele[19][3] != ele[21][2];
    ele[19][3] != ele[21][3];
    ele[19][3] != ele[21][4];
    ele[19][3] != ele[21][5];
    ele[19][3] != ele[22][0];
    ele[19][3] != ele[22][1];
    ele[19][3] != ele[22][2];
    ele[19][3] != ele[22][3];
    ele[19][3] != ele[22][4];
    ele[19][3] != ele[22][5];
    ele[19][3] != ele[23][0];
    ele[19][3] != ele[23][1];
    ele[19][3] != ele[23][2];
    ele[19][3] != ele[23][3];
    ele[19][3] != ele[23][4];
    ele[19][3] != ele[23][5];
    ele[19][3] != ele[24][3];
    ele[19][3] != ele[25][3];
    ele[19][3] != ele[26][3];
    ele[19][3] != ele[27][3];
    ele[19][3] != ele[28][3];
    ele[19][3] != ele[29][3];
    ele[19][3] != ele[30][3];
    ele[19][3] != ele[31][3];
    ele[19][3] != ele[32][3];
    ele[19][3] != ele[33][3];
    ele[19][3] != ele[34][3];
    ele[19][3] != ele[35][3];
    ele[19][30] != ele[19][31];
    ele[19][30] != ele[19][32];
    ele[19][30] != ele[19][33];
    ele[19][30] != ele[19][34];
    ele[19][30] != ele[19][35];
    ele[19][30] != ele[20][30];
    ele[19][30] != ele[20][31];
    ele[19][30] != ele[20][32];
    ele[19][30] != ele[20][33];
    ele[19][30] != ele[20][34];
    ele[19][30] != ele[20][35];
    ele[19][30] != ele[21][30];
    ele[19][30] != ele[21][31];
    ele[19][30] != ele[21][32];
    ele[19][30] != ele[21][33];
    ele[19][30] != ele[21][34];
    ele[19][30] != ele[21][35];
    ele[19][30] != ele[22][30];
    ele[19][30] != ele[22][31];
    ele[19][30] != ele[22][32];
    ele[19][30] != ele[22][33];
    ele[19][30] != ele[22][34];
    ele[19][30] != ele[22][35];
    ele[19][30] != ele[23][30];
    ele[19][30] != ele[23][31];
    ele[19][30] != ele[23][32];
    ele[19][30] != ele[23][33];
    ele[19][30] != ele[23][34];
    ele[19][30] != ele[23][35];
    ele[19][30] != ele[24][30];
    ele[19][30] != ele[25][30];
    ele[19][30] != ele[26][30];
    ele[19][30] != ele[27][30];
    ele[19][30] != ele[28][30];
    ele[19][30] != ele[29][30];
    ele[19][30] != ele[30][30];
    ele[19][30] != ele[31][30];
    ele[19][30] != ele[32][30];
    ele[19][30] != ele[33][30];
    ele[19][30] != ele[34][30];
    ele[19][30] != ele[35][30];
    ele[19][31] != ele[19][32];
    ele[19][31] != ele[19][33];
    ele[19][31] != ele[19][34];
    ele[19][31] != ele[19][35];
    ele[19][31] != ele[20][30];
    ele[19][31] != ele[20][31];
    ele[19][31] != ele[20][32];
    ele[19][31] != ele[20][33];
    ele[19][31] != ele[20][34];
    ele[19][31] != ele[20][35];
    ele[19][31] != ele[21][30];
    ele[19][31] != ele[21][31];
    ele[19][31] != ele[21][32];
    ele[19][31] != ele[21][33];
    ele[19][31] != ele[21][34];
    ele[19][31] != ele[21][35];
    ele[19][31] != ele[22][30];
    ele[19][31] != ele[22][31];
    ele[19][31] != ele[22][32];
    ele[19][31] != ele[22][33];
    ele[19][31] != ele[22][34];
    ele[19][31] != ele[22][35];
    ele[19][31] != ele[23][30];
    ele[19][31] != ele[23][31];
    ele[19][31] != ele[23][32];
    ele[19][31] != ele[23][33];
    ele[19][31] != ele[23][34];
    ele[19][31] != ele[23][35];
    ele[19][31] != ele[24][31];
    ele[19][31] != ele[25][31];
    ele[19][31] != ele[26][31];
    ele[19][31] != ele[27][31];
    ele[19][31] != ele[28][31];
    ele[19][31] != ele[29][31];
    ele[19][31] != ele[30][31];
    ele[19][31] != ele[31][31];
    ele[19][31] != ele[32][31];
    ele[19][31] != ele[33][31];
    ele[19][31] != ele[34][31];
    ele[19][31] != ele[35][31];
    ele[19][32] != ele[19][33];
    ele[19][32] != ele[19][34];
    ele[19][32] != ele[19][35];
    ele[19][32] != ele[20][30];
    ele[19][32] != ele[20][31];
    ele[19][32] != ele[20][32];
    ele[19][32] != ele[20][33];
    ele[19][32] != ele[20][34];
    ele[19][32] != ele[20][35];
    ele[19][32] != ele[21][30];
    ele[19][32] != ele[21][31];
    ele[19][32] != ele[21][32];
    ele[19][32] != ele[21][33];
    ele[19][32] != ele[21][34];
    ele[19][32] != ele[21][35];
    ele[19][32] != ele[22][30];
    ele[19][32] != ele[22][31];
    ele[19][32] != ele[22][32];
    ele[19][32] != ele[22][33];
    ele[19][32] != ele[22][34];
    ele[19][32] != ele[22][35];
    ele[19][32] != ele[23][30];
    ele[19][32] != ele[23][31];
    ele[19][32] != ele[23][32];
    ele[19][32] != ele[23][33];
    ele[19][32] != ele[23][34];
    ele[19][32] != ele[23][35];
    ele[19][32] != ele[24][32];
    ele[19][32] != ele[25][32];
    ele[19][32] != ele[26][32];
    ele[19][32] != ele[27][32];
    ele[19][32] != ele[28][32];
    ele[19][32] != ele[29][32];
    ele[19][32] != ele[30][32];
    ele[19][32] != ele[31][32];
    ele[19][32] != ele[32][32];
    ele[19][32] != ele[33][32];
    ele[19][32] != ele[34][32];
    ele[19][32] != ele[35][32];
    ele[19][33] != ele[19][34];
    ele[19][33] != ele[19][35];
    ele[19][33] != ele[20][30];
    ele[19][33] != ele[20][31];
    ele[19][33] != ele[20][32];
    ele[19][33] != ele[20][33];
    ele[19][33] != ele[20][34];
    ele[19][33] != ele[20][35];
    ele[19][33] != ele[21][30];
    ele[19][33] != ele[21][31];
    ele[19][33] != ele[21][32];
    ele[19][33] != ele[21][33];
    ele[19][33] != ele[21][34];
    ele[19][33] != ele[21][35];
    ele[19][33] != ele[22][30];
    ele[19][33] != ele[22][31];
    ele[19][33] != ele[22][32];
    ele[19][33] != ele[22][33];
    ele[19][33] != ele[22][34];
    ele[19][33] != ele[22][35];
    ele[19][33] != ele[23][30];
    ele[19][33] != ele[23][31];
    ele[19][33] != ele[23][32];
    ele[19][33] != ele[23][33];
    ele[19][33] != ele[23][34];
    ele[19][33] != ele[23][35];
    ele[19][33] != ele[24][33];
    ele[19][33] != ele[25][33];
    ele[19][33] != ele[26][33];
    ele[19][33] != ele[27][33];
    ele[19][33] != ele[28][33];
    ele[19][33] != ele[29][33];
    ele[19][33] != ele[30][33];
    ele[19][33] != ele[31][33];
    ele[19][33] != ele[32][33];
    ele[19][33] != ele[33][33];
    ele[19][33] != ele[34][33];
    ele[19][33] != ele[35][33];
    ele[19][34] != ele[19][35];
    ele[19][34] != ele[20][30];
    ele[19][34] != ele[20][31];
    ele[19][34] != ele[20][32];
    ele[19][34] != ele[20][33];
    ele[19][34] != ele[20][34];
    ele[19][34] != ele[20][35];
    ele[19][34] != ele[21][30];
    ele[19][34] != ele[21][31];
    ele[19][34] != ele[21][32];
    ele[19][34] != ele[21][33];
    ele[19][34] != ele[21][34];
    ele[19][34] != ele[21][35];
    ele[19][34] != ele[22][30];
    ele[19][34] != ele[22][31];
    ele[19][34] != ele[22][32];
    ele[19][34] != ele[22][33];
    ele[19][34] != ele[22][34];
    ele[19][34] != ele[22][35];
    ele[19][34] != ele[23][30];
    ele[19][34] != ele[23][31];
    ele[19][34] != ele[23][32];
    ele[19][34] != ele[23][33];
    ele[19][34] != ele[23][34];
    ele[19][34] != ele[23][35];
    ele[19][34] != ele[24][34];
    ele[19][34] != ele[25][34];
    ele[19][34] != ele[26][34];
    ele[19][34] != ele[27][34];
    ele[19][34] != ele[28][34];
    ele[19][34] != ele[29][34];
    ele[19][34] != ele[30][34];
    ele[19][34] != ele[31][34];
    ele[19][34] != ele[32][34];
    ele[19][34] != ele[33][34];
    ele[19][34] != ele[34][34];
    ele[19][34] != ele[35][34];
    ele[19][35] != ele[20][30];
    ele[19][35] != ele[20][31];
    ele[19][35] != ele[20][32];
    ele[19][35] != ele[20][33];
    ele[19][35] != ele[20][34];
    ele[19][35] != ele[20][35];
    ele[19][35] != ele[21][30];
    ele[19][35] != ele[21][31];
    ele[19][35] != ele[21][32];
    ele[19][35] != ele[21][33];
    ele[19][35] != ele[21][34];
    ele[19][35] != ele[21][35];
    ele[19][35] != ele[22][30];
    ele[19][35] != ele[22][31];
    ele[19][35] != ele[22][32];
    ele[19][35] != ele[22][33];
    ele[19][35] != ele[22][34];
    ele[19][35] != ele[22][35];
    ele[19][35] != ele[23][30];
    ele[19][35] != ele[23][31];
    ele[19][35] != ele[23][32];
    ele[19][35] != ele[23][33];
    ele[19][35] != ele[23][34];
    ele[19][35] != ele[23][35];
    ele[19][35] != ele[24][35];
    ele[19][35] != ele[25][35];
    ele[19][35] != ele[26][35];
    ele[19][35] != ele[27][35];
    ele[19][35] != ele[28][35];
    ele[19][35] != ele[29][35];
    ele[19][35] != ele[30][35];
    ele[19][35] != ele[31][35];
    ele[19][35] != ele[32][35];
    ele[19][35] != ele[33][35];
    ele[19][35] != ele[34][35];
    ele[19][35] != ele[35][35];
    ele[19][4] != ele[19][10];
    ele[19][4] != ele[19][11];
    ele[19][4] != ele[19][12];
    ele[19][4] != ele[19][13];
    ele[19][4] != ele[19][14];
    ele[19][4] != ele[19][15];
    ele[19][4] != ele[19][16];
    ele[19][4] != ele[19][17];
    ele[19][4] != ele[19][18];
    ele[19][4] != ele[19][19];
    ele[19][4] != ele[19][20];
    ele[19][4] != ele[19][21];
    ele[19][4] != ele[19][22];
    ele[19][4] != ele[19][23];
    ele[19][4] != ele[19][24];
    ele[19][4] != ele[19][25];
    ele[19][4] != ele[19][26];
    ele[19][4] != ele[19][27];
    ele[19][4] != ele[19][28];
    ele[19][4] != ele[19][29];
    ele[19][4] != ele[19][30];
    ele[19][4] != ele[19][31];
    ele[19][4] != ele[19][32];
    ele[19][4] != ele[19][33];
    ele[19][4] != ele[19][34];
    ele[19][4] != ele[19][35];
    ele[19][4] != ele[19][5];
    ele[19][4] != ele[19][6];
    ele[19][4] != ele[19][7];
    ele[19][4] != ele[19][8];
    ele[19][4] != ele[19][9];
    ele[19][4] != ele[20][0];
    ele[19][4] != ele[20][1];
    ele[19][4] != ele[20][2];
    ele[19][4] != ele[20][3];
    ele[19][4] != ele[20][4];
    ele[19][4] != ele[20][5];
    ele[19][4] != ele[21][0];
    ele[19][4] != ele[21][1];
    ele[19][4] != ele[21][2];
    ele[19][4] != ele[21][3];
    ele[19][4] != ele[21][4];
    ele[19][4] != ele[21][5];
    ele[19][4] != ele[22][0];
    ele[19][4] != ele[22][1];
    ele[19][4] != ele[22][2];
    ele[19][4] != ele[22][3];
    ele[19][4] != ele[22][4];
    ele[19][4] != ele[22][5];
    ele[19][4] != ele[23][0];
    ele[19][4] != ele[23][1];
    ele[19][4] != ele[23][2];
    ele[19][4] != ele[23][3];
    ele[19][4] != ele[23][4];
    ele[19][4] != ele[23][5];
    ele[19][4] != ele[24][4];
    ele[19][4] != ele[25][4];
    ele[19][4] != ele[26][4];
    ele[19][4] != ele[27][4];
    ele[19][4] != ele[28][4];
    ele[19][4] != ele[29][4];
    ele[19][4] != ele[30][4];
    ele[19][4] != ele[31][4];
    ele[19][4] != ele[32][4];
    ele[19][4] != ele[33][4];
    ele[19][4] != ele[34][4];
    ele[19][4] != ele[35][4];
    ele[19][5] != ele[19][10];
    ele[19][5] != ele[19][11];
    ele[19][5] != ele[19][12];
    ele[19][5] != ele[19][13];
    ele[19][5] != ele[19][14];
    ele[19][5] != ele[19][15];
    ele[19][5] != ele[19][16];
    ele[19][5] != ele[19][17];
    ele[19][5] != ele[19][18];
    ele[19][5] != ele[19][19];
    ele[19][5] != ele[19][20];
    ele[19][5] != ele[19][21];
    ele[19][5] != ele[19][22];
    ele[19][5] != ele[19][23];
    ele[19][5] != ele[19][24];
    ele[19][5] != ele[19][25];
    ele[19][5] != ele[19][26];
    ele[19][5] != ele[19][27];
    ele[19][5] != ele[19][28];
    ele[19][5] != ele[19][29];
    ele[19][5] != ele[19][30];
    ele[19][5] != ele[19][31];
    ele[19][5] != ele[19][32];
    ele[19][5] != ele[19][33];
    ele[19][5] != ele[19][34];
    ele[19][5] != ele[19][35];
    ele[19][5] != ele[19][6];
    ele[19][5] != ele[19][7];
    ele[19][5] != ele[19][8];
    ele[19][5] != ele[19][9];
    ele[19][5] != ele[20][0];
    ele[19][5] != ele[20][1];
    ele[19][5] != ele[20][2];
    ele[19][5] != ele[20][3];
    ele[19][5] != ele[20][4];
    ele[19][5] != ele[20][5];
    ele[19][5] != ele[21][0];
    ele[19][5] != ele[21][1];
    ele[19][5] != ele[21][2];
    ele[19][5] != ele[21][3];
    ele[19][5] != ele[21][4];
    ele[19][5] != ele[21][5];
    ele[19][5] != ele[22][0];
    ele[19][5] != ele[22][1];
    ele[19][5] != ele[22][2];
    ele[19][5] != ele[22][3];
    ele[19][5] != ele[22][4];
    ele[19][5] != ele[22][5];
    ele[19][5] != ele[23][0];
    ele[19][5] != ele[23][1];
    ele[19][5] != ele[23][2];
    ele[19][5] != ele[23][3];
    ele[19][5] != ele[23][4];
    ele[19][5] != ele[23][5];
    ele[19][5] != ele[24][5];
    ele[19][5] != ele[25][5];
    ele[19][5] != ele[26][5];
    ele[19][5] != ele[27][5];
    ele[19][5] != ele[28][5];
    ele[19][5] != ele[29][5];
    ele[19][5] != ele[30][5];
    ele[19][5] != ele[31][5];
    ele[19][5] != ele[32][5];
    ele[19][5] != ele[33][5];
    ele[19][5] != ele[34][5];
    ele[19][5] != ele[35][5];
    ele[19][6] != ele[19][10];
    ele[19][6] != ele[19][11];
    ele[19][6] != ele[19][12];
    ele[19][6] != ele[19][13];
    ele[19][6] != ele[19][14];
    ele[19][6] != ele[19][15];
    ele[19][6] != ele[19][16];
    ele[19][6] != ele[19][17];
    ele[19][6] != ele[19][18];
    ele[19][6] != ele[19][19];
    ele[19][6] != ele[19][20];
    ele[19][6] != ele[19][21];
    ele[19][6] != ele[19][22];
    ele[19][6] != ele[19][23];
    ele[19][6] != ele[19][24];
    ele[19][6] != ele[19][25];
    ele[19][6] != ele[19][26];
    ele[19][6] != ele[19][27];
    ele[19][6] != ele[19][28];
    ele[19][6] != ele[19][29];
    ele[19][6] != ele[19][30];
    ele[19][6] != ele[19][31];
    ele[19][6] != ele[19][32];
    ele[19][6] != ele[19][33];
    ele[19][6] != ele[19][34];
    ele[19][6] != ele[19][35];
    ele[19][6] != ele[19][7];
    ele[19][6] != ele[19][8];
    ele[19][6] != ele[19][9];
    ele[19][6] != ele[20][10];
    ele[19][6] != ele[20][11];
    ele[19][6] != ele[20][6];
    ele[19][6] != ele[20][7];
    ele[19][6] != ele[20][8];
    ele[19][6] != ele[20][9];
    ele[19][6] != ele[21][10];
    ele[19][6] != ele[21][11];
    ele[19][6] != ele[21][6];
    ele[19][6] != ele[21][7];
    ele[19][6] != ele[21][8];
    ele[19][6] != ele[21][9];
    ele[19][6] != ele[22][10];
    ele[19][6] != ele[22][11];
    ele[19][6] != ele[22][6];
    ele[19][6] != ele[22][7];
    ele[19][6] != ele[22][8];
    ele[19][6] != ele[22][9];
    ele[19][6] != ele[23][10];
    ele[19][6] != ele[23][11];
    ele[19][6] != ele[23][6];
    ele[19][6] != ele[23][7];
    ele[19][6] != ele[23][8];
    ele[19][6] != ele[23][9];
    ele[19][6] != ele[24][6];
    ele[19][6] != ele[25][6];
    ele[19][6] != ele[26][6];
    ele[19][6] != ele[27][6];
    ele[19][6] != ele[28][6];
    ele[19][6] != ele[29][6];
    ele[19][6] != ele[30][6];
    ele[19][6] != ele[31][6];
    ele[19][6] != ele[32][6];
    ele[19][6] != ele[33][6];
    ele[19][6] != ele[34][6];
    ele[19][6] != ele[35][6];
    ele[19][7] != ele[19][10];
    ele[19][7] != ele[19][11];
    ele[19][7] != ele[19][12];
    ele[19][7] != ele[19][13];
    ele[19][7] != ele[19][14];
    ele[19][7] != ele[19][15];
    ele[19][7] != ele[19][16];
    ele[19][7] != ele[19][17];
    ele[19][7] != ele[19][18];
    ele[19][7] != ele[19][19];
    ele[19][7] != ele[19][20];
    ele[19][7] != ele[19][21];
    ele[19][7] != ele[19][22];
    ele[19][7] != ele[19][23];
    ele[19][7] != ele[19][24];
    ele[19][7] != ele[19][25];
    ele[19][7] != ele[19][26];
    ele[19][7] != ele[19][27];
    ele[19][7] != ele[19][28];
    ele[19][7] != ele[19][29];
    ele[19][7] != ele[19][30];
    ele[19][7] != ele[19][31];
    ele[19][7] != ele[19][32];
    ele[19][7] != ele[19][33];
    ele[19][7] != ele[19][34];
    ele[19][7] != ele[19][35];
    ele[19][7] != ele[19][8];
    ele[19][7] != ele[19][9];
    ele[19][7] != ele[20][10];
    ele[19][7] != ele[20][11];
    ele[19][7] != ele[20][6];
    ele[19][7] != ele[20][7];
    ele[19][7] != ele[20][8];
    ele[19][7] != ele[20][9];
    ele[19][7] != ele[21][10];
    ele[19][7] != ele[21][11];
    ele[19][7] != ele[21][6];
    ele[19][7] != ele[21][7];
    ele[19][7] != ele[21][8];
    ele[19][7] != ele[21][9];
    ele[19][7] != ele[22][10];
    ele[19][7] != ele[22][11];
    ele[19][7] != ele[22][6];
    ele[19][7] != ele[22][7];
    ele[19][7] != ele[22][8];
    ele[19][7] != ele[22][9];
    ele[19][7] != ele[23][10];
    ele[19][7] != ele[23][11];
    ele[19][7] != ele[23][6];
    ele[19][7] != ele[23][7];
    ele[19][7] != ele[23][8];
    ele[19][7] != ele[23][9];
    ele[19][7] != ele[24][7];
    ele[19][7] != ele[25][7];
    ele[19][7] != ele[26][7];
    ele[19][7] != ele[27][7];
    ele[19][7] != ele[28][7];
    ele[19][7] != ele[29][7];
    ele[19][7] != ele[30][7];
    ele[19][7] != ele[31][7];
    ele[19][7] != ele[32][7];
    ele[19][7] != ele[33][7];
    ele[19][7] != ele[34][7];
    ele[19][7] != ele[35][7];
    ele[19][8] != ele[19][10];
    ele[19][8] != ele[19][11];
    ele[19][8] != ele[19][12];
    ele[19][8] != ele[19][13];
    ele[19][8] != ele[19][14];
    ele[19][8] != ele[19][15];
    ele[19][8] != ele[19][16];
    ele[19][8] != ele[19][17];
    ele[19][8] != ele[19][18];
    ele[19][8] != ele[19][19];
    ele[19][8] != ele[19][20];
    ele[19][8] != ele[19][21];
    ele[19][8] != ele[19][22];
    ele[19][8] != ele[19][23];
    ele[19][8] != ele[19][24];
    ele[19][8] != ele[19][25];
    ele[19][8] != ele[19][26];
    ele[19][8] != ele[19][27];
    ele[19][8] != ele[19][28];
    ele[19][8] != ele[19][29];
    ele[19][8] != ele[19][30];
    ele[19][8] != ele[19][31];
    ele[19][8] != ele[19][32];
    ele[19][8] != ele[19][33];
    ele[19][8] != ele[19][34];
    ele[19][8] != ele[19][35];
    ele[19][8] != ele[19][9];
    ele[19][8] != ele[20][10];
    ele[19][8] != ele[20][11];
    ele[19][8] != ele[20][6];
    ele[19][8] != ele[20][7];
    ele[19][8] != ele[20][8];
    ele[19][8] != ele[20][9];
    ele[19][8] != ele[21][10];
    ele[19][8] != ele[21][11];
    ele[19][8] != ele[21][6];
    ele[19][8] != ele[21][7];
    ele[19][8] != ele[21][8];
    ele[19][8] != ele[21][9];
    ele[19][8] != ele[22][10];
    ele[19][8] != ele[22][11];
    ele[19][8] != ele[22][6];
    ele[19][8] != ele[22][7];
    ele[19][8] != ele[22][8];
    ele[19][8] != ele[22][9];
    ele[19][8] != ele[23][10];
    ele[19][8] != ele[23][11];
    ele[19][8] != ele[23][6];
    ele[19][8] != ele[23][7];
    ele[19][8] != ele[23][8];
    ele[19][8] != ele[23][9];
    ele[19][8] != ele[24][8];
    ele[19][8] != ele[25][8];
    ele[19][8] != ele[26][8];
    ele[19][8] != ele[27][8];
    ele[19][8] != ele[28][8];
    ele[19][8] != ele[29][8];
    ele[19][8] != ele[30][8];
    ele[19][8] != ele[31][8];
    ele[19][8] != ele[32][8];
    ele[19][8] != ele[33][8];
    ele[19][8] != ele[34][8];
    ele[19][8] != ele[35][8];
    ele[19][9] != ele[19][10];
    ele[19][9] != ele[19][11];
    ele[19][9] != ele[19][12];
    ele[19][9] != ele[19][13];
    ele[19][9] != ele[19][14];
    ele[19][9] != ele[19][15];
    ele[19][9] != ele[19][16];
    ele[19][9] != ele[19][17];
    ele[19][9] != ele[19][18];
    ele[19][9] != ele[19][19];
    ele[19][9] != ele[19][20];
    ele[19][9] != ele[19][21];
    ele[19][9] != ele[19][22];
    ele[19][9] != ele[19][23];
    ele[19][9] != ele[19][24];
    ele[19][9] != ele[19][25];
    ele[19][9] != ele[19][26];
    ele[19][9] != ele[19][27];
    ele[19][9] != ele[19][28];
    ele[19][9] != ele[19][29];
    ele[19][9] != ele[19][30];
    ele[19][9] != ele[19][31];
    ele[19][9] != ele[19][32];
    ele[19][9] != ele[19][33];
    ele[19][9] != ele[19][34];
    ele[19][9] != ele[19][35];
    ele[19][9] != ele[20][10];
    ele[19][9] != ele[20][11];
    ele[19][9] != ele[20][6];
    ele[19][9] != ele[20][7];
    ele[19][9] != ele[20][8];
    ele[19][9] != ele[20][9];
    ele[19][9] != ele[21][10];
    ele[19][9] != ele[21][11];
    ele[19][9] != ele[21][6];
    ele[19][9] != ele[21][7];
    ele[19][9] != ele[21][8];
    ele[19][9] != ele[21][9];
    ele[19][9] != ele[22][10];
    ele[19][9] != ele[22][11];
    ele[19][9] != ele[22][6];
    ele[19][9] != ele[22][7];
    ele[19][9] != ele[22][8];
    ele[19][9] != ele[22][9];
    ele[19][9] != ele[23][10];
    ele[19][9] != ele[23][11];
    ele[19][9] != ele[23][6];
    ele[19][9] != ele[23][7];
    ele[19][9] != ele[23][8];
    ele[19][9] != ele[23][9];
    ele[19][9] != ele[24][9];
    ele[19][9] != ele[25][9];
    ele[19][9] != ele[26][9];
    ele[19][9] != ele[27][9];
    ele[19][9] != ele[28][9];
    ele[19][9] != ele[29][9];
    ele[19][9] != ele[30][9];
    ele[19][9] != ele[31][9];
    ele[19][9] != ele[32][9];
    ele[19][9] != ele[33][9];
    ele[19][9] != ele[34][9];
    ele[19][9] != ele[35][9];
    ele[2][0] != ele[10][0];
    ele[2][0] != ele[11][0];
    ele[2][0] != ele[12][0];
    ele[2][0] != ele[13][0];
    ele[2][0] != ele[14][0];
    ele[2][0] != ele[15][0];
    ele[2][0] != ele[16][0];
    ele[2][0] != ele[17][0];
    ele[2][0] != ele[18][0];
    ele[2][0] != ele[19][0];
    ele[2][0] != ele[2][1];
    ele[2][0] != ele[2][10];
    ele[2][0] != ele[2][11];
    ele[2][0] != ele[2][12];
    ele[2][0] != ele[2][13];
    ele[2][0] != ele[2][14];
    ele[2][0] != ele[2][15];
    ele[2][0] != ele[2][16];
    ele[2][0] != ele[2][17];
    ele[2][0] != ele[2][18];
    ele[2][0] != ele[2][19];
    ele[2][0] != ele[2][2];
    ele[2][0] != ele[2][20];
    ele[2][0] != ele[2][21];
    ele[2][0] != ele[2][22];
    ele[2][0] != ele[2][23];
    ele[2][0] != ele[2][24];
    ele[2][0] != ele[2][25];
    ele[2][0] != ele[2][26];
    ele[2][0] != ele[2][27];
    ele[2][0] != ele[2][28];
    ele[2][0] != ele[2][29];
    ele[2][0] != ele[2][3];
    ele[2][0] != ele[2][30];
    ele[2][0] != ele[2][31];
    ele[2][0] != ele[2][32];
    ele[2][0] != ele[2][33];
    ele[2][0] != ele[2][34];
    ele[2][0] != ele[2][35];
    ele[2][0] != ele[2][4];
    ele[2][0] != ele[2][5];
    ele[2][0] != ele[2][6];
    ele[2][0] != ele[2][7];
    ele[2][0] != ele[2][8];
    ele[2][0] != ele[2][9];
    ele[2][0] != ele[20][0];
    ele[2][0] != ele[21][0];
    ele[2][0] != ele[22][0];
    ele[2][0] != ele[23][0];
    ele[2][0] != ele[24][0];
    ele[2][0] != ele[25][0];
    ele[2][0] != ele[26][0];
    ele[2][0] != ele[27][0];
    ele[2][0] != ele[28][0];
    ele[2][0] != ele[29][0];
    ele[2][0] != ele[3][0];
    ele[2][0] != ele[3][1];
    ele[2][0] != ele[3][2];
    ele[2][0] != ele[3][3];
    ele[2][0] != ele[3][4];
    ele[2][0] != ele[3][5];
    ele[2][0] != ele[30][0];
    ele[2][0] != ele[31][0];
    ele[2][0] != ele[32][0];
    ele[2][0] != ele[33][0];
    ele[2][0] != ele[34][0];
    ele[2][0] != ele[35][0];
    ele[2][0] != ele[4][0];
    ele[2][0] != ele[4][1];
    ele[2][0] != ele[4][2];
    ele[2][0] != ele[4][3];
    ele[2][0] != ele[4][4];
    ele[2][0] != ele[4][5];
    ele[2][0] != ele[5][0];
    ele[2][0] != ele[5][1];
    ele[2][0] != ele[5][2];
    ele[2][0] != ele[5][3];
    ele[2][0] != ele[5][4];
    ele[2][0] != ele[5][5];
    ele[2][0] != ele[6][0];
    ele[2][0] != ele[7][0];
    ele[2][0] != ele[8][0];
    ele[2][0] != ele[9][0];
    ele[2][1] != ele[10][1];
    ele[2][1] != ele[11][1];
    ele[2][1] != ele[12][1];
    ele[2][1] != ele[13][1];
    ele[2][1] != ele[14][1];
    ele[2][1] != ele[15][1];
    ele[2][1] != ele[16][1];
    ele[2][1] != ele[17][1];
    ele[2][1] != ele[18][1];
    ele[2][1] != ele[19][1];
    ele[2][1] != ele[2][10];
    ele[2][1] != ele[2][11];
    ele[2][1] != ele[2][12];
    ele[2][1] != ele[2][13];
    ele[2][1] != ele[2][14];
    ele[2][1] != ele[2][15];
    ele[2][1] != ele[2][16];
    ele[2][1] != ele[2][17];
    ele[2][1] != ele[2][18];
    ele[2][1] != ele[2][19];
    ele[2][1] != ele[2][2];
    ele[2][1] != ele[2][20];
    ele[2][1] != ele[2][21];
    ele[2][1] != ele[2][22];
    ele[2][1] != ele[2][23];
    ele[2][1] != ele[2][24];
    ele[2][1] != ele[2][25];
    ele[2][1] != ele[2][26];
    ele[2][1] != ele[2][27];
    ele[2][1] != ele[2][28];
    ele[2][1] != ele[2][29];
    ele[2][1] != ele[2][3];
    ele[2][1] != ele[2][30];
    ele[2][1] != ele[2][31];
    ele[2][1] != ele[2][32];
    ele[2][1] != ele[2][33];
    ele[2][1] != ele[2][34];
    ele[2][1] != ele[2][35];
    ele[2][1] != ele[2][4];
    ele[2][1] != ele[2][5];
    ele[2][1] != ele[2][6];
    ele[2][1] != ele[2][7];
    ele[2][1] != ele[2][8];
    ele[2][1] != ele[2][9];
    ele[2][1] != ele[20][1];
    ele[2][1] != ele[21][1];
    ele[2][1] != ele[22][1];
    ele[2][1] != ele[23][1];
    ele[2][1] != ele[24][1];
    ele[2][1] != ele[25][1];
    ele[2][1] != ele[26][1];
    ele[2][1] != ele[27][1];
    ele[2][1] != ele[28][1];
    ele[2][1] != ele[29][1];
    ele[2][1] != ele[3][0];
    ele[2][1] != ele[3][1];
    ele[2][1] != ele[3][2];
    ele[2][1] != ele[3][3];
    ele[2][1] != ele[3][4];
    ele[2][1] != ele[3][5];
    ele[2][1] != ele[30][1];
    ele[2][1] != ele[31][1];
    ele[2][1] != ele[32][1];
    ele[2][1] != ele[33][1];
    ele[2][1] != ele[34][1];
    ele[2][1] != ele[35][1];
    ele[2][1] != ele[4][0];
    ele[2][1] != ele[4][1];
    ele[2][1] != ele[4][2];
    ele[2][1] != ele[4][3];
    ele[2][1] != ele[4][4];
    ele[2][1] != ele[4][5];
    ele[2][1] != ele[5][0];
    ele[2][1] != ele[5][1];
    ele[2][1] != ele[5][2];
    ele[2][1] != ele[5][3];
    ele[2][1] != ele[5][4];
    ele[2][1] != ele[5][5];
    ele[2][1] != ele[6][1];
    ele[2][1] != ele[7][1];
    ele[2][1] != ele[8][1];
    ele[2][1] != ele[9][1];
    ele[2][10] != ele[10][10];
    ele[2][10] != ele[11][10];
    ele[2][10] != ele[12][10];
    ele[2][10] != ele[13][10];
    ele[2][10] != ele[14][10];
    ele[2][10] != ele[15][10];
    ele[2][10] != ele[16][10];
    ele[2][10] != ele[17][10];
    ele[2][10] != ele[18][10];
    ele[2][10] != ele[19][10];
    ele[2][10] != ele[2][11];
    ele[2][10] != ele[2][12];
    ele[2][10] != ele[2][13];
    ele[2][10] != ele[2][14];
    ele[2][10] != ele[2][15];
    ele[2][10] != ele[2][16];
    ele[2][10] != ele[2][17];
    ele[2][10] != ele[2][18];
    ele[2][10] != ele[2][19];
    ele[2][10] != ele[2][20];
    ele[2][10] != ele[2][21];
    ele[2][10] != ele[2][22];
    ele[2][10] != ele[2][23];
    ele[2][10] != ele[2][24];
    ele[2][10] != ele[2][25];
    ele[2][10] != ele[2][26];
    ele[2][10] != ele[2][27];
    ele[2][10] != ele[2][28];
    ele[2][10] != ele[2][29];
    ele[2][10] != ele[2][30];
    ele[2][10] != ele[2][31];
    ele[2][10] != ele[2][32];
    ele[2][10] != ele[2][33];
    ele[2][10] != ele[2][34];
    ele[2][10] != ele[2][35];
    ele[2][10] != ele[20][10];
    ele[2][10] != ele[21][10];
    ele[2][10] != ele[22][10];
    ele[2][10] != ele[23][10];
    ele[2][10] != ele[24][10];
    ele[2][10] != ele[25][10];
    ele[2][10] != ele[26][10];
    ele[2][10] != ele[27][10];
    ele[2][10] != ele[28][10];
    ele[2][10] != ele[29][10];
    ele[2][10] != ele[3][10];
    ele[2][10] != ele[3][11];
    ele[2][10] != ele[3][6];
    ele[2][10] != ele[3][7];
    ele[2][10] != ele[3][8];
    ele[2][10] != ele[3][9];
    ele[2][10] != ele[30][10];
    ele[2][10] != ele[31][10];
    ele[2][10] != ele[32][10];
    ele[2][10] != ele[33][10];
    ele[2][10] != ele[34][10];
    ele[2][10] != ele[35][10];
    ele[2][10] != ele[4][10];
    ele[2][10] != ele[4][11];
    ele[2][10] != ele[4][6];
    ele[2][10] != ele[4][7];
    ele[2][10] != ele[4][8];
    ele[2][10] != ele[4][9];
    ele[2][10] != ele[5][10];
    ele[2][10] != ele[5][11];
    ele[2][10] != ele[5][6];
    ele[2][10] != ele[5][7];
    ele[2][10] != ele[5][8];
    ele[2][10] != ele[5][9];
    ele[2][10] != ele[6][10];
    ele[2][10] != ele[7][10];
    ele[2][10] != ele[8][10];
    ele[2][10] != ele[9][10];
    ele[2][11] != ele[10][11];
    ele[2][11] != ele[11][11];
    ele[2][11] != ele[12][11];
    ele[2][11] != ele[13][11];
    ele[2][11] != ele[14][11];
    ele[2][11] != ele[15][11];
    ele[2][11] != ele[16][11];
    ele[2][11] != ele[17][11];
    ele[2][11] != ele[18][11];
    ele[2][11] != ele[19][11];
    ele[2][11] != ele[2][12];
    ele[2][11] != ele[2][13];
    ele[2][11] != ele[2][14];
    ele[2][11] != ele[2][15];
    ele[2][11] != ele[2][16];
    ele[2][11] != ele[2][17];
    ele[2][11] != ele[2][18];
    ele[2][11] != ele[2][19];
    ele[2][11] != ele[2][20];
    ele[2][11] != ele[2][21];
    ele[2][11] != ele[2][22];
    ele[2][11] != ele[2][23];
    ele[2][11] != ele[2][24];
    ele[2][11] != ele[2][25];
    ele[2][11] != ele[2][26];
    ele[2][11] != ele[2][27];
    ele[2][11] != ele[2][28];
    ele[2][11] != ele[2][29];
    ele[2][11] != ele[2][30];
    ele[2][11] != ele[2][31];
    ele[2][11] != ele[2][32];
    ele[2][11] != ele[2][33];
    ele[2][11] != ele[2][34];
    ele[2][11] != ele[2][35];
    ele[2][11] != ele[20][11];
    ele[2][11] != ele[21][11];
    ele[2][11] != ele[22][11];
    ele[2][11] != ele[23][11];
    ele[2][11] != ele[24][11];
    ele[2][11] != ele[25][11];
    ele[2][11] != ele[26][11];
    ele[2][11] != ele[27][11];
    ele[2][11] != ele[28][11];
    ele[2][11] != ele[29][11];
    ele[2][11] != ele[3][10];
    ele[2][11] != ele[3][11];
    ele[2][11] != ele[3][6];
    ele[2][11] != ele[3][7];
    ele[2][11] != ele[3][8];
    ele[2][11] != ele[3][9];
    ele[2][11] != ele[30][11];
    ele[2][11] != ele[31][11];
    ele[2][11] != ele[32][11];
    ele[2][11] != ele[33][11];
    ele[2][11] != ele[34][11];
    ele[2][11] != ele[35][11];
    ele[2][11] != ele[4][10];
    ele[2][11] != ele[4][11];
    ele[2][11] != ele[4][6];
    ele[2][11] != ele[4][7];
    ele[2][11] != ele[4][8];
    ele[2][11] != ele[4][9];
    ele[2][11] != ele[5][10];
    ele[2][11] != ele[5][11];
    ele[2][11] != ele[5][6];
    ele[2][11] != ele[5][7];
    ele[2][11] != ele[5][8];
    ele[2][11] != ele[5][9];
    ele[2][11] != ele[6][11];
    ele[2][11] != ele[7][11];
    ele[2][11] != ele[8][11];
    ele[2][11] != ele[9][11];
    ele[2][12] != ele[10][12];
    ele[2][12] != ele[11][12];
    ele[2][12] != ele[12][12];
    ele[2][12] != ele[13][12];
    ele[2][12] != ele[14][12];
    ele[2][12] != ele[15][12];
    ele[2][12] != ele[16][12];
    ele[2][12] != ele[17][12];
    ele[2][12] != ele[18][12];
    ele[2][12] != ele[19][12];
    ele[2][12] != ele[2][13];
    ele[2][12] != ele[2][14];
    ele[2][12] != ele[2][15];
    ele[2][12] != ele[2][16];
    ele[2][12] != ele[2][17];
    ele[2][12] != ele[2][18];
    ele[2][12] != ele[2][19];
    ele[2][12] != ele[2][20];
    ele[2][12] != ele[2][21];
    ele[2][12] != ele[2][22];
    ele[2][12] != ele[2][23];
    ele[2][12] != ele[2][24];
    ele[2][12] != ele[2][25];
    ele[2][12] != ele[2][26];
    ele[2][12] != ele[2][27];
    ele[2][12] != ele[2][28];
    ele[2][12] != ele[2][29];
    ele[2][12] != ele[2][30];
    ele[2][12] != ele[2][31];
    ele[2][12] != ele[2][32];
    ele[2][12] != ele[2][33];
    ele[2][12] != ele[2][34];
    ele[2][12] != ele[2][35];
    ele[2][12] != ele[20][12];
    ele[2][12] != ele[21][12];
    ele[2][12] != ele[22][12];
    ele[2][12] != ele[23][12];
    ele[2][12] != ele[24][12];
    ele[2][12] != ele[25][12];
    ele[2][12] != ele[26][12];
    ele[2][12] != ele[27][12];
    ele[2][12] != ele[28][12];
    ele[2][12] != ele[29][12];
    ele[2][12] != ele[3][12];
    ele[2][12] != ele[3][13];
    ele[2][12] != ele[3][14];
    ele[2][12] != ele[3][15];
    ele[2][12] != ele[3][16];
    ele[2][12] != ele[3][17];
    ele[2][12] != ele[30][12];
    ele[2][12] != ele[31][12];
    ele[2][12] != ele[32][12];
    ele[2][12] != ele[33][12];
    ele[2][12] != ele[34][12];
    ele[2][12] != ele[35][12];
    ele[2][12] != ele[4][12];
    ele[2][12] != ele[4][13];
    ele[2][12] != ele[4][14];
    ele[2][12] != ele[4][15];
    ele[2][12] != ele[4][16];
    ele[2][12] != ele[4][17];
    ele[2][12] != ele[5][12];
    ele[2][12] != ele[5][13];
    ele[2][12] != ele[5][14];
    ele[2][12] != ele[5][15];
    ele[2][12] != ele[5][16];
    ele[2][12] != ele[5][17];
    ele[2][12] != ele[6][12];
    ele[2][12] != ele[7][12];
    ele[2][12] != ele[8][12];
    ele[2][12] != ele[9][12];
    ele[2][13] != ele[10][13];
    ele[2][13] != ele[11][13];
    ele[2][13] != ele[12][13];
    ele[2][13] != ele[13][13];
    ele[2][13] != ele[14][13];
    ele[2][13] != ele[15][13];
    ele[2][13] != ele[16][13];
    ele[2][13] != ele[17][13];
    ele[2][13] != ele[18][13];
    ele[2][13] != ele[19][13];
    ele[2][13] != ele[2][14];
    ele[2][13] != ele[2][15];
    ele[2][13] != ele[2][16];
    ele[2][13] != ele[2][17];
    ele[2][13] != ele[2][18];
    ele[2][13] != ele[2][19];
    ele[2][13] != ele[2][20];
    ele[2][13] != ele[2][21];
    ele[2][13] != ele[2][22];
    ele[2][13] != ele[2][23];
    ele[2][13] != ele[2][24];
    ele[2][13] != ele[2][25];
    ele[2][13] != ele[2][26];
    ele[2][13] != ele[2][27];
    ele[2][13] != ele[2][28];
    ele[2][13] != ele[2][29];
    ele[2][13] != ele[2][30];
    ele[2][13] != ele[2][31];
    ele[2][13] != ele[2][32];
    ele[2][13] != ele[2][33];
    ele[2][13] != ele[2][34];
    ele[2][13] != ele[2][35];
    ele[2][13] != ele[20][13];
    ele[2][13] != ele[21][13];
    ele[2][13] != ele[22][13];
    ele[2][13] != ele[23][13];
    ele[2][13] != ele[24][13];
    ele[2][13] != ele[25][13];
    ele[2][13] != ele[26][13];
    ele[2][13] != ele[27][13];
    ele[2][13] != ele[28][13];
    ele[2][13] != ele[29][13];
    ele[2][13] != ele[3][12];
    ele[2][13] != ele[3][13];
    ele[2][13] != ele[3][14];
    ele[2][13] != ele[3][15];
    ele[2][13] != ele[3][16];
    ele[2][13] != ele[3][17];
    ele[2][13] != ele[30][13];
    ele[2][13] != ele[31][13];
    ele[2][13] != ele[32][13];
    ele[2][13] != ele[33][13];
    ele[2][13] != ele[34][13];
    ele[2][13] != ele[35][13];
    ele[2][13] != ele[4][12];
    ele[2][13] != ele[4][13];
    ele[2][13] != ele[4][14];
    ele[2][13] != ele[4][15];
    ele[2][13] != ele[4][16];
    ele[2][13] != ele[4][17];
    ele[2][13] != ele[5][12];
    ele[2][13] != ele[5][13];
    ele[2][13] != ele[5][14];
    ele[2][13] != ele[5][15];
    ele[2][13] != ele[5][16];
    ele[2][13] != ele[5][17];
    ele[2][13] != ele[6][13];
    ele[2][13] != ele[7][13];
    ele[2][13] != ele[8][13];
    ele[2][13] != ele[9][13];
    ele[2][14] != ele[10][14];
    ele[2][14] != ele[11][14];
    ele[2][14] != ele[12][14];
    ele[2][14] != ele[13][14];
    ele[2][14] != ele[14][14];
    ele[2][14] != ele[15][14];
    ele[2][14] != ele[16][14];
    ele[2][14] != ele[17][14];
    ele[2][14] != ele[18][14];
    ele[2][14] != ele[19][14];
    ele[2][14] != ele[2][15];
    ele[2][14] != ele[2][16];
    ele[2][14] != ele[2][17];
    ele[2][14] != ele[2][18];
    ele[2][14] != ele[2][19];
    ele[2][14] != ele[2][20];
    ele[2][14] != ele[2][21];
    ele[2][14] != ele[2][22];
    ele[2][14] != ele[2][23];
    ele[2][14] != ele[2][24];
    ele[2][14] != ele[2][25];
    ele[2][14] != ele[2][26];
    ele[2][14] != ele[2][27];
    ele[2][14] != ele[2][28];
    ele[2][14] != ele[2][29];
    ele[2][14] != ele[2][30];
    ele[2][14] != ele[2][31];
    ele[2][14] != ele[2][32];
    ele[2][14] != ele[2][33];
    ele[2][14] != ele[2][34];
    ele[2][14] != ele[2][35];
    ele[2][14] != ele[20][14];
    ele[2][14] != ele[21][14];
    ele[2][14] != ele[22][14];
    ele[2][14] != ele[23][14];
    ele[2][14] != ele[24][14];
    ele[2][14] != ele[25][14];
    ele[2][14] != ele[26][14];
    ele[2][14] != ele[27][14];
    ele[2][14] != ele[28][14];
    ele[2][14] != ele[29][14];
    ele[2][14] != ele[3][12];
    ele[2][14] != ele[3][13];
    ele[2][14] != ele[3][14];
    ele[2][14] != ele[3][15];
    ele[2][14] != ele[3][16];
    ele[2][14] != ele[3][17];
    ele[2][14] != ele[30][14];
    ele[2][14] != ele[31][14];
    ele[2][14] != ele[32][14];
    ele[2][14] != ele[33][14];
    ele[2][14] != ele[34][14];
    ele[2][14] != ele[35][14];
    ele[2][14] != ele[4][12];
    ele[2][14] != ele[4][13];
    ele[2][14] != ele[4][14];
    ele[2][14] != ele[4][15];
    ele[2][14] != ele[4][16];
    ele[2][14] != ele[4][17];
    ele[2][14] != ele[5][12];
    ele[2][14] != ele[5][13];
    ele[2][14] != ele[5][14];
    ele[2][14] != ele[5][15];
    ele[2][14] != ele[5][16];
    ele[2][14] != ele[5][17];
    ele[2][14] != ele[6][14];
    ele[2][14] != ele[7][14];
    ele[2][14] != ele[8][14];
    ele[2][14] != ele[9][14];
    ele[2][15] != ele[10][15];
    ele[2][15] != ele[11][15];
    ele[2][15] != ele[12][15];
    ele[2][15] != ele[13][15];
    ele[2][15] != ele[14][15];
    ele[2][15] != ele[15][15];
    ele[2][15] != ele[16][15];
    ele[2][15] != ele[17][15];
    ele[2][15] != ele[18][15];
    ele[2][15] != ele[19][15];
    ele[2][15] != ele[2][16];
    ele[2][15] != ele[2][17];
    ele[2][15] != ele[2][18];
    ele[2][15] != ele[2][19];
    ele[2][15] != ele[2][20];
    ele[2][15] != ele[2][21];
    ele[2][15] != ele[2][22];
    ele[2][15] != ele[2][23];
    ele[2][15] != ele[2][24];
    ele[2][15] != ele[2][25];
    ele[2][15] != ele[2][26];
    ele[2][15] != ele[2][27];
    ele[2][15] != ele[2][28];
    ele[2][15] != ele[2][29];
    ele[2][15] != ele[2][30];
    ele[2][15] != ele[2][31];
    ele[2][15] != ele[2][32];
    ele[2][15] != ele[2][33];
    ele[2][15] != ele[2][34];
    ele[2][15] != ele[2][35];
    ele[2][15] != ele[20][15];
    ele[2][15] != ele[21][15];
    ele[2][15] != ele[22][15];
    ele[2][15] != ele[23][15];
    ele[2][15] != ele[24][15];
    ele[2][15] != ele[25][15];
    ele[2][15] != ele[26][15];
    ele[2][15] != ele[27][15];
    ele[2][15] != ele[28][15];
    ele[2][15] != ele[29][15];
    ele[2][15] != ele[3][12];
    ele[2][15] != ele[3][13];
    ele[2][15] != ele[3][14];
    ele[2][15] != ele[3][15];
    ele[2][15] != ele[3][16];
    ele[2][15] != ele[3][17];
    ele[2][15] != ele[30][15];
    ele[2][15] != ele[31][15];
    ele[2][15] != ele[32][15];
    ele[2][15] != ele[33][15];
    ele[2][15] != ele[34][15];
    ele[2][15] != ele[35][15];
    ele[2][15] != ele[4][12];
    ele[2][15] != ele[4][13];
    ele[2][15] != ele[4][14];
    ele[2][15] != ele[4][15];
    ele[2][15] != ele[4][16];
    ele[2][15] != ele[4][17];
    ele[2][15] != ele[5][12];
    ele[2][15] != ele[5][13];
    ele[2][15] != ele[5][14];
    ele[2][15] != ele[5][15];
    ele[2][15] != ele[5][16];
    ele[2][15] != ele[5][17];
    ele[2][15] != ele[6][15];
    ele[2][15] != ele[7][15];
    ele[2][15] != ele[8][15];
    ele[2][15] != ele[9][15];
    ele[2][16] != ele[10][16];
    ele[2][16] != ele[11][16];
    ele[2][16] != ele[12][16];
    ele[2][16] != ele[13][16];
    ele[2][16] != ele[14][16];
    ele[2][16] != ele[15][16];
    ele[2][16] != ele[16][16];
    ele[2][16] != ele[17][16];
    ele[2][16] != ele[18][16];
    ele[2][16] != ele[19][16];
    ele[2][16] != ele[2][17];
    ele[2][16] != ele[2][18];
    ele[2][16] != ele[2][19];
    ele[2][16] != ele[2][20];
    ele[2][16] != ele[2][21];
    ele[2][16] != ele[2][22];
    ele[2][16] != ele[2][23];
    ele[2][16] != ele[2][24];
    ele[2][16] != ele[2][25];
    ele[2][16] != ele[2][26];
    ele[2][16] != ele[2][27];
    ele[2][16] != ele[2][28];
    ele[2][16] != ele[2][29];
    ele[2][16] != ele[2][30];
    ele[2][16] != ele[2][31];
    ele[2][16] != ele[2][32];
    ele[2][16] != ele[2][33];
    ele[2][16] != ele[2][34];
    ele[2][16] != ele[2][35];
    ele[2][16] != ele[20][16];
    ele[2][16] != ele[21][16];
    ele[2][16] != ele[22][16];
    ele[2][16] != ele[23][16];
    ele[2][16] != ele[24][16];
    ele[2][16] != ele[25][16];
    ele[2][16] != ele[26][16];
    ele[2][16] != ele[27][16];
    ele[2][16] != ele[28][16];
    ele[2][16] != ele[29][16];
    ele[2][16] != ele[3][12];
    ele[2][16] != ele[3][13];
    ele[2][16] != ele[3][14];
    ele[2][16] != ele[3][15];
    ele[2][16] != ele[3][16];
    ele[2][16] != ele[3][17];
    ele[2][16] != ele[30][16];
    ele[2][16] != ele[31][16];
    ele[2][16] != ele[32][16];
    ele[2][16] != ele[33][16];
    ele[2][16] != ele[34][16];
    ele[2][16] != ele[35][16];
    ele[2][16] != ele[4][12];
    ele[2][16] != ele[4][13];
    ele[2][16] != ele[4][14];
    ele[2][16] != ele[4][15];
    ele[2][16] != ele[4][16];
    ele[2][16] != ele[4][17];
    ele[2][16] != ele[5][12];
    ele[2][16] != ele[5][13];
    ele[2][16] != ele[5][14];
    ele[2][16] != ele[5][15];
    ele[2][16] != ele[5][16];
    ele[2][16] != ele[5][17];
    ele[2][16] != ele[6][16];
    ele[2][16] != ele[7][16];
    ele[2][16] != ele[8][16];
    ele[2][16] != ele[9][16];
    ele[2][17] != ele[10][17];
    ele[2][17] != ele[11][17];
    ele[2][17] != ele[12][17];
    ele[2][17] != ele[13][17];
    ele[2][17] != ele[14][17];
    ele[2][17] != ele[15][17];
    ele[2][17] != ele[16][17];
    ele[2][17] != ele[17][17];
    ele[2][17] != ele[18][17];
    ele[2][17] != ele[19][17];
    ele[2][17] != ele[2][18];
    ele[2][17] != ele[2][19];
    ele[2][17] != ele[2][20];
    ele[2][17] != ele[2][21];
    ele[2][17] != ele[2][22];
    ele[2][17] != ele[2][23];
    ele[2][17] != ele[2][24];
    ele[2][17] != ele[2][25];
    ele[2][17] != ele[2][26];
    ele[2][17] != ele[2][27];
    ele[2][17] != ele[2][28];
    ele[2][17] != ele[2][29];
    ele[2][17] != ele[2][30];
    ele[2][17] != ele[2][31];
    ele[2][17] != ele[2][32];
    ele[2][17] != ele[2][33];
    ele[2][17] != ele[2][34];
    ele[2][17] != ele[2][35];
    ele[2][17] != ele[20][17];
    ele[2][17] != ele[21][17];
    ele[2][17] != ele[22][17];
    ele[2][17] != ele[23][17];
    ele[2][17] != ele[24][17];
    ele[2][17] != ele[25][17];
    ele[2][17] != ele[26][17];
    ele[2][17] != ele[27][17];
    ele[2][17] != ele[28][17];
    ele[2][17] != ele[29][17];
    ele[2][17] != ele[3][12];
    ele[2][17] != ele[3][13];
    ele[2][17] != ele[3][14];
    ele[2][17] != ele[3][15];
    ele[2][17] != ele[3][16];
    ele[2][17] != ele[3][17];
    ele[2][17] != ele[30][17];
    ele[2][17] != ele[31][17];
    ele[2][17] != ele[32][17];
    ele[2][17] != ele[33][17];
    ele[2][17] != ele[34][17];
    ele[2][17] != ele[35][17];
    ele[2][17] != ele[4][12];
    ele[2][17] != ele[4][13];
    ele[2][17] != ele[4][14];
    ele[2][17] != ele[4][15];
    ele[2][17] != ele[4][16];
    ele[2][17] != ele[4][17];
    ele[2][17] != ele[5][12];
    ele[2][17] != ele[5][13];
    ele[2][17] != ele[5][14];
    ele[2][17] != ele[5][15];
    ele[2][17] != ele[5][16];
    ele[2][17] != ele[5][17];
    ele[2][17] != ele[6][17];
    ele[2][17] != ele[7][17];
    ele[2][17] != ele[8][17];
    ele[2][17] != ele[9][17];
    ele[2][18] != ele[10][18];
    ele[2][18] != ele[11][18];
    ele[2][18] != ele[12][18];
    ele[2][18] != ele[13][18];
    ele[2][18] != ele[14][18];
    ele[2][18] != ele[15][18];
    ele[2][18] != ele[16][18];
    ele[2][18] != ele[17][18];
    ele[2][18] != ele[18][18];
    ele[2][18] != ele[19][18];
    ele[2][18] != ele[2][19];
    ele[2][18] != ele[2][20];
    ele[2][18] != ele[2][21];
    ele[2][18] != ele[2][22];
    ele[2][18] != ele[2][23];
    ele[2][18] != ele[2][24];
    ele[2][18] != ele[2][25];
    ele[2][18] != ele[2][26];
    ele[2][18] != ele[2][27];
    ele[2][18] != ele[2][28];
    ele[2][18] != ele[2][29];
    ele[2][18] != ele[2][30];
    ele[2][18] != ele[2][31];
    ele[2][18] != ele[2][32];
    ele[2][18] != ele[2][33];
    ele[2][18] != ele[2][34];
    ele[2][18] != ele[2][35];
    ele[2][18] != ele[20][18];
    ele[2][18] != ele[21][18];
    ele[2][18] != ele[22][18];
    ele[2][18] != ele[23][18];
    ele[2][18] != ele[24][18];
    ele[2][18] != ele[25][18];
    ele[2][18] != ele[26][18];
    ele[2][18] != ele[27][18];
    ele[2][18] != ele[28][18];
    ele[2][18] != ele[29][18];
    ele[2][18] != ele[3][18];
    ele[2][18] != ele[3][19];
    ele[2][18] != ele[3][20];
    ele[2][18] != ele[3][21];
    ele[2][18] != ele[3][22];
    ele[2][18] != ele[3][23];
    ele[2][18] != ele[30][18];
    ele[2][18] != ele[31][18];
    ele[2][18] != ele[32][18];
    ele[2][18] != ele[33][18];
    ele[2][18] != ele[34][18];
    ele[2][18] != ele[35][18];
    ele[2][18] != ele[4][18];
    ele[2][18] != ele[4][19];
    ele[2][18] != ele[4][20];
    ele[2][18] != ele[4][21];
    ele[2][18] != ele[4][22];
    ele[2][18] != ele[4][23];
    ele[2][18] != ele[5][18];
    ele[2][18] != ele[5][19];
    ele[2][18] != ele[5][20];
    ele[2][18] != ele[5][21];
    ele[2][18] != ele[5][22];
    ele[2][18] != ele[5][23];
    ele[2][18] != ele[6][18];
    ele[2][18] != ele[7][18];
    ele[2][18] != ele[8][18];
    ele[2][18] != ele[9][18];
    ele[2][19] != ele[10][19];
    ele[2][19] != ele[11][19];
    ele[2][19] != ele[12][19];
    ele[2][19] != ele[13][19];
    ele[2][19] != ele[14][19];
    ele[2][19] != ele[15][19];
    ele[2][19] != ele[16][19];
    ele[2][19] != ele[17][19];
    ele[2][19] != ele[18][19];
    ele[2][19] != ele[19][19];
    ele[2][19] != ele[2][20];
    ele[2][19] != ele[2][21];
    ele[2][19] != ele[2][22];
    ele[2][19] != ele[2][23];
    ele[2][19] != ele[2][24];
    ele[2][19] != ele[2][25];
    ele[2][19] != ele[2][26];
    ele[2][19] != ele[2][27];
    ele[2][19] != ele[2][28];
    ele[2][19] != ele[2][29];
    ele[2][19] != ele[2][30];
    ele[2][19] != ele[2][31];
    ele[2][19] != ele[2][32];
    ele[2][19] != ele[2][33];
    ele[2][19] != ele[2][34];
    ele[2][19] != ele[2][35];
    ele[2][19] != ele[20][19];
    ele[2][19] != ele[21][19];
    ele[2][19] != ele[22][19];
    ele[2][19] != ele[23][19];
    ele[2][19] != ele[24][19];
    ele[2][19] != ele[25][19];
    ele[2][19] != ele[26][19];
    ele[2][19] != ele[27][19];
    ele[2][19] != ele[28][19];
    ele[2][19] != ele[29][19];
    ele[2][19] != ele[3][18];
    ele[2][19] != ele[3][19];
    ele[2][19] != ele[3][20];
    ele[2][19] != ele[3][21];
    ele[2][19] != ele[3][22];
    ele[2][19] != ele[3][23];
    ele[2][19] != ele[30][19];
    ele[2][19] != ele[31][19];
    ele[2][19] != ele[32][19];
    ele[2][19] != ele[33][19];
    ele[2][19] != ele[34][19];
    ele[2][19] != ele[35][19];
    ele[2][19] != ele[4][18];
    ele[2][19] != ele[4][19];
    ele[2][19] != ele[4][20];
    ele[2][19] != ele[4][21];
    ele[2][19] != ele[4][22];
    ele[2][19] != ele[4][23];
    ele[2][19] != ele[5][18];
    ele[2][19] != ele[5][19];
    ele[2][19] != ele[5][20];
    ele[2][19] != ele[5][21];
    ele[2][19] != ele[5][22];
    ele[2][19] != ele[5][23];
    ele[2][19] != ele[6][19];
    ele[2][19] != ele[7][19];
    ele[2][19] != ele[8][19];
    ele[2][19] != ele[9][19];
    ele[2][2] != ele[10][2];
    ele[2][2] != ele[11][2];
    ele[2][2] != ele[12][2];
    ele[2][2] != ele[13][2];
    ele[2][2] != ele[14][2];
    ele[2][2] != ele[15][2];
    ele[2][2] != ele[16][2];
    ele[2][2] != ele[17][2];
    ele[2][2] != ele[18][2];
    ele[2][2] != ele[19][2];
    ele[2][2] != ele[2][10];
    ele[2][2] != ele[2][11];
    ele[2][2] != ele[2][12];
    ele[2][2] != ele[2][13];
    ele[2][2] != ele[2][14];
    ele[2][2] != ele[2][15];
    ele[2][2] != ele[2][16];
    ele[2][2] != ele[2][17];
    ele[2][2] != ele[2][18];
    ele[2][2] != ele[2][19];
    ele[2][2] != ele[2][20];
    ele[2][2] != ele[2][21];
    ele[2][2] != ele[2][22];
    ele[2][2] != ele[2][23];
    ele[2][2] != ele[2][24];
    ele[2][2] != ele[2][25];
    ele[2][2] != ele[2][26];
    ele[2][2] != ele[2][27];
    ele[2][2] != ele[2][28];
    ele[2][2] != ele[2][29];
    ele[2][2] != ele[2][3];
    ele[2][2] != ele[2][30];
    ele[2][2] != ele[2][31];
    ele[2][2] != ele[2][32];
    ele[2][2] != ele[2][33];
    ele[2][2] != ele[2][34];
    ele[2][2] != ele[2][35];
    ele[2][2] != ele[2][4];
    ele[2][2] != ele[2][5];
    ele[2][2] != ele[2][6];
    ele[2][2] != ele[2][7];
    ele[2][2] != ele[2][8];
    ele[2][2] != ele[2][9];
    ele[2][2] != ele[20][2];
    ele[2][2] != ele[21][2];
    ele[2][2] != ele[22][2];
    ele[2][2] != ele[23][2];
    ele[2][2] != ele[24][2];
    ele[2][2] != ele[25][2];
    ele[2][2] != ele[26][2];
    ele[2][2] != ele[27][2];
    ele[2][2] != ele[28][2];
    ele[2][2] != ele[29][2];
    ele[2][2] != ele[3][0];
    ele[2][2] != ele[3][1];
    ele[2][2] != ele[3][2];
    ele[2][2] != ele[3][3];
    ele[2][2] != ele[3][4];
    ele[2][2] != ele[3][5];
    ele[2][2] != ele[30][2];
    ele[2][2] != ele[31][2];
    ele[2][2] != ele[32][2];
    ele[2][2] != ele[33][2];
    ele[2][2] != ele[34][2];
    ele[2][2] != ele[35][2];
    ele[2][2] != ele[4][0];
    ele[2][2] != ele[4][1];
    ele[2][2] != ele[4][2];
    ele[2][2] != ele[4][3];
    ele[2][2] != ele[4][4];
    ele[2][2] != ele[4][5];
    ele[2][2] != ele[5][0];
    ele[2][2] != ele[5][1];
    ele[2][2] != ele[5][2];
    ele[2][2] != ele[5][3];
    ele[2][2] != ele[5][4];
    ele[2][2] != ele[5][5];
    ele[2][2] != ele[6][2];
    ele[2][2] != ele[7][2];
    ele[2][2] != ele[8][2];
    ele[2][2] != ele[9][2];
    ele[2][20] != ele[10][20];
    ele[2][20] != ele[11][20];
    ele[2][20] != ele[12][20];
    ele[2][20] != ele[13][20];
    ele[2][20] != ele[14][20];
    ele[2][20] != ele[15][20];
    ele[2][20] != ele[16][20];
    ele[2][20] != ele[17][20];
    ele[2][20] != ele[18][20];
    ele[2][20] != ele[19][20];
    ele[2][20] != ele[2][21];
    ele[2][20] != ele[2][22];
    ele[2][20] != ele[2][23];
    ele[2][20] != ele[2][24];
    ele[2][20] != ele[2][25];
    ele[2][20] != ele[2][26];
    ele[2][20] != ele[2][27];
    ele[2][20] != ele[2][28];
    ele[2][20] != ele[2][29];
    ele[2][20] != ele[2][30];
    ele[2][20] != ele[2][31];
    ele[2][20] != ele[2][32];
    ele[2][20] != ele[2][33];
    ele[2][20] != ele[2][34];
    ele[2][20] != ele[2][35];
    ele[2][20] != ele[20][20];
    ele[2][20] != ele[21][20];
    ele[2][20] != ele[22][20];
    ele[2][20] != ele[23][20];
    ele[2][20] != ele[24][20];
    ele[2][20] != ele[25][20];
    ele[2][20] != ele[26][20];
    ele[2][20] != ele[27][20];
    ele[2][20] != ele[28][20];
    ele[2][20] != ele[29][20];
    ele[2][20] != ele[3][18];
    ele[2][20] != ele[3][19];
    ele[2][20] != ele[3][20];
    ele[2][20] != ele[3][21];
    ele[2][20] != ele[3][22];
    ele[2][20] != ele[3][23];
    ele[2][20] != ele[30][20];
    ele[2][20] != ele[31][20];
    ele[2][20] != ele[32][20];
    ele[2][20] != ele[33][20];
    ele[2][20] != ele[34][20];
    ele[2][20] != ele[35][20];
    ele[2][20] != ele[4][18];
    ele[2][20] != ele[4][19];
    ele[2][20] != ele[4][20];
    ele[2][20] != ele[4][21];
    ele[2][20] != ele[4][22];
    ele[2][20] != ele[4][23];
    ele[2][20] != ele[5][18];
    ele[2][20] != ele[5][19];
    ele[2][20] != ele[5][20];
    ele[2][20] != ele[5][21];
    ele[2][20] != ele[5][22];
    ele[2][20] != ele[5][23];
    ele[2][20] != ele[6][20];
    ele[2][20] != ele[7][20];
    ele[2][20] != ele[8][20];
    ele[2][20] != ele[9][20];
    ele[2][21] != ele[10][21];
    ele[2][21] != ele[11][21];
    ele[2][21] != ele[12][21];
    ele[2][21] != ele[13][21];
    ele[2][21] != ele[14][21];
    ele[2][21] != ele[15][21];
    ele[2][21] != ele[16][21];
    ele[2][21] != ele[17][21];
    ele[2][21] != ele[18][21];
    ele[2][21] != ele[19][21];
    ele[2][21] != ele[2][22];
    ele[2][21] != ele[2][23];
    ele[2][21] != ele[2][24];
    ele[2][21] != ele[2][25];
    ele[2][21] != ele[2][26];
    ele[2][21] != ele[2][27];
    ele[2][21] != ele[2][28];
    ele[2][21] != ele[2][29];
    ele[2][21] != ele[2][30];
    ele[2][21] != ele[2][31];
    ele[2][21] != ele[2][32];
    ele[2][21] != ele[2][33];
    ele[2][21] != ele[2][34];
    ele[2][21] != ele[2][35];
    ele[2][21] != ele[20][21];
    ele[2][21] != ele[21][21];
    ele[2][21] != ele[22][21];
    ele[2][21] != ele[23][21];
    ele[2][21] != ele[24][21];
    ele[2][21] != ele[25][21];
    ele[2][21] != ele[26][21];
    ele[2][21] != ele[27][21];
    ele[2][21] != ele[28][21];
    ele[2][21] != ele[29][21];
    ele[2][21] != ele[3][18];
    ele[2][21] != ele[3][19];
    ele[2][21] != ele[3][20];
    ele[2][21] != ele[3][21];
    ele[2][21] != ele[3][22];
    ele[2][21] != ele[3][23];
    ele[2][21] != ele[30][21];
    ele[2][21] != ele[31][21];
    ele[2][21] != ele[32][21];
    ele[2][21] != ele[33][21];
    ele[2][21] != ele[34][21];
    ele[2][21] != ele[35][21];
    ele[2][21] != ele[4][18];
    ele[2][21] != ele[4][19];
    ele[2][21] != ele[4][20];
    ele[2][21] != ele[4][21];
    ele[2][21] != ele[4][22];
    ele[2][21] != ele[4][23];
    ele[2][21] != ele[5][18];
    ele[2][21] != ele[5][19];
    ele[2][21] != ele[5][20];
    ele[2][21] != ele[5][21];
    ele[2][21] != ele[5][22];
    ele[2][21] != ele[5][23];
    ele[2][21] != ele[6][21];
    ele[2][21] != ele[7][21];
    ele[2][21] != ele[8][21];
    ele[2][21] != ele[9][21];
    ele[2][22] != ele[10][22];
    ele[2][22] != ele[11][22];
    ele[2][22] != ele[12][22];
    ele[2][22] != ele[13][22];
    ele[2][22] != ele[14][22];
    ele[2][22] != ele[15][22];
    ele[2][22] != ele[16][22];
    ele[2][22] != ele[17][22];
    ele[2][22] != ele[18][22];
    ele[2][22] != ele[19][22];
    ele[2][22] != ele[2][23];
    ele[2][22] != ele[2][24];
    ele[2][22] != ele[2][25];
    ele[2][22] != ele[2][26];
    ele[2][22] != ele[2][27];
    ele[2][22] != ele[2][28];
    ele[2][22] != ele[2][29];
    ele[2][22] != ele[2][30];
    ele[2][22] != ele[2][31];
    ele[2][22] != ele[2][32];
    ele[2][22] != ele[2][33];
    ele[2][22] != ele[2][34];
    ele[2][22] != ele[2][35];
    ele[2][22] != ele[20][22];
    ele[2][22] != ele[21][22];
    ele[2][22] != ele[22][22];
    ele[2][22] != ele[23][22];
    ele[2][22] != ele[24][22];
    ele[2][22] != ele[25][22];
    ele[2][22] != ele[26][22];
    ele[2][22] != ele[27][22];
    ele[2][22] != ele[28][22];
    ele[2][22] != ele[29][22];
    ele[2][22] != ele[3][18];
    ele[2][22] != ele[3][19];
    ele[2][22] != ele[3][20];
    ele[2][22] != ele[3][21];
    ele[2][22] != ele[3][22];
    ele[2][22] != ele[3][23];
    ele[2][22] != ele[30][22];
    ele[2][22] != ele[31][22];
    ele[2][22] != ele[32][22];
    ele[2][22] != ele[33][22];
    ele[2][22] != ele[34][22];
    ele[2][22] != ele[35][22];
    ele[2][22] != ele[4][18];
    ele[2][22] != ele[4][19];
    ele[2][22] != ele[4][20];
    ele[2][22] != ele[4][21];
    ele[2][22] != ele[4][22];
    ele[2][22] != ele[4][23];
    ele[2][22] != ele[5][18];
    ele[2][22] != ele[5][19];
    ele[2][22] != ele[5][20];
    ele[2][22] != ele[5][21];
    ele[2][22] != ele[5][22];
    ele[2][22] != ele[5][23];
    ele[2][22] != ele[6][22];
    ele[2][22] != ele[7][22];
    ele[2][22] != ele[8][22];
    ele[2][22] != ele[9][22];
    ele[2][23] != ele[10][23];
    ele[2][23] != ele[11][23];
    ele[2][23] != ele[12][23];
    ele[2][23] != ele[13][23];
    ele[2][23] != ele[14][23];
    ele[2][23] != ele[15][23];
    ele[2][23] != ele[16][23];
    ele[2][23] != ele[17][23];
    ele[2][23] != ele[18][23];
    ele[2][23] != ele[19][23];
    ele[2][23] != ele[2][24];
    ele[2][23] != ele[2][25];
    ele[2][23] != ele[2][26];
    ele[2][23] != ele[2][27];
    ele[2][23] != ele[2][28];
    ele[2][23] != ele[2][29];
    ele[2][23] != ele[2][30];
    ele[2][23] != ele[2][31];
    ele[2][23] != ele[2][32];
    ele[2][23] != ele[2][33];
    ele[2][23] != ele[2][34];
    ele[2][23] != ele[2][35];
    ele[2][23] != ele[20][23];
    ele[2][23] != ele[21][23];
    ele[2][23] != ele[22][23];
    ele[2][23] != ele[23][23];
    ele[2][23] != ele[24][23];
    ele[2][23] != ele[25][23];
    ele[2][23] != ele[26][23];
    ele[2][23] != ele[27][23];
    ele[2][23] != ele[28][23];
    ele[2][23] != ele[29][23];
    ele[2][23] != ele[3][18];
    ele[2][23] != ele[3][19];
    ele[2][23] != ele[3][20];
    ele[2][23] != ele[3][21];
    ele[2][23] != ele[3][22];
    ele[2][23] != ele[3][23];
    ele[2][23] != ele[30][23];
    ele[2][23] != ele[31][23];
    ele[2][23] != ele[32][23];
    ele[2][23] != ele[33][23];
    ele[2][23] != ele[34][23];
    ele[2][23] != ele[35][23];
    ele[2][23] != ele[4][18];
    ele[2][23] != ele[4][19];
    ele[2][23] != ele[4][20];
    ele[2][23] != ele[4][21];
    ele[2][23] != ele[4][22];
    ele[2][23] != ele[4][23];
    ele[2][23] != ele[5][18];
    ele[2][23] != ele[5][19];
    ele[2][23] != ele[5][20];
    ele[2][23] != ele[5][21];
    ele[2][23] != ele[5][22];
    ele[2][23] != ele[5][23];
    ele[2][23] != ele[6][23];
    ele[2][23] != ele[7][23];
    ele[2][23] != ele[8][23];
    ele[2][23] != ele[9][23];
    ele[2][24] != ele[10][24];
    ele[2][24] != ele[11][24];
    ele[2][24] != ele[12][24];
    ele[2][24] != ele[13][24];
    ele[2][24] != ele[14][24];
    ele[2][24] != ele[15][24];
    ele[2][24] != ele[16][24];
    ele[2][24] != ele[17][24];
    ele[2][24] != ele[18][24];
    ele[2][24] != ele[19][24];
    ele[2][24] != ele[2][25];
    ele[2][24] != ele[2][26];
    ele[2][24] != ele[2][27];
    ele[2][24] != ele[2][28];
    ele[2][24] != ele[2][29];
    ele[2][24] != ele[2][30];
    ele[2][24] != ele[2][31];
    ele[2][24] != ele[2][32];
    ele[2][24] != ele[2][33];
    ele[2][24] != ele[2][34];
    ele[2][24] != ele[2][35];
    ele[2][24] != ele[20][24];
    ele[2][24] != ele[21][24];
    ele[2][24] != ele[22][24];
    ele[2][24] != ele[23][24];
    ele[2][24] != ele[24][24];
    ele[2][24] != ele[25][24];
    ele[2][24] != ele[26][24];
    ele[2][24] != ele[27][24];
    ele[2][24] != ele[28][24];
    ele[2][24] != ele[29][24];
    ele[2][24] != ele[3][24];
    ele[2][24] != ele[3][25];
    ele[2][24] != ele[3][26];
    ele[2][24] != ele[3][27];
    ele[2][24] != ele[3][28];
    ele[2][24] != ele[3][29];
    ele[2][24] != ele[30][24];
    ele[2][24] != ele[31][24];
    ele[2][24] != ele[32][24];
    ele[2][24] != ele[33][24];
    ele[2][24] != ele[34][24];
    ele[2][24] != ele[35][24];
    ele[2][24] != ele[4][24];
    ele[2][24] != ele[4][25];
    ele[2][24] != ele[4][26];
    ele[2][24] != ele[4][27];
    ele[2][24] != ele[4][28];
    ele[2][24] != ele[4][29];
    ele[2][24] != ele[5][24];
    ele[2][24] != ele[5][25];
    ele[2][24] != ele[5][26];
    ele[2][24] != ele[5][27];
    ele[2][24] != ele[5][28];
    ele[2][24] != ele[5][29];
    ele[2][24] != ele[6][24];
    ele[2][24] != ele[7][24];
    ele[2][24] != ele[8][24];
    ele[2][24] != ele[9][24];
    ele[2][25] != ele[10][25];
    ele[2][25] != ele[11][25];
    ele[2][25] != ele[12][25];
    ele[2][25] != ele[13][25];
    ele[2][25] != ele[14][25];
    ele[2][25] != ele[15][25];
    ele[2][25] != ele[16][25];
    ele[2][25] != ele[17][25];
    ele[2][25] != ele[18][25];
    ele[2][25] != ele[19][25];
    ele[2][25] != ele[2][26];
    ele[2][25] != ele[2][27];
    ele[2][25] != ele[2][28];
    ele[2][25] != ele[2][29];
    ele[2][25] != ele[2][30];
    ele[2][25] != ele[2][31];
    ele[2][25] != ele[2][32];
    ele[2][25] != ele[2][33];
    ele[2][25] != ele[2][34];
    ele[2][25] != ele[2][35];
    ele[2][25] != ele[20][25];
    ele[2][25] != ele[21][25];
    ele[2][25] != ele[22][25];
    ele[2][25] != ele[23][25];
    ele[2][25] != ele[24][25];
    ele[2][25] != ele[25][25];
    ele[2][25] != ele[26][25];
    ele[2][25] != ele[27][25];
    ele[2][25] != ele[28][25];
    ele[2][25] != ele[29][25];
    ele[2][25] != ele[3][24];
    ele[2][25] != ele[3][25];
    ele[2][25] != ele[3][26];
    ele[2][25] != ele[3][27];
    ele[2][25] != ele[3][28];
    ele[2][25] != ele[3][29];
    ele[2][25] != ele[30][25];
    ele[2][25] != ele[31][25];
    ele[2][25] != ele[32][25];
    ele[2][25] != ele[33][25];
    ele[2][25] != ele[34][25];
    ele[2][25] != ele[35][25];
    ele[2][25] != ele[4][24];
    ele[2][25] != ele[4][25];
    ele[2][25] != ele[4][26];
    ele[2][25] != ele[4][27];
    ele[2][25] != ele[4][28];
    ele[2][25] != ele[4][29];
    ele[2][25] != ele[5][24];
    ele[2][25] != ele[5][25];
    ele[2][25] != ele[5][26];
    ele[2][25] != ele[5][27];
    ele[2][25] != ele[5][28];
    ele[2][25] != ele[5][29];
    ele[2][25] != ele[6][25];
    ele[2][25] != ele[7][25];
    ele[2][25] != ele[8][25];
    ele[2][25] != ele[9][25];
    ele[2][26] != ele[10][26];
    ele[2][26] != ele[11][26];
    ele[2][26] != ele[12][26];
    ele[2][26] != ele[13][26];
    ele[2][26] != ele[14][26];
    ele[2][26] != ele[15][26];
    ele[2][26] != ele[16][26];
    ele[2][26] != ele[17][26];
    ele[2][26] != ele[18][26];
    ele[2][26] != ele[19][26];
    ele[2][26] != ele[2][27];
    ele[2][26] != ele[2][28];
    ele[2][26] != ele[2][29];
    ele[2][26] != ele[2][30];
    ele[2][26] != ele[2][31];
    ele[2][26] != ele[2][32];
    ele[2][26] != ele[2][33];
    ele[2][26] != ele[2][34];
    ele[2][26] != ele[2][35];
    ele[2][26] != ele[20][26];
    ele[2][26] != ele[21][26];
    ele[2][26] != ele[22][26];
    ele[2][26] != ele[23][26];
    ele[2][26] != ele[24][26];
    ele[2][26] != ele[25][26];
    ele[2][26] != ele[26][26];
    ele[2][26] != ele[27][26];
    ele[2][26] != ele[28][26];
    ele[2][26] != ele[29][26];
    ele[2][26] != ele[3][24];
    ele[2][26] != ele[3][25];
    ele[2][26] != ele[3][26];
    ele[2][26] != ele[3][27];
    ele[2][26] != ele[3][28];
    ele[2][26] != ele[3][29];
    ele[2][26] != ele[30][26];
    ele[2][26] != ele[31][26];
    ele[2][26] != ele[32][26];
    ele[2][26] != ele[33][26];
    ele[2][26] != ele[34][26];
    ele[2][26] != ele[35][26];
    ele[2][26] != ele[4][24];
    ele[2][26] != ele[4][25];
    ele[2][26] != ele[4][26];
    ele[2][26] != ele[4][27];
    ele[2][26] != ele[4][28];
    ele[2][26] != ele[4][29];
    ele[2][26] != ele[5][24];
    ele[2][26] != ele[5][25];
    ele[2][26] != ele[5][26];
    ele[2][26] != ele[5][27];
    ele[2][26] != ele[5][28];
    ele[2][26] != ele[5][29];
    ele[2][26] != ele[6][26];
    ele[2][26] != ele[7][26];
    ele[2][26] != ele[8][26];
    ele[2][26] != ele[9][26];
    ele[2][27] != ele[10][27];
    ele[2][27] != ele[11][27];
    ele[2][27] != ele[12][27];
    ele[2][27] != ele[13][27];
    ele[2][27] != ele[14][27];
    ele[2][27] != ele[15][27];
    ele[2][27] != ele[16][27];
    ele[2][27] != ele[17][27];
    ele[2][27] != ele[18][27];
    ele[2][27] != ele[19][27];
    ele[2][27] != ele[2][28];
    ele[2][27] != ele[2][29];
    ele[2][27] != ele[2][30];
    ele[2][27] != ele[2][31];
    ele[2][27] != ele[2][32];
    ele[2][27] != ele[2][33];
    ele[2][27] != ele[2][34];
    ele[2][27] != ele[2][35];
    ele[2][27] != ele[20][27];
    ele[2][27] != ele[21][27];
    ele[2][27] != ele[22][27];
    ele[2][27] != ele[23][27];
    ele[2][27] != ele[24][27];
    ele[2][27] != ele[25][27];
    ele[2][27] != ele[26][27];
    ele[2][27] != ele[27][27];
    ele[2][27] != ele[28][27];
    ele[2][27] != ele[29][27];
    ele[2][27] != ele[3][24];
    ele[2][27] != ele[3][25];
    ele[2][27] != ele[3][26];
    ele[2][27] != ele[3][27];
    ele[2][27] != ele[3][28];
    ele[2][27] != ele[3][29];
    ele[2][27] != ele[30][27];
    ele[2][27] != ele[31][27];
    ele[2][27] != ele[32][27];
    ele[2][27] != ele[33][27];
    ele[2][27] != ele[34][27];
    ele[2][27] != ele[35][27];
    ele[2][27] != ele[4][24];
    ele[2][27] != ele[4][25];
    ele[2][27] != ele[4][26];
    ele[2][27] != ele[4][27];
    ele[2][27] != ele[4][28];
    ele[2][27] != ele[4][29];
    ele[2][27] != ele[5][24];
    ele[2][27] != ele[5][25];
    ele[2][27] != ele[5][26];
    ele[2][27] != ele[5][27];
    ele[2][27] != ele[5][28];
    ele[2][27] != ele[5][29];
    ele[2][27] != ele[6][27];
    ele[2][27] != ele[7][27];
    ele[2][27] != ele[8][27];
    ele[2][27] != ele[9][27];
    ele[2][28] != ele[10][28];
    ele[2][28] != ele[11][28];
    ele[2][28] != ele[12][28];
    ele[2][28] != ele[13][28];
    ele[2][28] != ele[14][28];
    ele[2][28] != ele[15][28];
    ele[2][28] != ele[16][28];
    ele[2][28] != ele[17][28];
    ele[2][28] != ele[18][28];
    ele[2][28] != ele[19][28];
    ele[2][28] != ele[2][29];
    ele[2][28] != ele[2][30];
    ele[2][28] != ele[2][31];
    ele[2][28] != ele[2][32];
    ele[2][28] != ele[2][33];
    ele[2][28] != ele[2][34];
    ele[2][28] != ele[2][35];
    ele[2][28] != ele[20][28];
    ele[2][28] != ele[21][28];
    ele[2][28] != ele[22][28];
    ele[2][28] != ele[23][28];
    ele[2][28] != ele[24][28];
    ele[2][28] != ele[25][28];
    ele[2][28] != ele[26][28];
    ele[2][28] != ele[27][28];
    ele[2][28] != ele[28][28];
    ele[2][28] != ele[29][28];
    ele[2][28] != ele[3][24];
    ele[2][28] != ele[3][25];
    ele[2][28] != ele[3][26];
    ele[2][28] != ele[3][27];
    ele[2][28] != ele[3][28];
    ele[2][28] != ele[3][29];
    ele[2][28] != ele[30][28];
    ele[2][28] != ele[31][28];
    ele[2][28] != ele[32][28];
    ele[2][28] != ele[33][28];
    ele[2][28] != ele[34][28];
    ele[2][28] != ele[35][28];
    ele[2][28] != ele[4][24];
    ele[2][28] != ele[4][25];
    ele[2][28] != ele[4][26];
    ele[2][28] != ele[4][27];
    ele[2][28] != ele[4][28];
    ele[2][28] != ele[4][29];
    ele[2][28] != ele[5][24];
    ele[2][28] != ele[5][25];
    ele[2][28] != ele[5][26];
    ele[2][28] != ele[5][27];
    ele[2][28] != ele[5][28];
    ele[2][28] != ele[5][29];
    ele[2][28] != ele[6][28];
    ele[2][28] != ele[7][28];
    ele[2][28] != ele[8][28];
    ele[2][28] != ele[9][28];
    ele[2][29] != ele[10][29];
    ele[2][29] != ele[11][29];
    ele[2][29] != ele[12][29];
    ele[2][29] != ele[13][29];
    ele[2][29] != ele[14][29];
    ele[2][29] != ele[15][29];
    ele[2][29] != ele[16][29];
    ele[2][29] != ele[17][29];
    ele[2][29] != ele[18][29];
    ele[2][29] != ele[19][29];
    ele[2][29] != ele[2][30];
    ele[2][29] != ele[2][31];
    ele[2][29] != ele[2][32];
    ele[2][29] != ele[2][33];
    ele[2][29] != ele[2][34];
    ele[2][29] != ele[2][35];
    ele[2][29] != ele[20][29];
    ele[2][29] != ele[21][29];
    ele[2][29] != ele[22][29];
    ele[2][29] != ele[23][29];
    ele[2][29] != ele[24][29];
    ele[2][29] != ele[25][29];
    ele[2][29] != ele[26][29];
    ele[2][29] != ele[27][29];
    ele[2][29] != ele[28][29];
    ele[2][29] != ele[29][29];
    ele[2][29] != ele[3][24];
    ele[2][29] != ele[3][25];
    ele[2][29] != ele[3][26];
    ele[2][29] != ele[3][27];
    ele[2][29] != ele[3][28];
    ele[2][29] != ele[3][29];
    ele[2][29] != ele[30][29];
    ele[2][29] != ele[31][29];
    ele[2][29] != ele[32][29];
    ele[2][29] != ele[33][29];
    ele[2][29] != ele[34][29];
    ele[2][29] != ele[35][29];
    ele[2][29] != ele[4][24];
    ele[2][29] != ele[4][25];
    ele[2][29] != ele[4][26];
    ele[2][29] != ele[4][27];
    ele[2][29] != ele[4][28];
    ele[2][29] != ele[4][29];
    ele[2][29] != ele[5][24];
    ele[2][29] != ele[5][25];
    ele[2][29] != ele[5][26];
    ele[2][29] != ele[5][27];
    ele[2][29] != ele[5][28];
    ele[2][29] != ele[5][29];
    ele[2][29] != ele[6][29];
    ele[2][29] != ele[7][29];
    ele[2][29] != ele[8][29];
    ele[2][29] != ele[9][29];
    ele[2][3] != ele[10][3];
    ele[2][3] != ele[11][3];
    ele[2][3] != ele[12][3];
    ele[2][3] != ele[13][3];
    ele[2][3] != ele[14][3];
    ele[2][3] != ele[15][3];
    ele[2][3] != ele[16][3];
    ele[2][3] != ele[17][3];
    ele[2][3] != ele[18][3];
    ele[2][3] != ele[19][3];
    ele[2][3] != ele[2][10];
    ele[2][3] != ele[2][11];
    ele[2][3] != ele[2][12];
    ele[2][3] != ele[2][13];
    ele[2][3] != ele[2][14];
    ele[2][3] != ele[2][15];
    ele[2][3] != ele[2][16];
    ele[2][3] != ele[2][17];
    ele[2][3] != ele[2][18];
    ele[2][3] != ele[2][19];
    ele[2][3] != ele[2][20];
    ele[2][3] != ele[2][21];
    ele[2][3] != ele[2][22];
    ele[2][3] != ele[2][23];
    ele[2][3] != ele[2][24];
    ele[2][3] != ele[2][25];
    ele[2][3] != ele[2][26];
    ele[2][3] != ele[2][27];
    ele[2][3] != ele[2][28];
    ele[2][3] != ele[2][29];
    ele[2][3] != ele[2][30];
    ele[2][3] != ele[2][31];
    ele[2][3] != ele[2][32];
    ele[2][3] != ele[2][33];
    ele[2][3] != ele[2][34];
    ele[2][3] != ele[2][35];
    ele[2][3] != ele[2][4];
    ele[2][3] != ele[2][5];
    ele[2][3] != ele[2][6];
    ele[2][3] != ele[2][7];
    ele[2][3] != ele[2][8];
    ele[2][3] != ele[2][9];
    ele[2][3] != ele[20][3];
    ele[2][3] != ele[21][3];
    ele[2][3] != ele[22][3];
    ele[2][3] != ele[23][3];
    ele[2][3] != ele[24][3];
    ele[2][3] != ele[25][3];
    ele[2][3] != ele[26][3];
    ele[2][3] != ele[27][3];
    ele[2][3] != ele[28][3];
    ele[2][3] != ele[29][3];
    ele[2][3] != ele[3][0];
    ele[2][3] != ele[3][1];
    ele[2][3] != ele[3][2];
    ele[2][3] != ele[3][3];
    ele[2][3] != ele[3][4];
    ele[2][3] != ele[3][5];
    ele[2][3] != ele[30][3];
    ele[2][3] != ele[31][3];
    ele[2][3] != ele[32][3];
    ele[2][3] != ele[33][3];
    ele[2][3] != ele[34][3];
    ele[2][3] != ele[35][3];
    ele[2][3] != ele[4][0];
    ele[2][3] != ele[4][1];
    ele[2][3] != ele[4][2];
    ele[2][3] != ele[4][3];
    ele[2][3] != ele[4][4];
    ele[2][3] != ele[4][5];
    ele[2][3] != ele[5][0];
    ele[2][3] != ele[5][1];
    ele[2][3] != ele[5][2];
    ele[2][3] != ele[5][3];
    ele[2][3] != ele[5][4];
    ele[2][3] != ele[5][5];
    ele[2][3] != ele[6][3];
    ele[2][3] != ele[7][3];
    ele[2][3] != ele[8][3];
    ele[2][3] != ele[9][3];
    ele[2][30] != ele[10][30];
    ele[2][30] != ele[11][30];
    ele[2][30] != ele[12][30];
    ele[2][30] != ele[13][30];
    ele[2][30] != ele[14][30];
    ele[2][30] != ele[15][30];
    ele[2][30] != ele[16][30];
    ele[2][30] != ele[17][30];
    ele[2][30] != ele[18][30];
    ele[2][30] != ele[19][30];
    ele[2][30] != ele[2][31];
    ele[2][30] != ele[2][32];
    ele[2][30] != ele[2][33];
    ele[2][30] != ele[2][34];
    ele[2][30] != ele[2][35];
    ele[2][30] != ele[20][30];
    ele[2][30] != ele[21][30];
    ele[2][30] != ele[22][30];
    ele[2][30] != ele[23][30];
    ele[2][30] != ele[24][30];
    ele[2][30] != ele[25][30];
    ele[2][30] != ele[26][30];
    ele[2][30] != ele[27][30];
    ele[2][30] != ele[28][30];
    ele[2][30] != ele[29][30];
    ele[2][30] != ele[3][30];
    ele[2][30] != ele[3][31];
    ele[2][30] != ele[3][32];
    ele[2][30] != ele[3][33];
    ele[2][30] != ele[3][34];
    ele[2][30] != ele[3][35];
    ele[2][30] != ele[30][30];
    ele[2][30] != ele[31][30];
    ele[2][30] != ele[32][30];
    ele[2][30] != ele[33][30];
    ele[2][30] != ele[34][30];
    ele[2][30] != ele[35][30];
    ele[2][30] != ele[4][30];
    ele[2][30] != ele[4][31];
    ele[2][30] != ele[4][32];
    ele[2][30] != ele[4][33];
    ele[2][30] != ele[4][34];
    ele[2][30] != ele[4][35];
    ele[2][30] != ele[5][30];
    ele[2][30] != ele[5][31];
    ele[2][30] != ele[5][32];
    ele[2][30] != ele[5][33];
    ele[2][30] != ele[5][34];
    ele[2][30] != ele[5][35];
    ele[2][30] != ele[6][30];
    ele[2][30] != ele[7][30];
    ele[2][30] != ele[8][30];
    ele[2][30] != ele[9][30];
    ele[2][31] != ele[10][31];
    ele[2][31] != ele[11][31];
    ele[2][31] != ele[12][31];
    ele[2][31] != ele[13][31];
    ele[2][31] != ele[14][31];
    ele[2][31] != ele[15][31];
    ele[2][31] != ele[16][31];
    ele[2][31] != ele[17][31];
    ele[2][31] != ele[18][31];
    ele[2][31] != ele[19][31];
    ele[2][31] != ele[2][32];
    ele[2][31] != ele[2][33];
    ele[2][31] != ele[2][34];
    ele[2][31] != ele[2][35];
    ele[2][31] != ele[20][31];
    ele[2][31] != ele[21][31];
    ele[2][31] != ele[22][31];
    ele[2][31] != ele[23][31];
    ele[2][31] != ele[24][31];
    ele[2][31] != ele[25][31];
    ele[2][31] != ele[26][31];
    ele[2][31] != ele[27][31];
    ele[2][31] != ele[28][31];
    ele[2][31] != ele[29][31];
    ele[2][31] != ele[3][30];
    ele[2][31] != ele[3][31];
    ele[2][31] != ele[3][32];
    ele[2][31] != ele[3][33];
    ele[2][31] != ele[3][34];
    ele[2][31] != ele[3][35];
    ele[2][31] != ele[30][31];
    ele[2][31] != ele[31][31];
    ele[2][31] != ele[32][31];
    ele[2][31] != ele[33][31];
    ele[2][31] != ele[34][31];
    ele[2][31] != ele[35][31];
    ele[2][31] != ele[4][30];
    ele[2][31] != ele[4][31];
    ele[2][31] != ele[4][32];
    ele[2][31] != ele[4][33];
    ele[2][31] != ele[4][34];
    ele[2][31] != ele[4][35];
    ele[2][31] != ele[5][30];
    ele[2][31] != ele[5][31];
    ele[2][31] != ele[5][32];
    ele[2][31] != ele[5][33];
    ele[2][31] != ele[5][34];
    ele[2][31] != ele[5][35];
    ele[2][31] != ele[6][31];
    ele[2][31] != ele[7][31];
    ele[2][31] != ele[8][31];
    ele[2][31] != ele[9][31];
    ele[2][32] != ele[10][32];
    ele[2][32] != ele[11][32];
    ele[2][32] != ele[12][32];
    ele[2][32] != ele[13][32];
    ele[2][32] != ele[14][32];
    ele[2][32] != ele[15][32];
    ele[2][32] != ele[16][32];
    ele[2][32] != ele[17][32];
    ele[2][32] != ele[18][32];
    ele[2][32] != ele[19][32];
    ele[2][32] != ele[2][33];
    ele[2][32] != ele[2][34];
    ele[2][32] != ele[2][35];
    ele[2][32] != ele[20][32];
    ele[2][32] != ele[21][32];
    ele[2][32] != ele[22][32];
    ele[2][32] != ele[23][32];
    ele[2][32] != ele[24][32];
    ele[2][32] != ele[25][32];
    ele[2][32] != ele[26][32];
    ele[2][32] != ele[27][32];
    ele[2][32] != ele[28][32];
    ele[2][32] != ele[29][32];
    ele[2][32] != ele[3][30];
    ele[2][32] != ele[3][31];
    ele[2][32] != ele[3][32];
    ele[2][32] != ele[3][33];
    ele[2][32] != ele[3][34];
    ele[2][32] != ele[3][35];
    ele[2][32] != ele[30][32];
    ele[2][32] != ele[31][32];
    ele[2][32] != ele[32][32];
    ele[2][32] != ele[33][32];
    ele[2][32] != ele[34][32];
    ele[2][32] != ele[35][32];
    ele[2][32] != ele[4][30];
    ele[2][32] != ele[4][31];
    ele[2][32] != ele[4][32];
    ele[2][32] != ele[4][33];
    ele[2][32] != ele[4][34];
    ele[2][32] != ele[4][35];
    ele[2][32] != ele[5][30];
    ele[2][32] != ele[5][31];
    ele[2][32] != ele[5][32];
    ele[2][32] != ele[5][33];
    ele[2][32] != ele[5][34];
    ele[2][32] != ele[5][35];
    ele[2][32] != ele[6][32];
    ele[2][32] != ele[7][32];
    ele[2][32] != ele[8][32];
    ele[2][32] != ele[9][32];
    ele[2][33] != ele[10][33];
    ele[2][33] != ele[11][33];
    ele[2][33] != ele[12][33];
    ele[2][33] != ele[13][33];
    ele[2][33] != ele[14][33];
    ele[2][33] != ele[15][33];
    ele[2][33] != ele[16][33];
    ele[2][33] != ele[17][33];
    ele[2][33] != ele[18][33];
    ele[2][33] != ele[19][33];
    ele[2][33] != ele[2][34];
    ele[2][33] != ele[2][35];
    ele[2][33] != ele[20][33];
    ele[2][33] != ele[21][33];
    ele[2][33] != ele[22][33];
    ele[2][33] != ele[23][33];
    ele[2][33] != ele[24][33];
    ele[2][33] != ele[25][33];
    ele[2][33] != ele[26][33];
    ele[2][33] != ele[27][33];
    ele[2][33] != ele[28][33];
    ele[2][33] != ele[29][33];
    ele[2][33] != ele[3][30];
    ele[2][33] != ele[3][31];
    ele[2][33] != ele[3][32];
    ele[2][33] != ele[3][33];
    ele[2][33] != ele[3][34];
    ele[2][33] != ele[3][35];
    ele[2][33] != ele[30][33];
    ele[2][33] != ele[31][33];
    ele[2][33] != ele[32][33];
    ele[2][33] != ele[33][33];
    ele[2][33] != ele[34][33];
    ele[2][33] != ele[35][33];
    ele[2][33] != ele[4][30];
    ele[2][33] != ele[4][31];
    ele[2][33] != ele[4][32];
    ele[2][33] != ele[4][33];
    ele[2][33] != ele[4][34];
    ele[2][33] != ele[4][35];
    ele[2][33] != ele[5][30];
    ele[2][33] != ele[5][31];
    ele[2][33] != ele[5][32];
    ele[2][33] != ele[5][33];
    ele[2][33] != ele[5][34];
    ele[2][33] != ele[5][35];
    ele[2][33] != ele[6][33];
    ele[2][33] != ele[7][33];
    ele[2][33] != ele[8][33];
    ele[2][33] != ele[9][33];
    ele[2][34] != ele[10][34];
    ele[2][34] != ele[11][34];
    ele[2][34] != ele[12][34];
    ele[2][34] != ele[13][34];
    ele[2][34] != ele[14][34];
    ele[2][34] != ele[15][34];
    ele[2][34] != ele[16][34];
    ele[2][34] != ele[17][34];
    ele[2][34] != ele[18][34];
    ele[2][34] != ele[19][34];
    ele[2][34] != ele[2][35];
    ele[2][34] != ele[20][34];
    ele[2][34] != ele[21][34];
    ele[2][34] != ele[22][34];
    ele[2][34] != ele[23][34];
    ele[2][34] != ele[24][34];
    ele[2][34] != ele[25][34];
    ele[2][34] != ele[26][34];
    ele[2][34] != ele[27][34];
    ele[2][34] != ele[28][34];
    ele[2][34] != ele[29][34];
    ele[2][34] != ele[3][30];
    ele[2][34] != ele[3][31];
    ele[2][34] != ele[3][32];
    ele[2][34] != ele[3][33];
    ele[2][34] != ele[3][34];
    ele[2][34] != ele[3][35];
    ele[2][34] != ele[30][34];
    ele[2][34] != ele[31][34];
    ele[2][34] != ele[32][34];
    ele[2][34] != ele[33][34];
    ele[2][34] != ele[34][34];
    ele[2][34] != ele[35][34];
    ele[2][34] != ele[4][30];
    ele[2][34] != ele[4][31];
    ele[2][34] != ele[4][32];
    ele[2][34] != ele[4][33];
    ele[2][34] != ele[4][34];
    ele[2][34] != ele[4][35];
    ele[2][34] != ele[5][30];
    ele[2][34] != ele[5][31];
    ele[2][34] != ele[5][32];
    ele[2][34] != ele[5][33];
    ele[2][34] != ele[5][34];
    ele[2][34] != ele[5][35];
    ele[2][34] != ele[6][34];
    ele[2][34] != ele[7][34];
    ele[2][34] != ele[8][34];
    ele[2][34] != ele[9][34];
    ele[2][35] != ele[10][35];
    ele[2][35] != ele[11][35];
    ele[2][35] != ele[12][35];
    ele[2][35] != ele[13][35];
    ele[2][35] != ele[14][35];
    ele[2][35] != ele[15][35];
    ele[2][35] != ele[16][35];
    ele[2][35] != ele[17][35];
    ele[2][35] != ele[18][35];
    ele[2][35] != ele[19][35];
    ele[2][35] != ele[20][35];
    ele[2][35] != ele[21][35];
    ele[2][35] != ele[22][35];
    ele[2][35] != ele[23][35];
    ele[2][35] != ele[24][35];
    ele[2][35] != ele[25][35];
    ele[2][35] != ele[26][35];
    ele[2][35] != ele[27][35];
    ele[2][35] != ele[28][35];
    ele[2][35] != ele[29][35];
    ele[2][35] != ele[3][30];
    ele[2][35] != ele[3][31];
    ele[2][35] != ele[3][32];
    ele[2][35] != ele[3][33];
    ele[2][35] != ele[3][34];
    ele[2][35] != ele[3][35];
    ele[2][35] != ele[30][35];
    ele[2][35] != ele[31][35];
    ele[2][35] != ele[32][35];
    ele[2][35] != ele[33][35];
    ele[2][35] != ele[34][35];
    ele[2][35] != ele[35][35];
    ele[2][35] != ele[4][30];
    ele[2][35] != ele[4][31];
    ele[2][35] != ele[4][32];
    ele[2][35] != ele[4][33];
    ele[2][35] != ele[4][34];
    ele[2][35] != ele[4][35];
    ele[2][35] != ele[5][30];
    ele[2][35] != ele[5][31];
    ele[2][35] != ele[5][32];
    ele[2][35] != ele[5][33];
    ele[2][35] != ele[5][34];
    ele[2][35] != ele[5][35];
    ele[2][35] != ele[6][35];
    ele[2][35] != ele[7][35];
    ele[2][35] != ele[8][35];
    ele[2][35] != ele[9][35];
    ele[2][4] != ele[10][4];
    ele[2][4] != ele[11][4];
    ele[2][4] != ele[12][4];
    ele[2][4] != ele[13][4];
    ele[2][4] != ele[14][4];
    ele[2][4] != ele[15][4];
    ele[2][4] != ele[16][4];
    ele[2][4] != ele[17][4];
    ele[2][4] != ele[18][4];
    ele[2][4] != ele[19][4];
    ele[2][4] != ele[2][10];
    ele[2][4] != ele[2][11];
    ele[2][4] != ele[2][12];
    ele[2][4] != ele[2][13];
    ele[2][4] != ele[2][14];
    ele[2][4] != ele[2][15];
    ele[2][4] != ele[2][16];
    ele[2][4] != ele[2][17];
    ele[2][4] != ele[2][18];
    ele[2][4] != ele[2][19];
    ele[2][4] != ele[2][20];
    ele[2][4] != ele[2][21];
    ele[2][4] != ele[2][22];
    ele[2][4] != ele[2][23];
    ele[2][4] != ele[2][24];
    ele[2][4] != ele[2][25];
    ele[2][4] != ele[2][26];
    ele[2][4] != ele[2][27];
    ele[2][4] != ele[2][28];
    ele[2][4] != ele[2][29];
    ele[2][4] != ele[2][30];
    ele[2][4] != ele[2][31];
    ele[2][4] != ele[2][32];
    ele[2][4] != ele[2][33];
    ele[2][4] != ele[2][34];
    ele[2][4] != ele[2][35];
    ele[2][4] != ele[2][5];
    ele[2][4] != ele[2][6];
    ele[2][4] != ele[2][7];
    ele[2][4] != ele[2][8];
    ele[2][4] != ele[2][9];
    ele[2][4] != ele[20][4];
    ele[2][4] != ele[21][4];
    ele[2][4] != ele[22][4];
    ele[2][4] != ele[23][4];
    ele[2][4] != ele[24][4];
    ele[2][4] != ele[25][4];
    ele[2][4] != ele[26][4];
    ele[2][4] != ele[27][4];
    ele[2][4] != ele[28][4];
    ele[2][4] != ele[29][4];
    ele[2][4] != ele[3][0];
    ele[2][4] != ele[3][1];
    ele[2][4] != ele[3][2];
    ele[2][4] != ele[3][3];
    ele[2][4] != ele[3][4];
    ele[2][4] != ele[3][5];
    ele[2][4] != ele[30][4];
    ele[2][4] != ele[31][4];
    ele[2][4] != ele[32][4];
    ele[2][4] != ele[33][4];
    ele[2][4] != ele[34][4];
    ele[2][4] != ele[35][4];
    ele[2][4] != ele[4][0];
    ele[2][4] != ele[4][1];
    ele[2][4] != ele[4][2];
    ele[2][4] != ele[4][3];
    ele[2][4] != ele[4][4];
    ele[2][4] != ele[4][5];
    ele[2][4] != ele[5][0];
    ele[2][4] != ele[5][1];
    ele[2][4] != ele[5][2];
    ele[2][4] != ele[5][3];
    ele[2][4] != ele[5][4];
    ele[2][4] != ele[5][5];
    ele[2][4] != ele[6][4];
    ele[2][4] != ele[7][4];
    ele[2][4] != ele[8][4];
    ele[2][4] != ele[9][4];
    ele[2][5] != ele[10][5];
    ele[2][5] != ele[11][5];
    ele[2][5] != ele[12][5];
    ele[2][5] != ele[13][5];
    ele[2][5] != ele[14][5];
    ele[2][5] != ele[15][5];
    ele[2][5] != ele[16][5];
    ele[2][5] != ele[17][5];
    ele[2][5] != ele[18][5];
    ele[2][5] != ele[19][5];
    ele[2][5] != ele[2][10];
    ele[2][5] != ele[2][11];
    ele[2][5] != ele[2][12];
    ele[2][5] != ele[2][13];
    ele[2][5] != ele[2][14];
    ele[2][5] != ele[2][15];
    ele[2][5] != ele[2][16];
    ele[2][5] != ele[2][17];
    ele[2][5] != ele[2][18];
    ele[2][5] != ele[2][19];
    ele[2][5] != ele[2][20];
    ele[2][5] != ele[2][21];
    ele[2][5] != ele[2][22];
    ele[2][5] != ele[2][23];
    ele[2][5] != ele[2][24];
    ele[2][5] != ele[2][25];
    ele[2][5] != ele[2][26];
    ele[2][5] != ele[2][27];
    ele[2][5] != ele[2][28];
    ele[2][5] != ele[2][29];
    ele[2][5] != ele[2][30];
    ele[2][5] != ele[2][31];
    ele[2][5] != ele[2][32];
    ele[2][5] != ele[2][33];
    ele[2][5] != ele[2][34];
    ele[2][5] != ele[2][35];
    ele[2][5] != ele[2][6];
    ele[2][5] != ele[2][7];
    ele[2][5] != ele[2][8];
    ele[2][5] != ele[2][9];
    ele[2][5] != ele[20][5];
    ele[2][5] != ele[21][5];
    ele[2][5] != ele[22][5];
    ele[2][5] != ele[23][5];
    ele[2][5] != ele[24][5];
    ele[2][5] != ele[25][5];
    ele[2][5] != ele[26][5];
    ele[2][5] != ele[27][5];
    ele[2][5] != ele[28][5];
    ele[2][5] != ele[29][5];
    ele[2][5] != ele[3][0];
    ele[2][5] != ele[3][1];
    ele[2][5] != ele[3][2];
    ele[2][5] != ele[3][3];
    ele[2][5] != ele[3][4];
    ele[2][5] != ele[3][5];
    ele[2][5] != ele[30][5];
    ele[2][5] != ele[31][5];
    ele[2][5] != ele[32][5];
    ele[2][5] != ele[33][5];
    ele[2][5] != ele[34][5];
    ele[2][5] != ele[35][5];
    ele[2][5] != ele[4][0];
    ele[2][5] != ele[4][1];
    ele[2][5] != ele[4][2];
    ele[2][5] != ele[4][3];
    ele[2][5] != ele[4][4];
    ele[2][5] != ele[4][5];
    ele[2][5] != ele[5][0];
    ele[2][5] != ele[5][1];
    ele[2][5] != ele[5][2];
    ele[2][5] != ele[5][3];
    ele[2][5] != ele[5][4];
    ele[2][5] != ele[5][5];
    ele[2][5] != ele[6][5];
    ele[2][5] != ele[7][5];
    ele[2][5] != ele[8][5];
    ele[2][5] != ele[9][5];
    ele[2][6] != ele[10][6];
    ele[2][6] != ele[11][6];
    ele[2][6] != ele[12][6];
    ele[2][6] != ele[13][6];
    ele[2][6] != ele[14][6];
    ele[2][6] != ele[15][6];
    ele[2][6] != ele[16][6];
    ele[2][6] != ele[17][6];
    ele[2][6] != ele[18][6];
    ele[2][6] != ele[19][6];
    ele[2][6] != ele[2][10];
    ele[2][6] != ele[2][11];
    ele[2][6] != ele[2][12];
    ele[2][6] != ele[2][13];
    ele[2][6] != ele[2][14];
    ele[2][6] != ele[2][15];
    ele[2][6] != ele[2][16];
    ele[2][6] != ele[2][17];
    ele[2][6] != ele[2][18];
    ele[2][6] != ele[2][19];
    ele[2][6] != ele[2][20];
    ele[2][6] != ele[2][21];
    ele[2][6] != ele[2][22];
    ele[2][6] != ele[2][23];
    ele[2][6] != ele[2][24];
    ele[2][6] != ele[2][25];
    ele[2][6] != ele[2][26];
    ele[2][6] != ele[2][27];
    ele[2][6] != ele[2][28];
    ele[2][6] != ele[2][29];
    ele[2][6] != ele[2][30];
    ele[2][6] != ele[2][31];
    ele[2][6] != ele[2][32];
    ele[2][6] != ele[2][33];
    ele[2][6] != ele[2][34];
    ele[2][6] != ele[2][35];
    ele[2][6] != ele[2][7];
    ele[2][6] != ele[2][8];
    ele[2][6] != ele[2][9];
    ele[2][6] != ele[20][6];
    ele[2][6] != ele[21][6];
    ele[2][6] != ele[22][6];
    ele[2][6] != ele[23][6];
    ele[2][6] != ele[24][6];
    ele[2][6] != ele[25][6];
    ele[2][6] != ele[26][6];
    ele[2][6] != ele[27][6];
    ele[2][6] != ele[28][6];
    ele[2][6] != ele[29][6];
    ele[2][6] != ele[3][10];
    ele[2][6] != ele[3][11];
    ele[2][6] != ele[3][6];
    ele[2][6] != ele[3][7];
    ele[2][6] != ele[3][8];
    ele[2][6] != ele[3][9];
    ele[2][6] != ele[30][6];
    ele[2][6] != ele[31][6];
    ele[2][6] != ele[32][6];
    ele[2][6] != ele[33][6];
    ele[2][6] != ele[34][6];
    ele[2][6] != ele[35][6];
    ele[2][6] != ele[4][10];
    ele[2][6] != ele[4][11];
    ele[2][6] != ele[4][6];
    ele[2][6] != ele[4][7];
    ele[2][6] != ele[4][8];
    ele[2][6] != ele[4][9];
    ele[2][6] != ele[5][10];
    ele[2][6] != ele[5][11];
    ele[2][6] != ele[5][6];
    ele[2][6] != ele[5][7];
    ele[2][6] != ele[5][8];
    ele[2][6] != ele[5][9];
    ele[2][6] != ele[6][6];
    ele[2][6] != ele[7][6];
    ele[2][6] != ele[8][6];
    ele[2][6] != ele[9][6];
    ele[2][7] != ele[10][7];
    ele[2][7] != ele[11][7];
    ele[2][7] != ele[12][7];
    ele[2][7] != ele[13][7];
    ele[2][7] != ele[14][7];
    ele[2][7] != ele[15][7];
    ele[2][7] != ele[16][7];
    ele[2][7] != ele[17][7];
    ele[2][7] != ele[18][7];
    ele[2][7] != ele[19][7];
    ele[2][7] != ele[2][10];
    ele[2][7] != ele[2][11];
    ele[2][7] != ele[2][12];
    ele[2][7] != ele[2][13];
    ele[2][7] != ele[2][14];
    ele[2][7] != ele[2][15];
    ele[2][7] != ele[2][16];
    ele[2][7] != ele[2][17];
    ele[2][7] != ele[2][18];
    ele[2][7] != ele[2][19];
    ele[2][7] != ele[2][20];
    ele[2][7] != ele[2][21];
    ele[2][7] != ele[2][22];
    ele[2][7] != ele[2][23];
    ele[2][7] != ele[2][24];
    ele[2][7] != ele[2][25];
    ele[2][7] != ele[2][26];
    ele[2][7] != ele[2][27];
    ele[2][7] != ele[2][28];
    ele[2][7] != ele[2][29];
    ele[2][7] != ele[2][30];
    ele[2][7] != ele[2][31];
    ele[2][7] != ele[2][32];
    ele[2][7] != ele[2][33];
    ele[2][7] != ele[2][34];
    ele[2][7] != ele[2][35];
    ele[2][7] != ele[2][8];
    ele[2][7] != ele[2][9];
    ele[2][7] != ele[20][7];
    ele[2][7] != ele[21][7];
    ele[2][7] != ele[22][7];
    ele[2][7] != ele[23][7];
    ele[2][7] != ele[24][7];
    ele[2][7] != ele[25][7];
    ele[2][7] != ele[26][7];
    ele[2][7] != ele[27][7];
    ele[2][7] != ele[28][7];
    ele[2][7] != ele[29][7];
    ele[2][7] != ele[3][10];
    ele[2][7] != ele[3][11];
    ele[2][7] != ele[3][6];
    ele[2][7] != ele[3][7];
    ele[2][7] != ele[3][8];
    ele[2][7] != ele[3][9];
    ele[2][7] != ele[30][7];
    ele[2][7] != ele[31][7];
    ele[2][7] != ele[32][7];
    ele[2][7] != ele[33][7];
    ele[2][7] != ele[34][7];
    ele[2][7] != ele[35][7];
    ele[2][7] != ele[4][10];
    ele[2][7] != ele[4][11];
    ele[2][7] != ele[4][6];
    ele[2][7] != ele[4][7];
    ele[2][7] != ele[4][8];
    ele[2][7] != ele[4][9];
    ele[2][7] != ele[5][10];
    ele[2][7] != ele[5][11];
    ele[2][7] != ele[5][6];
    ele[2][7] != ele[5][7];
    ele[2][7] != ele[5][8];
    ele[2][7] != ele[5][9];
    ele[2][7] != ele[6][7];
    ele[2][7] != ele[7][7];
    ele[2][7] != ele[8][7];
    ele[2][7] != ele[9][7];
    ele[2][8] != ele[10][8];
    ele[2][8] != ele[11][8];
    ele[2][8] != ele[12][8];
    ele[2][8] != ele[13][8];
    ele[2][8] != ele[14][8];
    ele[2][8] != ele[15][8];
    ele[2][8] != ele[16][8];
    ele[2][8] != ele[17][8];
    ele[2][8] != ele[18][8];
    ele[2][8] != ele[19][8];
    ele[2][8] != ele[2][10];
    ele[2][8] != ele[2][11];
    ele[2][8] != ele[2][12];
    ele[2][8] != ele[2][13];
    ele[2][8] != ele[2][14];
    ele[2][8] != ele[2][15];
    ele[2][8] != ele[2][16];
    ele[2][8] != ele[2][17];
    ele[2][8] != ele[2][18];
    ele[2][8] != ele[2][19];
    ele[2][8] != ele[2][20];
    ele[2][8] != ele[2][21];
    ele[2][8] != ele[2][22];
    ele[2][8] != ele[2][23];
    ele[2][8] != ele[2][24];
    ele[2][8] != ele[2][25];
    ele[2][8] != ele[2][26];
    ele[2][8] != ele[2][27];
    ele[2][8] != ele[2][28];
    ele[2][8] != ele[2][29];
    ele[2][8] != ele[2][30];
    ele[2][8] != ele[2][31];
    ele[2][8] != ele[2][32];
    ele[2][8] != ele[2][33];
    ele[2][8] != ele[2][34];
    ele[2][8] != ele[2][35];
    ele[2][8] != ele[2][9];
    ele[2][8] != ele[20][8];
    ele[2][8] != ele[21][8];
    ele[2][8] != ele[22][8];
    ele[2][8] != ele[23][8];
    ele[2][8] != ele[24][8];
    ele[2][8] != ele[25][8];
    ele[2][8] != ele[26][8];
    ele[2][8] != ele[27][8];
    ele[2][8] != ele[28][8];
    ele[2][8] != ele[29][8];
    ele[2][8] != ele[3][10];
    ele[2][8] != ele[3][11];
    ele[2][8] != ele[3][6];
    ele[2][8] != ele[3][7];
    ele[2][8] != ele[3][8];
    ele[2][8] != ele[3][9];
    ele[2][8] != ele[30][8];
    ele[2][8] != ele[31][8];
    ele[2][8] != ele[32][8];
    ele[2][8] != ele[33][8];
    ele[2][8] != ele[34][8];
    ele[2][8] != ele[35][8];
    ele[2][8] != ele[4][10];
    ele[2][8] != ele[4][11];
    ele[2][8] != ele[4][6];
    ele[2][8] != ele[4][7];
    ele[2][8] != ele[4][8];
    ele[2][8] != ele[4][9];
    ele[2][8] != ele[5][10];
    ele[2][8] != ele[5][11];
    ele[2][8] != ele[5][6];
    ele[2][8] != ele[5][7];
    ele[2][8] != ele[5][8];
    ele[2][8] != ele[5][9];
    ele[2][8] != ele[6][8];
    ele[2][8] != ele[7][8];
    ele[2][8] != ele[8][8];
    ele[2][8] != ele[9][8];
    ele[2][9] != ele[10][9];
    ele[2][9] != ele[11][9];
    ele[2][9] != ele[12][9];
    ele[2][9] != ele[13][9];
    ele[2][9] != ele[14][9];
    ele[2][9] != ele[15][9];
    ele[2][9] != ele[16][9];
    ele[2][9] != ele[17][9];
    ele[2][9] != ele[18][9];
    ele[2][9] != ele[19][9];
    ele[2][9] != ele[2][10];
    ele[2][9] != ele[2][11];
    ele[2][9] != ele[2][12];
    ele[2][9] != ele[2][13];
    ele[2][9] != ele[2][14];
    ele[2][9] != ele[2][15];
    ele[2][9] != ele[2][16];
    ele[2][9] != ele[2][17];
    ele[2][9] != ele[2][18];
    ele[2][9] != ele[2][19];
    ele[2][9] != ele[2][20];
    ele[2][9] != ele[2][21];
    ele[2][9] != ele[2][22];
    ele[2][9] != ele[2][23];
    ele[2][9] != ele[2][24];
    ele[2][9] != ele[2][25];
    ele[2][9] != ele[2][26];
    ele[2][9] != ele[2][27];
    ele[2][9] != ele[2][28];
    ele[2][9] != ele[2][29];
    ele[2][9] != ele[2][30];
    ele[2][9] != ele[2][31];
    ele[2][9] != ele[2][32];
    ele[2][9] != ele[2][33];
    ele[2][9] != ele[2][34];
    ele[2][9] != ele[2][35];
    ele[2][9] != ele[20][9];
    ele[2][9] != ele[21][9];
    ele[2][9] != ele[22][9];
    ele[2][9] != ele[23][9];
    ele[2][9] != ele[24][9];
    ele[2][9] != ele[25][9];
    ele[2][9] != ele[26][9];
    ele[2][9] != ele[27][9];
    ele[2][9] != ele[28][9];
    ele[2][9] != ele[29][9];
    ele[2][9] != ele[3][10];
    ele[2][9] != ele[3][11];
    ele[2][9] != ele[3][6];
    ele[2][9] != ele[3][7];
    ele[2][9] != ele[3][8];
    ele[2][9] != ele[3][9];
    ele[2][9] != ele[30][9];
    ele[2][9] != ele[31][9];
    ele[2][9] != ele[32][9];
    ele[2][9] != ele[33][9];
    ele[2][9] != ele[34][9];
    ele[2][9] != ele[35][9];
    ele[2][9] != ele[4][10];
    ele[2][9] != ele[4][11];
    ele[2][9] != ele[4][6];
    ele[2][9] != ele[4][7];
    ele[2][9] != ele[4][8];
    ele[2][9] != ele[4][9];
    ele[2][9] != ele[5][10];
    ele[2][9] != ele[5][11];
    ele[2][9] != ele[5][6];
    ele[2][9] != ele[5][7];
    ele[2][9] != ele[5][8];
    ele[2][9] != ele[5][9];
    ele[2][9] != ele[6][9];
    ele[2][9] != ele[7][9];
    ele[2][9] != ele[8][9];
    ele[2][9] != ele[9][9];
    ele[20][0] != ele[20][1];
    ele[20][0] != ele[20][10];
    ele[20][0] != ele[20][11];
    ele[20][0] != ele[20][12];
    ele[20][0] != ele[20][13];
    ele[20][0] != ele[20][14];
    ele[20][0] != ele[20][15];
    ele[20][0] != ele[20][16];
    ele[20][0] != ele[20][17];
    ele[20][0] != ele[20][18];
    ele[20][0] != ele[20][19];
    ele[20][0] != ele[20][2];
    ele[20][0] != ele[20][20];
    ele[20][0] != ele[20][21];
    ele[20][0] != ele[20][22];
    ele[20][0] != ele[20][23];
    ele[20][0] != ele[20][24];
    ele[20][0] != ele[20][25];
    ele[20][0] != ele[20][26];
    ele[20][0] != ele[20][27];
    ele[20][0] != ele[20][28];
    ele[20][0] != ele[20][29];
    ele[20][0] != ele[20][3];
    ele[20][0] != ele[20][30];
    ele[20][0] != ele[20][31];
    ele[20][0] != ele[20][32];
    ele[20][0] != ele[20][33];
    ele[20][0] != ele[20][34];
    ele[20][0] != ele[20][35];
    ele[20][0] != ele[20][4];
    ele[20][0] != ele[20][5];
    ele[20][0] != ele[20][6];
    ele[20][0] != ele[20][7];
    ele[20][0] != ele[20][8];
    ele[20][0] != ele[20][9];
    ele[20][0] != ele[21][0];
    ele[20][0] != ele[21][1];
    ele[20][0] != ele[21][2];
    ele[20][0] != ele[21][3];
    ele[20][0] != ele[21][4];
    ele[20][0] != ele[21][5];
    ele[20][0] != ele[22][0];
    ele[20][0] != ele[22][1];
    ele[20][0] != ele[22][2];
    ele[20][0] != ele[22][3];
    ele[20][0] != ele[22][4];
    ele[20][0] != ele[22][5];
    ele[20][0] != ele[23][0];
    ele[20][0] != ele[23][1];
    ele[20][0] != ele[23][2];
    ele[20][0] != ele[23][3];
    ele[20][0] != ele[23][4];
    ele[20][0] != ele[23][5];
    ele[20][0] != ele[24][0];
    ele[20][0] != ele[25][0];
    ele[20][0] != ele[26][0];
    ele[20][0] != ele[27][0];
    ele[20][0] != ele[28][0];
    ele[20][0] != ele[29][0];
    ele[20][0] != ele[30][0];
    ele[20][0] != ele[31][0];
    ele[20][0] != ele[32][0];
    ele[20][0] != ele[33][0];
    ele[20][0] != ele[34][0];
    ele[20][0] != ele[35][0];
    ele[20][1] != ele[20][10];
    ele[20][1] != ele[20][11];
    ele[20][1] != ele[20][12];
    ele[20][1] != ele[20][13];
    ele[20][1] != ele[20][14];
    ele[20][1] != ele[20][15];
    ele[20][1] != ele[20][16];
    ele[20][1] != ele[20][17];
    ele[20][1] != ele[20][18];
    ele[20][1] != ele[20][19];
    ele[20][1] != ele[20][2];
    ele[20][1] != ele[20][20];
    ele[20][1] != ele[20][21];
    ele[20][1] != ele[20][22];
    ele[20][1] != ele[20][23];
    ele[20][1] != ele[20][24];
    ele[20][1] != ele[20][25];
    ele[20][1] != ele[20][26];
    ele[20][1] != ele[20][27];
    ele[20][1] != ele[20][28];
    ele[20][1] != ele[20][29];
    ele[20][1] != ele[20][3];
    ele[20][1] != ele[20][30];
    ele[20][1] != ele[20][31];
    ele[20][1] != ele[20][32];
    ele[20][1] != ele[20][33];
    ele[20][1] != ele[20][34];
    ele[20][1] != ele[20][35];
    ele[20][1] != ele[20][4];
    ele[20][1] != ele[20][5];
    ele[20][1] != ele[20][6];
    ele[20][1] != ele[20][7];
    ele[20][1] != ele[20][8];
    ele[20][1] != ele[20][9];
    ele[20][1] != ele[21][0];
    ele[20][1] != ele[21][1];
    ele[20][1] != ele[21][2];
    ele[20][1] != ele[21][3];
    ele[20][1] != ele[21][4];
    ele[20][1] != ele[21][5];
    ele[20][1] != ele[22][0];
    ele[20][1] != ele[22][1];
    ele[20][1] != ele[22][2];
    ele[20][1] != ele[22][3];
    ele[20][1] != ele[22][4];
    ele[20][1] != ele[22][5];
    ele[20][1] != ele[23][0];
    ele[20][1] != ele[23][1];
    ele[20][1] != ele[23][2];
    ele[20][1] != ele[23][3];
    ele[20][1] != ele[23][4];
    ele[20][1] != ele[23][5];
    ele[20][1] != ele[24][1];
    ele[20][1] != ele[25][1];
    ele[20][1] != ele[26][1];
    ele[20][1] != ele[27][1];
    ele[20][1] != ele[28][1];
    ele[20][1] != ele[29][1];
    ele[20][1] != ele[30][1];
    ele[20][1] != ele[31][1];
    ele[20][1] != ele[32][1];
    ele[20][1] != ele[33][1];
    ele[20][1] != ele[34][1];
    ele[20][1] != ele[35][1];
    ele[20][10] != ele[20][11];
    ele[20][10] != ele[20][12];
    ele[20][10] != ele[20][13];
    ele[20][10] != ele[20][14];
    ele[20][10] != ele[20][15];
    ele[20][10] != ele[20][16];
    ele[20][10] != ele[20][17];
    ele[20][10] != ele[20][18];
    ele[20][10] != ele[20][19];
    ele[20][10] != ele[20][20];
    ele[20][10] != ele[20][21];
    ele[20][10] != ele[20][22];
    ele[20][10] != ele[20][23];
    ele[20][10] != ele[20][24];
    ele[20][10] != ele[20][25];
    ele[20][10] != ele[20][26];
    ele[20][10] != ele[20][27];
    ele[20][10] != ele[20][28];
    ele[20][10] != ele[20][29];
    ele[20][10] != ele[20][30];
    ele[20][10] != ele[20][31];
    ele[20][10] != ele[20][32];
    ele[20][10] != ele[20][33];
    ele[20][10] != ele[20][34];
    ele[20][10] != ele[20][35];
    ele[20][10] != ele[21][10];
    ele[20][10] != ele[21][11];
    ele[20][10] != ele[21][6];
    ele[20][10] != ele[21][7];
    ele[20][10] != ele[21][8];
    ele[20][10] != ele[21][9];
    ele[20][10] != ele[22][10];
    ele[20][10] != ele[22][11];
    ele[20][10] != ele[22][6];
    ele[20][10] != ele[22][7];
    ele[20][10] != ele[22][8];
    ele[20][10] != ele[22][9];
    ele[20][10] != ele[23][10];
    ele[20][10] != ele[23][11];
    ele[20][10] != ele[23][6];
    ele[20][10] != ele[23][7];
    ele[20][10] != ele[23][8];
    ele[20][10] != ele[23][9];
    ele[20][10] != ele[24][10];
    ele[20][10] != ele[25][10];
    ele[20][10] != ele[26][10];
    ele[20][10] != ele[27][10];
    ele[20][10] != ele[28][10];
    ele[20][10] != ele[29][10];
    ele[20][10] != ele[30][10];
    ele[20][10] != ele[31][10];
    ele[20][10] != ele[32][10];
    ele[20][10] != ele[33][10];
    ele[20][10] != ele[34][10];
    ele[20][10] != ele[35][10];
    ele[20][11] != ele[20][12];
    ele[20][11] != ele[20][13];
    ele[20][11] != ele[20][14];
    ele[20][11] != ele[20][15];
    ele[20][11] != ele[20][16];
    ele[20][11] != ele[20][17];
    ele[20][11] != ele[20][18];
    ele[20][11] != ele[20][19];
    ele[20][11] != ele[20][20];
    ele[20][11] != ele[20][21];
    ele[20][11] != ele[20][22];
    ele[20][11] != ele[20][23];
    ele[20][11] != ele[20][24];
    ele[20][11] != ele[20][25];
    ele[20][11] != ele[20][26];
    ele[20][11] != ele[20][27];
    ele[20][11] != ele[20][28];
    ele[20][11] != ele[20][29];
    ele[20][11] != ele[20][30];
    ele[20][11] != ele[20][31];
    ele[20][11] != ele[20][32];
    ele[20][11] != ele[20][33];
    ele[20][11] != ele[20][34];
    ele[20][11] != ele[20][35];
    ele[20][11] != ele[21][10];
    ele[20][11] != ele[21][11];
    ele[20][11] != ele[21][6];
    ele[20][11] != ele[21][7];
    ele[20][11] != ele[21][8];
    ele[20][11] != ele[21][9];
    ele[20][11] != ele[22][10];
    ele[20][11] != ele[22][11];
    ele[20][11] != ele[22][6];
    ele[20][11] != ele[22][7];
    ele[20][11] != ele[22][8];
    ele[20][11] != ele[22][9];
    ele[20][11] != ele[23][10];
    ele[20][11] != ele[23][11];
    ele[20][11] != ele[23][6];
    ele[20][11] != ele[23][7];
    ele[20][11] != ele[23][8];
    ele[20][11] != ele[23][9];
    ele[20][11] != ele[24][11];
    ele[20][11] != ele[25][11];
    ele[20][11] != ele[26][11];
    ele[20][11] != ele[27][11];
    ele[20][11] != ele[28][11];
    ele[20][11] != ele[29][11];
    ele[20][11] != ele[30][11];
    ele[20][11] != ele[31][11];
    ele[20][11] != ele[32][11];
    ele[20][11] != ele[33][11];
    ele[20][11] != ele[34][11];
    ele[20][11] != ele[35][11];
    ele[20][12] != ele[20][13];
    ele[20][12] != ele[20][14];
    ele[20][12] != ele[20][15];
    ele[20][12] != ele[20][16];
    ele[20][12] != ele[20][17];
    ele[20][12] != ele[20][18];
    ele[20][12] != ele[20][19];
    ele[20][12] != ele[20][20];
    ele[20][12] != ele[20][21];
    ele[20][12] != ele[20][22];
    ele[20][12] != ele[20][23];
    ele[20][12] != ele[20][24];
    ele[20][12] != ele[20][25];
    ele[20][12] != ele[20][26];
    ele[20][12] != ele[20][27];
    ele[20][12] != ele[20][28];
    ele[20][12] != ele[20][29];
    ele[20][12] != ele[20][30];
    ele[20][12] != ele[20][31];
    ele[20][12] != ele[20][32];
    ele[20][12] != ele[20][33];
    ele[20][12] != ele[20][34];
    ele[20][12] != ele[20][35];
    ele[20][12] != ele[21][12];
    ele[20][12] != ele[21][13];
    ele[20][12] != ele[21][14];
    ele[20][12] != ele[21][15];
    ele[20][12] != ele[21][16];
    ele[20][12] != ele[21][17];
    ele[20][12] != ele[22][12];
    ele[20][12] != ele[22][13];
    ele[20][12] != ele[22][14];
    ele[20][12] != ele[22][15];
    ele[20][12] != ele[22][16];
    ele[20][12] != ele[22][17];
    ele[20][12] != ele[23][12];
    ele[20][12] != ele[23][13];
    ele[20][12] != ele[23][14];
    ele[20][12] != ele[23][15];
    ele[20][12] != ele[23][16];
    ele[20][12] != ele[23][17];
    ele[20][12] != ele[24][12];
    ele[20][12] != ele[25][12];
    ele[20][12] != ele[26][12];
    ele[20][12] != ele[27][12];
    ele[20][12] != ele[28][12];
    ele[20][12] != ele[29][12];
    ele[20][12] != ele[30][12];
    ele[20][12] != ele[31][12];
    ele[20][12] != ele[32][12];
    ele[20][12] != ele[33][12];
    ele[20][12] != ele[34][12];
    ele[20][12] != ele[35][12];
    ele[20][13] != ele[20][14];
    ele[20][13] != ele[20][15];
    ele[20][13] != ele[20][16];
    ele[20][13] != ele[20][17];
    ele[20][13] != ele[20][18];
    ele[20][13] != ele[20][19];
    ele[20][13] != ele[20][20];
    ele[20][13] != ele[20][21];
    ele[20][13] != ele[20][22];
    ele[20][13] != ele[20][23];
    ele[20][13] != ele[20][24];
    ele[20][13] != ele[20][25];
    ele[20][13] != ele[20][26];
    ele[20][13] != ele[20][27];
    ele[20][13] != ele[20][28];
    ele[20][13] != ele[20][29];
    ele[20][13] != ele[20][30];
    ele[20][13] != ele[20][31];
    ele[20][13] != ele[20][32];
    ele[20][13] != ele[20][33];
    ele[20][13] != ele[20][34];
    ele[20][13] != ele[20][35];
    ele[20][13] != ele[21][12];
    ele[20][13] != ele[21][13];
    ele[20][13] != ele[21][14];
    ele[20][13] != ele[21][15];
    ele[20][13] != ele[21][16];
    ele[20][13] != ele[21][17];
    ele[20][13] != ele[22][12];
    ele[20][13] != ele[22][13];
    ele[20][13] != ele[22][14];
    ele[20][13] != ele[22][15];
    ele[20][13] != ele[22][16];
    ele[20][13] != ele[22][17];
    ele[20][13] != ele[23][12];
    ele[20][13] != ele[23][13];
    ele[20][13] != ele[23][14];
    ele[20][13] != ele[23][15];
    ele[20][13] != ele[23][16];
    ele[20][13] != ele[23][17];
    ele[20][13] != ele[24][13];
    ele[20][13] != ele[25][13];
    ele[20][13] != ele[26][13];
    ele[20][13] != ele[27][13];
    ele[20][13] != ele[28][13];
    ele[20][13] != ele[29][13];
    ele[20][13] != ele[30][13];
    ele[20][13] != ele[31][13];
    ele[20][13] != ele[32][13];
    ele[20][13] != ele[33][13];
    ele[20][13] != ele[34][13];
    ele[20][13] != ele[35][13];
    ele[20][14] != ele[20][15];
    ele[20][14] != ele[20][16];
    ele[20][14] != ele[20][17];
    ele[20][14] != ele[20][18];
    ele[20][14] != ele[20][19];
    ele[20][14] != ele[20][20];
    ele[20][14] != ele[20][21];
    ele[20][14] != ele[20][22];
    ele[20][14] != ele[20][23];
    ele[20][14] != ele[20][24];
    ele[20][14] != ele[20][25];
    ele[20][14] != ele[20][26];
    ele[20][14] != ele[20][27];
    ele[20][14] != ele[20][28];
    ele[20][14] != ele[20][29];
    ele[20][14] != ele[20][30];
    ele[20][14] != ele[20][31];
    ele[20][14] != ele[20][32];
    ele[20][14] != ele[20][33];
    ele[20][14] != ele[20][34];
    ele[20][14] != ele[20][35];
    ele[20][14] != ele[21][12];
    ele[20][14] != ele[21][13];
    ele[20][14] != ele[21][14];
    ele[20][14] != ele[21][15];
    ele[20][14] != ele[21][16];
    ele[20][14] != ele[21][17];
    ele[20][14] != ele[22][12];
    ele[20][14] != ele[22][13];
    ele[20][14] != ele[22][14];
    ele[20][14] != ele[22][15];
    ele[20][14] != ele[22][16];
    ele[20][14] != ele[22][17];
    ele[20][14] != ele[23][12];
    ele[20][14] != ele[23][13];
    ele[20][14] != ele[23][14];
    ele[20][14] != ele[23][15];
    ele[20][14] != ele[23][16];
    ele[20][14] != ele[23][17];
    ele[20][14] != ele[24][14];
    ele[20][14] != ele[25][14];
    ele[20][14] != ele[26][14];
    ele[20][14] != ele[27][14];
    ele[20][14] != ele[28][14];
    ele[20][14] != ele[29][14];
    ele[20][14] != ele[30][14];
    ele[20][14] != ele[31][14];
    ele[20][14] != ele[32][14];
    ele[20][14] != ele[33][14];
    ele[20][14] != ele[34][14];
    ele[20][14] != ele[35][14];
    ele[20][15] != ele[20][16];
    ele[20][15] != ele[20][17];
    ele[20][15] != ele[20][18];
    ele[20][15] != ele[20][19];
    ele[20][15] != ele[20][20];
    ele[20][15] != ele[20][21];
    ele[20][15] != ele[20][22];
    ele[20][15] != ele[20][23];
    ele[20][15] != ele[20][24];
    ele[20][15] != ele[20][25];
    ele[20][15] != ele[20][26];
    ele[20][15] != ele[20][27];
    ele[20][15] != ele[20][28];
    ele[20][15] != ele[20][29];
    ele[20][15] != ele[20][30];
    ele[20][15] != ele[20][31];
    ele[20][15] != ele[20][32];
    ele[20][15] != ele[20][33];
    ele[20][15] != ele[20][34];
    ele[20][15] != ele[20][35];
    ele[20][15] != ele[21][12];
    ele[20][15] != ele[21][13];
    ele[20][15] != ele[21][14];
    ele[20][15] != ele[21][15];
    ele[20][15] != ele[21][16];
    ele[20][15] != ele[21][17];
    ele[20][15] != ele[22][12];
    ele[20][15] != ele[22][13];
    ele[20][15] != ele[22][14];
    ele[20][15] != ele[22][15];
    ele[20][15] != ele[22][16];
    ele[20][15] != ele[22][17];
    ele[20][15] != ele[23][12];
    ele[20][15] != ele[23][13];
    ele[20][15] != ele[23][14];
    ele[20][15] != ele[23][15];
    ele[20][15] != ele[23][16];
    ele[20][15] != ele[23][17];
    ele[20][15] != ele[24][15];
    ele[20][15] != ele[25][15];
    ele[20][15] != ele[26][15];
    ele[20][15] != ele[27][15];
    ele[20][15] != ele[28][15];
    ele[20][15] != ele[29][15];
    ele[20][15] != ele[30][15];
    ele[20][15] != ele[31][15];
    ele[20][15] != ele[32][15];
    ele[20][15] != ele[33][15];
    ele[20][15] != ele[34][15];
    ele[20][15] != ele[35][15];
    ele[20][16] != ele[20][17];
    ele[20][16] != ele[20][18];
    ele[20][16] != ele[20][19];
    ele[20][16] != ele[20][20];
    ele[20][16] != ele[20][21];
    ele[20][16] != ele[20][22];
    ele[20][16] != ele[20][23];
    ele[20][16] != ele[20][24];
    ele[20][16] != ele[20][25];
    ele[20][16] != ele[20][26];
    ele[20][16] != ele[20][27];
    ele[20][16] != ele[20][28];
    ele[20][16] != ele[20][29];
    ele[20][16] != ele[20][30];
    ele[20][16] != ele[20][31];
    ele[20][16] != ele[20][32];
    ele[20][16] != ele[20][33];
    ele[20][16] != ele[20][34];
    ele[20][16] != ele[20][35];
    ele[20][16] != ele[21][12];
    ele[20][16] != ele[21][13];
    ele[20][16] != ele[21][14];
    ele[20][16] != ele[21][15];
    ele[20][16] != ele[21][16];
    ele[20][16] != ele[21][17];
    ele[20][16] != ele[22][12];
    ele[20][16] != ele[22][13];
    ele[20][16] != ele[22][14];
    ele[20][16] != ele[22][15];
    ele[20][16] != ele[22][16];
    ele[20][16] != ele[22][17];
    ele[20][16] != ele[23][12];
    ele[20][16] != ele[23][13];
    ele[20][16] != ele[23][14];
    ele[20][16] != ele[23][15];
    ele[20][16] != ele[23][16];
    ele[20][16] != ele[23][17];
    ele[20][16] != ele[24][16];
    ele[20][16] != ele[25][16];
    ele[20][16] != ele[26][16];
    ele[20][16] != ele[27][16];
    ele[20][16] != ele[28][16];
    ele[20][16] != ele[29][16];
    ele[20][16] != ele[30][16];
    ele[20][16] != ele[31][16];
    ele[20][16] != ele[32][16];
    ele[20][16] != ele[33][16];
    ele[20][16] != ele[34][16];
    ele[20][16] != ele[35][16];
    ele[20][17] != ele[20][18];
    ele[20][17] != ele[20][19];
    ele[20][17] != ele[20][20];
    ele[20][17] != ele[20][21];
    ele[20][17] != ele[20][22];
    ele[20][17] != ele[20][23];
    ele[20][17] != ele[20][24];
    ele[20][17] != ele[20][25];
    ele[20][17] != ele[20][26];
    ele[20][17] != ele[20][27];
    ele[20][17] != ele[20][28];
    ele[20][17] != ele[20][29];
    ele[20][17] != ele[20][30];
    ele[20][17] != ele[20][31];
    ele[20][17] != ele[20][32];
    ele[20][17] != ele[20][33];
    ele[20][17] != ele[20][34];
    ele[20][17] != ele[20][35];
    ele[20][17] != ele[21][12];
    ele[20][17] != ele[21][13];
    ele[20][17] != ele[21][14];
    ele[20][17] != ele[21][15];
    ele[20][17] != ele[21][16];
    ele[20][17] != ele[21][17];
    ele[20][17] != ele[22][12];
    ele[20][17] != ele[22][13];
    ele[20][17] != ele[22][14];
    ele[20][17] != ele[22][15];
    ele[20][17] != ele[22][16];
    ele[20][17] != ele[22][17];
    ele[20][17] != ele[23][12];
    ele[20][17] != ele[23][13];
    ele[20][17] != ele[23][14];
    ele[20][17] != ele[23][15];
    ele[20][17] != ele[23][16];
    ele[20][17] != ele[23][17];
    ele[20][17] != ele[24][17];
    ele[20][17] != ele[25][17];
    ele[20][17] != ele[26][17];
    ele[20][17] != ele[27][17];
    ele[20][17] != ele[28][17];
    ele[20][17] != ele[29][17];
    ele[20][17] != ele[30][17];
    ele[20][17] != ele[31][17];
    ele[20][17] != ele[32][17];
    ele[20][17] != ele[33][17];
    ele[20][17] != ele[34][17];
    ele[20][17] != ele[35][17];
    ele[20][18] != ele[20][19];
    ele[20][18] != ele[20][20];
    ele[20][18] != ele[20][21];
    ele[20][18] != ele[20][22];
    ele[20][18] != ele[20][23];
    ele[20][18] != ele[20][24];
    ele[20][18] != ele[20][25];
    ele[20][18] != ele[20][26];
    ele[20][18] != ele[20][27];
    ele[20][18] != ele[20][28];
    ele[20][18] != ele[20][29];
    ele[20][18] != ele[20][30];
    ele[20][18] != ele[20][31];
    ele[20][18] != ele[20][32];
    ele[20][18] != ele[20][33];
    ele[20][18] != ele[20][34];
    ele[20][18] != ele[20][35];
    ele[20][18] != ele[21][18];
    ele[20][18] != ele[21][19];
    ele[20][18] != ele[21][20];
    ele[20][18] != ele[21][21];
    ele[20][18] != ele[21][22];
    ele[20][18] != ele[21][23];
    ele[20][18] != ele[22][18];
    ele[20][18] != ele[22][19];
    ele[20][18] != ele[22][20];
    ele[20][18] != ele[22][21];
    ele[20][18] != ele[22][22];
    ele[20][18] != ele[22][23];
    ele[20][18] != ele[23][18];
    ele[20][18] != ele[23][19];
    ele[20][18] != ele[23][20];
    ele[20][18] != ele[23][21];
    ele[20][18] != ele[23][22];
    ele[20][18] != ele[23][23];
    ele[20][18] != ele[24][18];
    ele[20][18] != ele[25][18];
    ele[20][18] != ele[26][18];
    ele[20][18] != ele[27][18];
    ele[20][18] != ele[28][18];
    ele[20][18] != ele[29][18];
    ele[20][18] != ele[30][18];
    ele[20][18] != ele[31][18];
    ele[20][18] != ele[32][18];
    ele[20][18] != ele[33][18];
    ele[20][18] != ele[34][18];
    ele[20][18] != ele[35][18];
    ele[20][19] != ele[20][20];
    ele[20][19] != ele[20][21];
    ele[20][19] != ele[20][22];
    ele[20][19] != ele[20][23];
    ele[20][19] != ele[20][24];
    ele[20][19] != ele[20][25];
    ele[20][19] != ele[20][26];
    ele[20][19] != ele[20][27];
    ele[20][19] != ele[20][28];
    ele[20][19] != ele[20][29];
    ele[20][19] != ele[20][30];
    ele[20][19] != ele[20][31];
    ele[20][19] != ele[20][32];
    ele[20][19] != ele[20][33];
    ele[20][19] != ele[20][34];
    ele[20][19] != ele[20][35];
    ele[20][19] != ele[21][18];
    ele[20][19] != ele[21][19];
    ele[20][19] != ele[21][20];
    ele[20][19] != ele[21][21];
    ele[20][19] != ele[21][22];
    ele[20][19] != ele[21][23];
    ele[20][19] != ele[22][18];
    ele[20][19] != ele[22][19];
    ele[20][19] != ele[22][20];
    ele[20][19] != ele[22][21];
    ele[20][19] != ele[22][22];
    ele[20][19] != ele[22][23];
    ele[20][19] != ele[23][18];
    ele[20][19] != ele[23][19];
    ele[20][19] != ele[23][20];
    ele[20][19] != ele[23][21];
    ele[20][19] != ele[23][22];
    ele[20][19] != ele[23][23];
    ele[20][19] != ele[24][19];
    ele[20][19] != ele[25][19];
    ele[20][19] != ele[26][19];
    ele[20][19] != ele[27][19];
    ele[20][19] != ele[28][19];
    ele[20][19] != ele[29][19];
    ele[20][19] != ele[30][19];
    ele[20][19] != ele[31][19];
    ele[20][19] != ele[32][19];
    ele[20][19] != ele[33][19];
    ele[20][19] != ele[34][19];
    ele[20][19] != ele[35][19];
    ele[20][2] != ele[20][10];
    ele[20][2] != ele[20][11];
    ele[20][2] != ele[20][12];
    ele[20][2] != ele[20][13];
    ele[20][2] != ele[20][14];
    ele[20][2] != ele[20][15];
    ele[20][2] != ele[20][16];
    ele[20][2] != ele[20][17];
    ele[20][2] != ele[20][18];
    ele[20][2] != ele[20][19];
    ele[20][2] != ele[20][20];
    ele[20][2] != ele[20][21];
    ele[20][2] != ele[20][22];
    ele[20][2] != ele[20][23];
    ele[20][2] != ele[20][24];
    ele[20][2] != ele[20][25];
    ele[20][2] != ele[20][26];
    ele[20][2] != ele[20][27];
    ele[20][2] != ele[20][28];
    ele[20][2] != ele[20][29];
    ele[20][2] != ele[20][3];
    ele[20][2] != ele[20][30];
    ele[20][2] != ele[20][31];
    ele[20][2] != ele[20][32];
    ele[20][2] != ele[20][33];
    ele[20][2] != ele[20][34];
    ele[20][2] != ele[20][35];
    ele[20][2] != ele[20][4];
    ele[20][2] != ele[20][5];
    ele[20][2] != ele[20][6];
    ele[20][2] != ele[20][7];
    ele[20][2] != ele[20][8];
    ele[20][2] != ele[20][9];
    ele[20][2] != ele[21][0];
    ele[20][2] != ele[21][1];
    ele[20][2] != ele[21][2];
    ele[20][2] != ele[21][3];
    ele[20][2] != ele[21][4];
    ele[20][2] != ele[21][5];
    ele[20][2] != ele[22][0];
    ele[20][2] != ele[22][1];
    ele[20][2] != ele[22][2];
    ele[20][2] != ele[22][3];
    ele[20][2] != ele[22][4];
    ele[20][2] != ele[22][5];
    ele[20][2] != ele[23][0];
    ele[20][2] != ele[23][1];
    ele[20][2] != ele[23][2];
    ele[20][2] != ele[23][3];
    ele[20][2] != ele[23][4];
    ele[20][2] != ele[23][5];
    ele[20][2] != ele[24][2];
    ele[20][2] != ele[25][2];
    ele[20][2] != ele[26][2];
    ele[20][2] != ele[27][2];
    ele[20][2] != ele[28][2];
    ele[20][2] != ele[29][2];
    ele[20][2] != ele[30][2];
    ele[20][2] != ele[31][2];
    ele[20][2] != ele[32][2];
    ele[20][2] != ele[33][2];
    ele[20][2] != ele[34][2];
    ele[20][2] != ele[35][2];
    ele[20][20] != ele[20][21];
    ele[20][20] != ele[20][22];
    ele[20][20] != ele[20][23];
    ele[20][20] != ele[20][24];
    ele[20][20] != ele[20][25];
    ele[20][20] != ele[20][26];
    ele[20][20] != ele[20][27];
    ele[20][20] != ele[20][28];
    ele[20][20] != ele[20][29];
    ele[20][20] != ele[20][30];
    ele[20][20] != ele[20][31];
    ele[20][20] != ele[20][32];
    ele[20][20] != ele[20][33];
    ele[20][20] != ele[20][34];
    ele[20][20] != ele[20][35];
    ele[20][20] != ele[21][18];
    ele[20][20] != ele[21][19];
    ele[20][20] != ele[21][20];
    ele[20][20] != ele[21][21];
    ele[20][20] != ele[21][22];
    ele[20][20] != ele[21][23];
    ele[20][20] != ele[22][18];
    ele[20][20] != ele[22][19];
    ele[20][20] != ele[22][20];
    ele[20][20] != ele[22][21];
    ele[20][20] != ele[22][22];
    ele[20][20] != ele[22][23];
    ele[20][20] != ele[23][18];
    ele[20][20] != ele[23][19];
    ele[20][20] != ele[23][20];
    ele[20][20] != ele[23][21];
    ele[20][20] != ele[23][22];
    ele[20][20] != ele[23][23];
    ele[20][20] != ele[24][20];
    ele[20][20] != ele[25][20];
    ele[20][20] != ele[26][20];
    ele[20][20] != ele[27][20];
    ele[20][20] != ele[28][20];
    ele[20][20] != ele[29][20];
    ele[20][20] != ele[30][20];
    ele[20][20] != ele[31][20];
    ele[20][20] != ele[32][20];
    ele[20][20] != ele[33][20];
    ele[20][20] != ele[34][20];
    ele[20][20] != ele[35][20];
    ele[20][21] != ele[20][22];
    ele[20][21] != ele[20][23];
    ele[20][21] != ele[20][24];
    ele[20][21] != ele[20][25];
    ele[20][21] != ele[20][26];
    ele[20][21] != ele[20][27];
    ele[20][21] != ele[20][28];
    ele[20][21] != ele[20][29];
    ele[20][21] != ele[20][30];
    ele[20][21] != ele[20][31];
    ele[20][21] != ele[20][32];
    ele[20][21] != ele[20][33];
    ele[20][21] != ele[20][34];
    ele[20][21] != ele[20][35];
    ele[20][21] != ele[21][18];
    ele[20][21] != ele[21][19];
    ele[20][21] != ele[21][20];
    ele[20][21] != ele[21][21];
    ele[20][21] != ele[21][22];
    ele[20][21] != ele[21][23];
    ele[20][21] != ele[22][18];
    ele[20][21] != ele[22][19];
    ele[20][21] != ele[22][20];
    ele[20][21] != ele[22][21];
    ele[20][21] != ele[22][22];
    ele[20][21] != ele[22][23];
    ele[20][21] != ele[23][18];
    ele[20][21] != ele[23][19];
    ele[20][21] != ele[23][20];
    ele[20][21] != ele[23][21];
    ele[20][21] != ele[23][22];
    ele[20][21] != ele[23][23];
    ele[20][21] != ele[24][21];
    ele[20][21] != ele[25][21];
    ele[20][21] != ele[26][21];
    ele[20][21] != ele[27][21];
    ele[20][21] != ele[28][21];
    ele[20][21] != ele[29][21];
    ele[20][21] != ele[30][21];
    ele[20][21] != ele[31][21];
    ele[20][21] != ele[32][21];
    ele[20][21] != ele[33][21];
    ele[20][21] != ele[34][21];
    ele[20][21] != ele[35][21];
    ele[20][22] != ele[20][23];
    ele[20][22] != ele[20][24];
    ele[20][22] != ele[20][25];
    ele[20][22] != ele[20][26];
    ele[20][22] != ele[20][27];
    ele[20][22] != ele[20][28];
    ele[20][22] != ele[20][29];
    ele[20][22] != ele[20][30];
    ele[20][22] != ele[20][31];
    ele[20][22] != ele[20][32];
    ele[20][22] != ele[20][33];
    ele[20][22] != ele[20][34];
    ele[20][22] != ele[20][35];
    ele[20][22] != ele[21][18];
    ele[20][22] != ele[21][19];
    ele[20][22] != ele[21][20];
    ele[20][22] != ele[21][21];
    ele[20][22] != ele[21][22];
    ele[20][22] != ele[21][23];
    ele[20][22] != ele[22][18];
    ele[20][22] != ele[22][19];
    ele[20][22] != ele[22][20];
    ele[20][22] != ele[22][21];
    ele[20][22] != ele[22][22];
    ele[20][22] != ele[22][23];
    ele[20][22] != ele[23][18];
    ele[20][22] != ele[23][19];
    ele[20][22] != ele[23][20];
    ele[20][22] != ele[23][21];
    ele[20][22] != ele[23][22];
    ele[20][22] != ele[23][23];
    ele[20][22] != ele[24][22];
    ele[20][22] != ele[25][22];
    ele[20][22] != ele[26][22];
    ele[20][22] != ele[27][22];
    ele[20][22] != ele[28][22];
    ele[20][22] != ele[29][22];
    ele[20][22] != ele[30][22];
    ele[20][22] != ele[31][22];
    ele[20][22] != ele[32][22];
    ele[20][22] != ele[33][22];
    ele[20][22] != ele[34][22];
    ele[20][22] != ele[35][22];
    ele[20][23] != ele[20][24];
    ele[20][23] != ele[20][25];
    ele[20][23] != ele[20][26];
    ele[20][23] != ele[20][27];
    ele[20][23] != ele[20][28];
    ele[20][23] != ele[20][29];
    ele[20][23] != ele[20][30];
    ele[20][23] != ele[20][31];
    ele[20][23] != ele[20][32];
    ele[20][23] != ele[20][33];
    ele[20][23] != ele[20][34];
    ele[20][23] != ele[20][35];
    ele[20][23] != ele[21][18];
    ele[20][23] != ele[21][19];
    ele[20][23] != ele[21][20];
    ele[20][23] != ele[21][21];
    ele[20][23] != ele[21][22];
    ele[20][23] != ele[21][23];
    ele[20][23] != ele[22][18];
    ele[20][23] != ele[22][19];
    ele[20][23] != ele[22][20];
    ele[20][23] != ele[22][21];
    ele[20][23] != ele[22][22];
    ele[20][23] != ele[22][23];
    ele[20][23] != ele[23][18];
    ele[20][23] != ele[23][19];
    ele[20][23] != ele[23][20];
    ele[20][23] != ele[23][21];
    ele[20][23] != ele[23][22];
    ele[20][23] != ele[23][23];
    ele[20][23] != ele[24][23];
    ele[20][23] != ele[25][23];
    ele[20][23] != ele[26][23];
    ele[20][23] != ele[27][23];
    ele[20][23] != ele[28][23];
    ele[20][23] != ele[29][23];
    ele[20][23] != ele[30][23];
    ele[20][23] != ele[31][23];
    ele[20][23] != ele[32][23];
    ele[20][23] != ele[33][23];
    ele[20][23] != ele[34][23];
    ele[20][23] != ele[35][23];
    ele[20][24] != ele[20][25];
    ele[20][24] != ele[20][26];
    ele[20][24] != ele[20][27];
    ele[20][24] != ele[20][28];
    ele[20][24] != ele[20][29];
    ele[20][24] != ele[20][30];
    ele[20][24] != ele[20][31];
    ele[20][24] != ele[20][32];
    ele[20][24] != ele[20][33];
    ele[20][24] != ele[20][34];
    ele[20][24] != ele[20][35];
    ele[20][24] != ele[21][24];
    ele[20][24] != ele[21][25];
    ele[20][24] != ele[21][26];
    ele[20][24] != ele[21][27];
    ele[20][24] != ele[21][28];
    ele[20][24] != ele[21][29];
    ele[20][24] != ele[22][24];
    ele[20][24] != ele[22][25];
    ele[20][24] != ele[22][26];
    ele[20][24] != ele[22][27];
    ele[20][24] != ele[22][28];
    ele[20][24] != ele[22][29];
    ele[20][24] != ele[23][24];
    ele[20][24] != ele[23][25];
    ele[20][24] != ele[23][26];
    ele[20][24] != ele[23][27];
    ele[20][24] != ele[23][28];
    ele[20][24] != ele[23][29];
    ele[20][24] != ele[24][24];
    ele[20][24] != ele[25][24];
    ele[20][24] != ele[26][24];
    ele[20][24] != ele[27][24];
    ele[20][24] != ele[28][24];
    ele[20][24] != ele[29][24];
    ele[20][24] != ele[30][24];
    ele[20][24] != ele[31][24];
    ele[20][24] != ele[32][24];
    ele[20][24] != ele[33][24];
    ele[20][24] != ele[34][24];
    ele[20][24] != ele[35][24];
    ele[20][25] != ele[20][26];
    ele[20][25] != ele[20][27];
    ele[20][25] != ele[20][28];
    ele[20][25] != ele[20][29];
    ele[20][25] != ele[20][30];
    ele[20][25] != ele[20][31];
    ele[20][25] != ele[20][32];
    ele[20][25] != ele[20][33];
    ele[20][25] != ele[20][34];
    ele[20][25] != ele[20][35];
    ele[20][25] != ele[21][24];
    ele[20][25] != ele[21][25];
    ele[20][25] != ele[21][26];
    ele[20][25] != ele[21][27];
    ele[20][25] != ele[21][28];
    ele[20][25] != ele[21][29];
    ele[20][25] != ele[22][24];
    ele[20][25] != ele[22][25];
    ele[20][25] != ele[22][26];
    ele[20][25] != ele[22][27];
    ele[20][25] != ele[22][28];
    ele[20][25] != ele[22][29];
    ele[20][25] != ele[23][24];
    ele[20][25] != ele[23][25];
    ele[20][25] != ele[23][26];
    ele[20][25] != ele[23][27];
    ele[20][25] != ele[23][28];
    ele[20][25] != ele[23][29];
    ele[20][25] != ele[24][25];
    ele[20][25] != ele[25][25];
    ele[20][25] != ele[26][25];
    ele[20][25] != ele[27][25];
    ele[20][25] != ele[28][25];
    ele[20][25] != ele[29][25];
    ele[20][25] != ele[30][25];
    ele[20][25] != ele[31][25];
    ele[20][25] != ele[32][25];
    ele[20][25] != ele[33][25];
    ele[20][25] != ele[34][25];
    ele[20][25] != ele[35][25];
    ele[20][26] != ele[20][27];
    ele[20][26] != ele[20][28];
    ele[20][26] != ele[20][29];
    ele[20][26] != ele[20][30];
    ele[20][26] != ele[20][31];
    ele[20][26] != ele[20][32];
    ele[20][26] != ele[20][33];
    ele[20][26] != ele[20][34];
    ele[20][26] != ele[20][35];
    ele[20][26] != ele[21][24];
    ele[20][26] != ele[21][25];
    ele[20][26] != ele[21][26];
    ele[20][26] != ele[21][27];
    ele[20][26] != ele[21][28];
    ele[20][26] != ele[21][29];
    ele[20][26] != ele[22][24];
    ele[20][26] != ele[22][25];
    ele[20][26] != ele[22][26];
    ele[20][26] != ele[22][27];
    ele[20][26] != ele[22][28];
    ele[20][26] != ele[22][29];
    ele[20][26] != ele[23][24];
    ele[20][26] != ele[23][25];
    ele[20][26] != ele[23][26];
    ele[20][26] != ele[23][27];
    ele[20][26] != ele[23][28];
    ele[20][26] != ele[23][29];
    ele[20][26] != ele[24][26];
    ele[20][26] != ele[25][26];
    ele[20][26] != ele[26][26];
    ele[20][26] != ele[27][26];
    ele[20][26] != ele[28][26];
    ele[20][26] != ele[29][26];
    ele[20][26] != ele[30][26];
    ele[20][26] != ele[31][26];
    ele[20][26] != ele[32][26];
    ele[20][26] != ele[33][26];
    ele[20][26] != ele[34][26];
    ele[20][26] != ele[35][26];
    ele[20][27] != ele[20][28];
    ele[20][27] != ele[20][29];
    ele[20][27] != ele[20][30];
    ele[20][27] != ele[20][31];
    ele[20][27] != ele[20][32];
    ele[20][27] != ele[20][33];
    ele[20][27] != ele[20][34];
    ele[20][27] != ele[20][35];
    ele[20][27] != ele[21][24];
    ele[20][27] != ele[21][25];
    ele[20][27] != ele[21][26];
    ele[20][27] != ele[21][27];
    ele[20][27] != ele[21][28];
    ele[20][27] != ele[21][29];
    ele[20][27] != ele[22][24];
    ele[20][27] != ele[22][25];
    ele[20][27] != ele[22][26];
    ele[20][27] != ele[22][27];
    ele[20][27] != ele[22][28];
    ele[20][27] != ele[22][29];
    ele[20][27] != ele[23][24];
    ele[20][27] != ele[23][25];
    ele[20][27] != ele[23][26];
    ele[20][27] != ele[23][27];
    ele[20][27] != ele[23][28];
    ele[20][27] != ele[23][29];
    ele[20][27] != ele[24][27];
    ele[20][27] != ele[25][27];
    ele[20][27] != ele[26][27];
    ele[20][27] != ele[27][27];
    ele[20][27] != ele[28][27];
    ele[20][27] != ele[29][27];
    ele[20][27] != ele[30][27];
    ele[20][27] != ele[31][27];
    ele[20][27] != ele[32][27];
    ele[20][27] != ele[33][27];
    ele[20][27] != ele[34][27];
    ele[20][27] != ele[35][27];
    ele[20][28] != ele[20][29];
    ele[20][28] != ele[20][30];
    ele[20][28] != ele[20][31];
    ele[20][28] != ele[20][32];
    ele[20][28] != ele[20][33];
    ele[20][28] != ele[20][34];
    ele[20][28] != ele[20][35];
    ele[20][28] != ele[21][24];
    ele[20][28] != ele[21][25];
    ele[20][28] != ele[21][26];
    ele[20][28] != ele[21][27];
    ele[20][28] != ele[21][28];
    ele[20][28] != ele[21][29];
    ele[20][28] != ele[22][24];
    ele[20][28] != ele[22][25];
    ele[20][28] != ele[22][26];
    ele[20][28] != ele[22][27];
    ele[20][28] != ele[22][28];
    ele[20][28] != ele[22][29];
    ele[20][28] != ele[23][24];
    ele[20][28] != ele[23][25];
    ele[20][28] != ele[23][26];
    ele[20][28] != ele[23][27];
    ele[20][28] != ele[23][28];
    ele[20][28] != ele[23][29];
    ele[20][28] != ele[24][28];
    ele[20][28] != ele[25][28];
    ele[20][28] != ele[26][28];
    ele[20][28] != ele[27][28];
    ele[20][28] != ele[28][28];
    ele[20][28] != ele[29][28];
    ele[20][28] != ele[30][28];
    ele[20][28] != ele[31][28];
    ele[20][28] != ele[32][28];
    ele[20][28] != ele[33][28];
    ele[20][28] != ele[34][28];
    ele[20][28] != ele[35][28];
    ele[20][29] != ele[20][30];
    ele[20][29] != ele[20][31];
    ele[20][29] != ele[20][32];
    ele[20][29] != ele[20][33];
    ele[20][29] != ele[20][34];
    ele[20][29] != ele[20][35];
    ele[20][29] != ele[21][24];
    ele[20][29] != ele[21][25];
    ele[20][29] != ele[21][26];
    ele[20][29] != ele[21][27];
    ele[20][29] != ele[21][28];
    ele[20][29] != ele[21][29];
    ele[20][29] != ele[22][24];
    ele[20][29] != ele[22][25];
    ele[20][29] != ele[22][26];
    ele[20][29] != ele[22][27];
    ele[20][29] != ele[22][28];
    ele[20][29] != ele[22][29];
    ele[20][29] != ele[23][24];
    ele[20][29] != ele[23][25];
    ele[20][29] != ele[23][26];
    ele[20][29] != ele[23][27];
    ele[20][29] != ele[23][28];
    ele[20][29] != ele[23][29];
    ele[20][29] != ele[24][29];
    ele[20][29] != ele[25][29];
    ele[20][29] != ele[26][29];
    ele[20][29] != ele[27][29];
    ele[20][29] != ele[28][29];
    ele[20][29] != ele[29][29];
    ele[20][29] != ele[30][29];
    ele[20][29] != ele[31][29];
    ele[20][29] != ele[32][29];
    ele[20][29] != ele[33][29];
    ele[20][29] != ele[34][29];
    ele[20][29] != ele[35][29];
    ele[20][3] != ele[20][10];
    ele[20][3] != ele[20][11];
    ele[20][3] != ele[20][12];
    ele[20][3] != ele[20][13];
    ele[20][3] != ele[20][14];
    ele[20][3] != ele[20][15];
    ele[20][3] != ele[20][16];
    ele[20][3] != ele[20][17];
    ele[20][3] != ele[20][18];
    ele[20][3] != ele[20][19];
    ele[20][3] != ele[20][20];
    ele[20][3] != ele[20][21];
    ele[20][3] != ele[20][22];
    ele[20][3] != ele[20][23];
    ele[20][3] != ele[20][24];
    ele[20][3] != ele[20][25];
    ele[20][3] != ele[20][26];
    ele[20][3] != ele[20][27];
    ele[20][3] != ele[20][28];
    ele[20][3] != ele[20][29];
    ele[20][3] != ele[20][30];
    ele[20][3] != ele[20][31];
    ele[20][3] != ele[20][32];
    ele[20][3] != ele[20][33];
    ele[20][3] != ele[20][34];
    ele[20][3] != ele[20][35];
    ele[20][3] != ele[20][4];
    ele[20][3] != ele[20][5];
    ele[20][3] != ele[20][6];
    ele[20][3] != ele[20][7];
    ele[20][3] != ele[20][8];
    ele[20][3] != ele[20][9];
    ele[20][3] != ele[21][0];
    ele[20][3] != ele[21][1];
    ele[20][3] != ele[21][2];
    ele[20][3] != ele[21][3];
    ele[20][3] != ele[21][4];
    ele[20][3] != ele[21][5];
    ele[20][3] != ele[22][0];
    ele[20][3] != ele[22][1];
    ele[20][3] != ele[22][2];
    ele[20][3] != ele[22][3];
    ele[20][3] != ele[22][4];
    ele[20][3] != ele[22][5];
    ele[20][3] != ele[23][0];
    ele[20][3] != ele[23][1];
    ele[20][3] != ele[23][2];
    ele[20][3] != ele[23][3];
    ele[20][3] != ele[23][4];
    ele[20][3] != ele[23][5];
    ele[20][3] != ele[24][3];
    ele[20][3] != ele[25][3];
    ele[20][3] != ele[26][3];
    ele[20][3] != ele[27][3];
    ele[20][3] != ele[28][3];
    ele[20][3] != ele[29][3];
    ele[20][3] != ele[30][3];
    ele[20][3] != ele[31][3];
    ele[20][3] != ele[32][3];
    ele[20][3] != ele[33][3];
    ele[20][3] != ele[34][3];
    ele[20][3] != ele[35][3];
    ele[20][30] != ele[20][31];
    ele[20][30] != ele[20][32];
    ele[20][30] != ele[20][33];
    ele[20][30] != ele[20][34];
    ele[20][30] != ele[20][35];
    ele[20][30] != ele[21][30];
    ele[20][30] != ele[21][31];
    ele[20][30] != ele[21][32];
    ele[20][30] != ele[21][33];
    ele[20][30] != ele[21][34];
    ele[20][30] != ele[21][35];
    ele[20][30] != ele[22][30];
    ele[20][30] != ele[22][31];
    ele[20][30] != ele[22][32];
    ele[20][30] != ele[22][33];
    ele[20][30] != ele[22][34];
    ele[20][30] != ele[22][35];
    ele[20][30] != ele[23][30];
    ele[20][30] != ele[23][31];
    ele[20][30] != ele[23][32];
    ele[20][30] != ele[23][33];
    ele[20][30] != ele[23][34];
    ele[20][30] != ele[23][35];
    ele[20][30] != ele[24][30];
    ele[20][30] != ele[25][30];
    ele[20][30] != ele[26][30];
    ele[20][30] != ele[27][30];
    ele[20][30] != ele[28][30];
    ele[20][30] != ele[29][30];
    ele[20][30] != ele[30][30];
    ele[20][30] != ele[31][30];
    ele[20][30] != ele[32][30];
    ele[20][30] != ele[33][30];
    ele[20][30] != ele[34][30];
    ele[20][30] != ele[35][30];
    ele[20][31] != ele[20][32];
    ele[20][31] != ele[20][33];
    ele[20][31] != ele[20][34];
    ele[20][31] != ele[20][35];
    ele[20][31] != ele[21][30];
    ele[20][31] != ele[21][31];
    ele[20][31] != ele[21][32];
    ele[20][31] != ele[21][33];
    ele[20][31] != ele[21][34];
    ele[20][31] != ele[21][35];
    ele[20][31] != ele[22][30];
    ele[20][31] != ele[22][31];
    ele[20][31] != ele[22][32];
    ele[20][31] != ele[22][33];
    ele[20][31] != ele[22][34];
    ele[20][31] != ele[22][35];
    ele[20][31] != ele[23][30];
    ele[20][31] != ele[23][31];
    ele[20][31] != ele[23][32];
    ele[20][31] != ele[23][33];
    ele[20][31] != ele[23][34];
    ele[20][31] != ele[23][35];
    ele[20][31] != ele[24][31];
    ele[20][31] != ele[25][31];
    ele[20][31] != ele[26][31];
    ele[20][31] != ele[27][31];
    ele[20][31] != ele[28][31];
    ele[20][31] != ele[29][31];
    ele[20][31] != ele[30][31];
    ele[20][31] != ele[31][31];
    ele[20][31] != ele[32][31];
    ele[20][31] != ele[33][31];
    ele[20][31] != ele[34][31];
    ele[20][31] != ele[35][31];
    ele[20][32] != ele[20][33];
    ele[20][32] != ele[20][34];
    ele[20][32] != ele[20][35];
    ele[20][32] != ele[21][30];
    ele[20][32] != ele[21][31];
    ele[20][32] != ele[21][32];
    ele[20][32] != ele[21][33];
    ele[20][32] != ele[21][34];
    ele[20][32] != ele[21][35];
    ele[20][32] != ele[22][30];
    ele[20][32] != ele[22][31];
    ele[20][32] != ele[22][32];
    ele[20][32] != ele[22][33];
    ele[20][32] != ele[22][34];
    ele[20][32] != ele[22][35];
    ele[20][32] != ele[23][30];
    ele[20][32] != ele[23][31];
    ele[20][32] != ele[23][32];
    ele[20][32] != ele[23][33];
    ele[20][32] != ele[23][34];
    ele[20][32] != ele[23][35];
    ele[20][32] != ele[24][32];
    ele[20][32] != ele[25][32];
    ele[20][32] != ele[26][32];
    ele[20][32] != ele[27][32];
    ele[20][32] != ele[28][32];
    ele[20][32] != ele[29][32];
    ele[20][32] != ele[30][32];
    ele[20][32] != ele[31][32];
    ele[20][32] != ele[32][32];
    ele[20][32] != ele[33][32];
    ele[20][32] != ele[34][32];
    ele[20][32] != ele[35][32];
    ele[20][33] != ele[20][34];
    ele[20][33] != ele[20][35];
    ele[20][33] != ele[21][30];
    ele[20][33] != ele[21][31];
    ele[20][33] != ele[21][32];
    ele[20][33] != ele[21][33];
    ele[20][33] != ele[21][34];
    ele[20][33] != ele[21][35];
    ele[20][33] != ele[22][30];
    ele[20][33] != ele[22][31];
    ele[20][33] != ele[22][32];
    ele[20][33] != ele[22][33];
    ele[20][33] != ele[22][34];
    ele[20][33] != ele[22][35];
    ele[20][33] != ele[23][30];
    ele[20][33] != ele[23][31];
    ele[20][33] != ele[23][32];
    ele[20][33] != ele[23][33];
    ele[20][33] != ele[23][34];
    ele[20][33] != ele[23][35];
    ele[20][33] != ele[24][33];
    ele[20][33] != ele[25][33];
    ele[20][33] != ele[26][33];
    ele[20][33] != ele[27][33];
    ele[20][33] != ele[28][33];
    ele[20][33] != ele[29][33];
    ele[20][33] != ele[30][33];
    ele[20][33] != ele[31][33];
    ele[20][33] != ele[32][33];
    ele[20][33] != ele[33][33];
    ele[20][33] != ele[34][33];
    ele[20][33] != ele[35][33];
    ele[20][34] != ele[20][35];
    ele[20][34] != ele[21][30];
    ele[20][34] != ele[21][31];
    ele[20][34] != ele[21][32];
    ele[20][34] != ele[21][33];
    ele[20][34] != ele[21][34];
    ele[20][34] != ele[21][35];
    ele[20][34] != ele[22][30];
    ele[20][34] != ele[22][31];
    ele[20][34] != ele[22][32];
    ele[20][34] != ele[22][33];
    ele[20][34] != ele[22][34];
    ele[20][34] != ele[22][35];
    ele[20][34] != ele[23][30];
    ele[20][34] != ele[23][31];
    ele[20][34] != ele[23][32];
    ele[20][34] != ele[23][33];
    ele[20][34] != ele[23][34];
    ele[20][34] != ele[23][35];
    ele[20][34] != ele[24][34];
    ele[20][34] != ele[25][34];
    ele[20][34] != ele[26][34];
    ele[20][34] != ele[27][34];
    ele[20][34] != ele[28][34];
    ele[20][34] != ele[29][34];
    ele[20][34] != ele[30][34];
    ele[20][34] != ele[31][34];
    ele[20][34] != ele[32][34];
    ele[20][34] != ele[33][34];
    ele[20][34] != ele[34][34];
    ele[20][34] != ele[35][34];
    ele[20][35] != ele[21][30];
    ele[20][35] != ele[21][31];
    ele[20][35] != ele[21][32];
    ele[20][35] != ele[21][33];
    ele[20][35] != ele[21][34];
    ele[20][35] != ele[21][35];
    ele[20][35] != ele[22][30];
    ele[20][35] != ele[22][31];
    ele[20][35] != ele[22][32];
    ele[20][35] != ele[22][33];
    ele[20][35] != ele[22][34];
    ele[20][35] != ele[22][35];
    ele[20][35] != ele[23][30];
    ele[20][35] != ele[23][31];
    ele[20][35] != ele[23][32];
    ele[20][35] != ele[23][33];
    ele[20][35] != ele[23][34];
    ele[20][35] != ele[23][35];
    ele[20][35] != ele[24][35];
    ele[20][35] != ele[25][35];
    ele[20][35] != ele[26][35];
    ele[20][35] != ele[27][35];
    ele[20][35] != ele[28][35];
    ele[20][35] != ele[29][35];
    ele[20][35] != ele[30][35];
    ele[20][35] != ele[31][35];
    ele[20][35] != ele[32][35];
    ele[20][35] != ele[33][35];
    ele[20][35] != ele[34][35];
    ele[20][35] != ele[35][35];
    ele[20][4] != ele[20][10];
    ele[20][4] != ele[20][11];
    ele[20][4] != ele[20][12];
    ele[20][4] != ele[20][13];
    ele[20][4] != ele[20][14];
    ele[20][4] != ele[20][15];
    ele[20][4] != ele[20][16];
    ele[20][4] != ele[20][17];
    ele[20][4] != ele[20][18];
    ele[20][4] != ele[20][19];
    ele[20][4] != ele[20][20];
    ele[20][4] != ele[20][21];
    ele[20][4] != ele[20][22];
    ele[20][4] != ele[20][23];
    ele[20][4] != ele[20][24];
    ele[20][4] != ele[20][25];
    ele[20][4] != ele[20][26];
    ele[20][4] != ele[20][27];
    ele[20][4] != ele[20][28];
    ele[20][4] != ele[20][29];
    ele[20][4] != ele[20][30];
    ele[20][4] != ele[20][31];
    ele[20][4] != ele[20][32];
    ele[20][4] != ele[20][33];
    ele[20][4] != ele[20][34];
    ele[20][4] != ele[20][35];
    ele[20][4] != ele[20][5];
    ele[20][4] != ele[20][6];
    ele[20][4] != ele[20][7];
    ele[20][4] != ele[20][8];
    ele[20][4] != ele[20][9];
    ele[20][4] != ele[21][0];
    ele[20][4] != ele[21][1];
    ele[20][4] != ele[21][2];
    ele[20][4] != ele[21][3];
    ele[20][4] != ele[21][4];
    ele[20][4] != ele[21][5];
    ele[20][4] != ele[22][0];
    ele[20][4] != ele[22][1];
    ele[20][4] != ele[22][2];
    ele[20][4] != ele[22][3];
    ele[20][4] != ele[22][4];
    ele[20][4] != ele[22][5];
    ele[20][4] != ele[23][0];
    ele[20][4] != ele[23][1];
    ele[20][4] != ele[23][2];
    ele[20][4] != ele[23][3];
    ele[20][4] != ele[23][4];
    ele[20][4] != ele[23][5];
    ele[20][4] != ele[24][4];
    ele[20][4] != ele[25][4];
    ele[20][4] != ele[26][4];
    ele[20][4] != ele[27][4];
    ele[20][4] != ele[28][4];
    ele[20][4] != ele[29][4];
    ele[20][4] != ele[30][4];
    ele[20][4] != ele[31][4];
    ele[20][4] != ele[32][4];
    ele[20][4] != ele[33][4];
    ele[20][4] != ele[34][4];
    ele[20][4] != ele[35][4];
    ele[20][5] != ele[20][10];
    ele[20][5] != ele[20][11];
    ele[20][5] != ele[20][12];
    ele[20][5] != ele[20][13];
    ele[20][5] != ele[20][14];
    ele[20][5] != ele[20][15];
    ele[20][5] != ele[20][16];
    ele[20][5] != ele[20][17];
    ele[20][5] != ele[20][18];
    ele[20][5] != ele[20][19];
    ele[20][5] != ele[20][20];
    ele[20][5] != ele[20][21];
    ele[20][5] != ele[20][22];
    ele[20][5] != ele[20][23];
    ele[20][5] != ele[20][24];
    ele[20][5] != ele[20][25];
    ele[20][5] != ele[20][26];
    ele[20][5] != ele[20][27];
    ele[20][5] != ele[20][28];
    ele[20][5] != ele[20][29];
    ele[20][5] != ele[20][30];
    ele[20][5] != ele[20][31];
    ele[20][5] != ele[20][32];
    ele[20][5] != ele[20][33];
    ele[20][5] != ele[20][34];
    ele[20][5] != ele[20][35];
    ele[20][5] != ele[20][6];
    ele[20][5] != ele[20][7];
    ele[20][5] != ele[20][8];
    ele[20][5] != ele[20][9];
    ele[20][5] != ele[21][0];
    ele[20][5] != ele[21][1];
    ele[20][5] != ele[21][2];
    ele[20][5] != ele[21][3];
    ele[20][5] != ele[21][4];
    ele[20][5] != ele[21][5];
    ele[20][5] != ele[22][0];
    ele[20][5] != ele[22][1];
    ele[20][5] != ele[22][2];
    ele[20][5] != ele[22][3];
    ele[20][5] != ele[22][4];
    ele[20][5] != ele[22][5];
    ele[20][5] != ele[23][0];
    ele[20][5] != ele[23][1];
    ele[20][5] != ele[23][2];
    ele[20][5] != ele[23][3];
    ele[20][5] != ele[23][4];
    ele[20][5] != ele[23][5];
    ele[20][5] != ele[24][5];
    ele[20][5] != ele[25][5];
    ele[20][5] != ele[26][5];
    ele[20][5] != ele[27][5];
    ele[20][5] != ele[28][5];
    ele[20][5] != ele[29][5];
    ele[20][5] != ele[30][5];
    ele[20][5] != ele[31][5];
    ele[20][5] != ele[32][5];
    ele[20][5] != ele[33][5];
    ele[20][5] != ele[34][5];
    ele[20][5] != ele[35][5];
    ele[20][6] != ele[20][10];
    ele[20][6] != ele[20][11];
    ele[20][6] != ele[20][12];
    ele[20][6] != ele[20][13];
    ele[20][6] != ele[20][14];
    ele[20][6] != ele[20][15];
    ele[20][6] != ele[20][16];
    ele[20][6] != ele[20][17];
    ele[20][6] != ele[20][18];
    ele[20][6] != ele[20][19];
    ele[20][6] != ele[20][20];
    ele[20][6] != ele[20][21];
    ele[20][6] != ele[20][22];
    ele[20][6] != ele[20][23];
    ele[20][6] != ele[20][24];
    ele[20][6] != ele[20][25];
    ele[20][6] != ele[20][26];
    ele[20][6] != ele[20][27];
    ele[20][6] != ele[20][28];
    ele[20][6] != ele[20][29];
    ele[20][6] != ele[20][30];
    ele[20][6] != ele[20][31];
    ele[20][6] != ele[20][32];
    ele[20][6] != ele[20][33];
    ele[20][6] != ele[20][34];
    ele[20][6] != ele[20][35];
    ele[20][6] != ele[20][7];
    ele[20][6] != ele[20][8];
    ele[20][6] != ele[20][9];
    ele[20][6] != ele[21][10];
    ele[20][6] != ele[21][11];
    ele[20][6] != ele[21][6];
    ele[20][6] != ele[21][7];
    ele[20][6] != ele[21][8];
    ele[20][6] != ele[21][9];
    ele[20][6] != ele[22][10];
    ele[20][6] != ele[22][11];
    ele[20][6] != ele[22][6];
    ele[20][6] != ele[22][7];
    ele[20][6] != ele[22][8];
    ele[20][6] != ele[22][9];
    ele[20][6] != ele[23][10];
    ele[20][6] != ele[23][11];
    ele[20][6] != ele[23][6];
    ele[20][6] != ele[23][7];
    ele[20][6] != ele[23][8];
    ele[20][6] != ele[23][9];
    ele[20][6] != ele[24][6];
    ele[20][6] != ele[25][6];
    ele[20][6] != ele[26][6];
    ele[20][6] != ele[27][6];
    ele[20][6] != ele[28][6];
    ele[20][6] != ele[29][6];
    ele[20][6] != ele[30][6];
    ele[20][6] != ele[31][6];
    ele[20][6] != ele[32][6];
    ele[20][6] != ele[33][6];
    ele[20][6] != ele[34][6];
    ele[20][6] != ele[35][6];
    ele[20][7] != ele[20][10];
    ele[20][7] != ele[20][11];
    ele[20][7] != ele[20][12];
    ele[20][7] != ele[20][13];
    ele[20][7] != ele[20][14];
    ele[20][7] != ele[20][15];
    ele[20][7] != ele[20][16];
    ele[20][7] != ele[20][17];
    ele[20][7] != ele[20][18];
    ele[20][7] != ele[20][19];
    ele[20][7] != ele[20][20];
    ele[20][7] != ele[20][21];
    ele[20][7] != ele[20][22];
    ele[20][7] != ele[20][23];
    ele[20][7] != ele[20][24];
    ele[20][7] != ele[20][25];
    ele[20][7] != ele[20][26];
    ele[20][7] != ele[20][27];
    ele[20][7] != ele[20][28];
    ele[20][7] != ele[20][29];
    ele[20][7] != ele[20][30];
    ele[20][7] != ele[20][31];
    ele[20][7] != ele[20][32];
    ele[20][7] != ele[20][33];
    ele[20][7] != ele[20][34];
    ele[20][7] != ele[20][35];
    ele[20][7] != ele[20][8];
    ele[20][7] != ele[20][9];
    ele[20][7] != ele[21][10];
    ele[20][7] != ele[21][11];
    ele[20][7] != ele[21][6];
    ele[20][7] != ele[21][7];
    ele[20][7] != ele[21][8];
    ele[20][7] != ele[21][9];
    ele[20][7] != ele[22][10];
    ele[20][7] != ele[22][11];
    ele[20][7] != ele[22][6];
    ele[20][7] != ele[22][7];
    ele[20][7] != ele[22][8];
    ele[20][7] != ele[22][9];
    ele[20][7] != ele[23][10];
    ele[20][7] != ele[23][11];
    ele[20][7] != ele[23][6];
    ele[20][7] != ele[23][7];
    ele[20][7] != ele[23][8];
    ele[20][7] != ele[23][9];
    ele[20][7] != ele[24][7];
    ele[20][7] != ele[25][7];
    ele[20][7] != ele[26][7];
    ele[20][7] != ele[27][7];
    ele[20][7] != ele[28][7];
    ele[20][7] != ele[29][7];
    ele[20][7] != ele[30][7];
    ele[20][7] != ele[31][7];
    ele[20][7] != ele[32][7];
    ele[20][7] != ele[33][7];
    ele[20][7] != ele[34][7];
    ele[20][7] != ele[35][7];
    ele[20][8] != ele[20][10];
    ele[20][8] != ele[20][11];
    ele[20][8] != ele[20][12];
    ele[20][8] != ele[20][13];
    ele[20][8] != ele[20][14];
    ele[20][8] != ele[20][15];
    ele[20][8] != ele[20][16];
    ele[20][8] != ele[20][17];
    ele[20][8] != ele[20][18];
    ele[20][8] != ele[20][19];
    ele[20][8] != ele[20][20];
    ele[20][8] != ele[20][21];
    ele[20][8] != ele[20][22];
    ele[20][8] != ele[20][23];
    ele[20][8] != ele[20][24];
    ele[20][8] != ele[20][25];
    ele[20][8] != ele[20][26];
    ele[20][8] != ele[20][27];
    ele[20][8] != ele[20][28];
    ele[20][8] != ele[20][29];
    ele[20][8] != ele[20][30];
    ele[20][8] != ele[20][31];
    ele[20][8] != ele[20][32];
    ele[20][8] != ele[20][33];
    ele[20][8] != ele[20][34];
    ele[20][8] != ele[20][35];
    ele[20][8] != ele[20][9];
    ele[20][8] != ele[21][10];
    ele[20][8] != ele[21][11];
    ele[20][8] != ele[21][6];
    ele[20][8] != ele[21][7];
    ele[20][8] != ele[21][8];
    ele[20][8] != ele[21][9];
    ele[20][8] != ele[22][10];
    ele[20][8] != ele[22][11];
    ele[20][8] != ele[22][6];
    ele[20][8] != ele[22][7];
    ele[20][8] != ele[22][8];
    ele[20][8] != ele[22][9];
    ele[20][8] != ele[23][10];
    ele[20][8] != ele[23][11];
    ele[20][8] != ele[23][6];
    ele[20][8] != ele[23][7];
    ele[20][8] != ele[23][8];
    ele[20][8] != ele[23][9];
    ele[20][8] != ele[24][8];
    ele[20][8] != ele[25][8];
    ele[20][8] != ele[26][8];
    ele[20][8] != ele[27][8];
    ele[20][8] != ele[28][8];
    ele[20][8] != ele[29][8];
    ele[20][8] != ele[30][8];
    ele[20][8] != ele[31][8];
    ele[20][8] != ele[32][8];
    ele[20][8] != ele[33][8];
    ele[20][8] != ele[34][8];
    ele[20][8] != ele[35][8];
    ele[20][9] != ele[20][10];
    ele[20][9] != ele[20][11];
    ele[20][9] != ele[20][12];
    ele[20][9] != ele[20][13];
    ele[20][9] != ele[20][14];
    ele[20][9] != ele[20][15];
    ele[20][9] != ele[20][16];
    ele[20][9] != ele[20][17];
    ele[20][9] != ele[20][18];
    ele[20][9] != ele[20][19];
    ele[20][9] != ele[20][20];
    ele[20][9] != ele[20][21];
    ele[20][9] != ele[20][22];
    ele[20][9] != ele[20][23];
    ele[20][9] != ele[20][24];
    ele[20][9] != ele[20][25];
    ele[20][9] != ele[20][26];
    ele[20][9] != ele[20][27];
    ele[20][9] != ele[20][28];
    ele[20][9] != ele[20][29];
    ele[20][9] != ele[20][30];
    ele[20][9] != ele[20][31];
    ele[20][9] != ele[20][32];
    ele[20][9] != ele[20][33];
    ele[20][9] != ele[20][34];
    ele[20][9] != ele[20][35];
    ele[20][9] != ele[21][10];
    ele[20][9] != ele[21][11];
    ele[20][9] != ele[21][6];
    ele[20][9] != ele[21][7];
    ele[20][9] != ele[21][8];
    ele[20][9] != ele[21][9];
    ele[20][9] != ele[22][10];
    ele[20][9] != ele[22][11];
    ele[20][9] != ele[22][6];
    ele[20][9] != ele[22][7];
    ele[20][9] != ele[22][8];
    ele[20][9] != ele[22][9];
    ele[20][9] != ele[23][10];
    ele[20][9] != ele[23][11];
    ele[20][9] != ele[23][6];
    ele[20][9] != ele[23][7];
    ele[20][9] != ele[23][8];
    ele[20][9] != ele[23][9];
    ele[20][9] != ele[24][9];
    ele[20][9] != ele[25][9];
    ele[20][9] != ele[26][9];
    ele[20][9] != ele[27][9];
    ele[20][9] != ele[28][9];
    ele[20][9] != ele[29][9];
    ele[20][9] != ele[30][9];
    ele[20][9] != ele[31][9];
    ele[20][9] != ele[32][9];
    ele[20][9] != ele[33][9];
    ele[20][9] != ele[34][9];
    ele[20][9] != ele[35][9];
    ele[21][0] != ele[21][1];
    ele[21][0] != ele[21][10];
    ele[21][0] != ele[21][11];
    ele[21][0] != ele[21][12];
    ele[21][0] != ele[21][13];
    ele[21][0] != ele[21][14];
    ele[21][0] != ele[21][15];
    ele[21][0] != ele[21][16];
    ele[21][0] != ele[21][17];
    ele[21][0] != ele[21][18];
    ele[21][0] != ele[21][19];
    ele[21][0] != ele[21][2];
    ele[21][0] != ele[21][20];
    ele[21][0] != ele[21][21];
    ele[21][0] != ele[21][22];
    ele[21][0] != ele[21][23];
    ele[21][0] != ele[21][24];
    ele[21][0] != ele[21][25];
    ele[21][0] != ele[21][26];
    ele[21][0] != ele[21][27];
    ele[21][0] != ele[21][28];
    ele[21][0] != ele[21][29];
    ele[21][0] != ele[21][3];
    ele[21][0] != ele[21][30];
    ele[21][0] != ele[21][31];
    ele[21][0] != ele[21][32];
    ele[21][0] != ele[21][33];
    ele[21][0] != ele[21][34];
    ele[21][0] != ele[21][35];
    ele[21][0] != ele[21][4];
    ele[21][0] != ele[21][5];
    ele[21][0] != ele[21][6];
    ele[21][0] != ele[21][7];
    ele[21][0] != ele[21][8];
    ele[21][0] != ele[21][9];
    ele[21][0] != ele[22][0];
    ele[21][0] != ele[22][1];
    ele[21][0] != ele[22][2];
    ele[21][0] != ele[22][3];
    ele[21][0] != ele[22][4];
    ele[21][0] != ele[22][5];
    ele[21][0] != ele[23][0];
    ele[21][0] != ele[23][1];
    ele[21][0] != ele[23][2];
    ele[21][0] != ele[23][3];
    ele[21][0] != ele[23][4];
    ele[21][0] != ele[23][5];
    ele[21][0] != ele[24][0];
    ele[21][0] != ele[25][0];
    ele[21][0] != ele[26][0];
    ele[21][0] != ele[27][0];
    ele[21][0] != ele[28][0];
    ele[21][0] != ele[29][0];
    ele[21][0] != ele[30][0];
    ele[21][0] != ele[31][0];
    ele[21][0] != ele[32][0];
    ele[21][0] != ele[33][0];
    ele[21][0] != ele[34][0];
    ele[21][0] != ele[35][0];
    ele[21][1] != ele[21][10];
    ele[21][1] != ele[21][11];
    ele[21][1] != ele[21][12];
    ele[21][1] != ele[21][13];
    ele[21][1] != ele[21][14];
    ele[21][1] != ele[21][15];
    ele[21][1] != ele[21][16];
    ele[21][1] != ele[21][17];
    ele[21][1] != ele[21][18];
    ele[21][1] != ele[21][19];
    ele[21][1] != ele[21][2];
    ele[21][1] != ele[21][20];
    ele[21][1] != ele[21][21];
    ele[21][1] != ele[21][22];
    ele[21][1] != ele[21][23];
    ele[21][1] != ele[21][24];
    ele[21][1] != ele[21][25];
    ele[21][1] != ele[21][26];
    ele[21][1] != ele[21][27];
    ele[21][1] != ele[21][28];
    ele[21][1] != ele[21][29];
    ele[21][1] != ele[21][3];
    ele[21][1] != ele[21][30];
    ele[21][1] != ele[21][31];
    ele[21][1] != ele[21][32];
    ele[21][1] != ele[21][33];
    ele[21][1] != ele[21][34];
    ele[21][1] != ele[21][35];
    ele[21][1] != ele[21][4];
    ele[21][1] != ele[21][5];
    ele[21][1] != ele[21][6];
    ele[21][1] != ele[21][7];
    ele[21][1] != ele[21][8];
    ele[21][1] != ele[21][9];
    ele[21][1] != ele[22][0];
    ele[21][1] != ele[22][1];
    ele[21][1] != ele[22][2];
    ele[21][1] != ele[22][3];
    ele[21][1] != ele[22][4];
    ele[21][1] != ele[22][5];
    ele[21][1] != ele[23][0];
    ele[21][1] != ele[23][1];
    ele[21][1] != ele[23][2];
    ele[21][1] != ele[23][3];
    ele[21][1] != ele[23][4];
    ele[21][1] != ele[23][5];
    ele[21][1] != ele[24][1];
    ele[21][1] != ele[25][1];
    ele[21][1] != ele[26][1];
    ele[21][1] != ele[27][1];
    ele[21][1] != ele[28][1];
    ele[21][1] != ele[29][1];
    ele[21][1] != ele[30][1];
    ele[21][1] != ele[31][1];
    ele[21][1] != ele[32][1];
    ele[21][1] != ele[33][1];
    ele[21][1] != ele[34][1];
    ele[21][1] != ele[35][1];
    ele[21][10] != ele[21][11];
    ele[21][10] != ele[21][12];
    ele[21][10] != ele[21][13];
    ele[21][10] != ele[21][14];
    ele[21][10] != ele[21][15];
    ele[21][10] != ele[21][16];
    ele[21][10] != ele[21][17];
    ele[21][10] != ele[21][18];
    ele[21][10] != ele[21][19];
    ele[21][10] != ele[21][20];
    ele[21][10] != ele[21][21];
    ele[21][10] != ele[21][22];
    ele[21][10] != ele[21][23];
    ele[21][10] != ele[21][24];
    ele[21][10] != ele[21][25];
    ele[21][10] != ele[21][26];
    ele[21][10] != ele[21][27];
    ele[21][10] != ele[21][28];
    ele[21][10] != ele[21][29];
    ele[21][10] != ele[21][30];
    ele[21][10] != ele[21][31];
    ele[21][10] != ele[21][32];
    ele[21][10] != ele[21][33];
    ele[21][10] != ele[21][34];
    ele[21][10] != ele[21][35];
    ele[21][10] != ele[22][10];
    ele[21][10] != ele[22][11];
    ele[21][10] != ele[22][6];
    ele[21][10] != ele[22][7];
    ele[21][10] != ele[22][8];
    ele[21][10] != ele[22][9];
    ele[21][10] != ele[23][10];
    ele[21][10] != ele[23][11];
    ele[21][10] != ele[23][6];
    ele[21][10] != ele[23][7];
    ele[21][10] != ele[23][8];
    ele[21][10] != ele[23][9];
    ele[21][10] != ele[24][10];
    ele[21][10] != ele[25][10];
    ele[21][10] != ele[26][10];
    ele[21][10] != ele[27][10];
    ele[21][10] != ele[28][10];
    ele[21][10] != ele[29][10];
    ele[21][10] != ele[30][10];
    ele[21][10] != ele[31][10];
    ele[21][10] != ele[32][10];
    ele[21][10] != ele[33][10];
    ele[21][10] != ele[34][10];
    ele[21][10] != ele[35][10];
    ele[21][11] != ele[21][12];
    ele[21][11] != ele[21][13];
    ele[21][11] != ele[21][14];
    ele[21][11] != ele[21][15];
    ele[21][11] != ele[21][16];
    ele[21][11] != ele[21][17];
    ele[21][11] != ele[21][18];
    ele[21][11] != ele[21][19];
    ele[21][11] != ele[21][20];
    ele[21][11] != ele[21][21];
    ele[21][11] != ele[21][22];
    ele[21][11] != ele[21][23];
    ele[21][11] != ele[21][24];
    ele[21][11] != ele[21][25];
    ele[21][11] != ele[21][26];
    ele[21][11] != ele[21][27];
    ele[21][11] != ele[21][28];
    ele[21][11] != ele[21][29];
    ele[21][11] != ele[21][30];
    ele[21][11] != ele[21][31];
    ele[21][11] != ele[21][32];
    ele[21][11] != ele[21][33];
    ele[21][11] != ele[21][34];
    ele[21][11] != ele[21][35];
    ele[21][11] != ele[22][10];
    ele[21][11] != ele[22][11];
    ele[21][11] != ele[22][6];
    ele[21][11] != ele[22][7];
    ele[21][11] != ele[22][8];
    ele[21][11] != ele[22][9];
    ele[21][11] != ele[23][10];
    ele[21][11] != ele[23][11];
    ele[21][11] != ele[23][6];
    ele[21][11] != ele[23][7];
    ele[21][11] != ele[23][8];
    ele[21][11] != ele[23][9];
    ele[21][11] != ele[24][11];
    ele[21][11] != ele[25][11];
    ele[21][11] != ele[26][11];
    ele[21][11] != ele[27][11];
    ele[21][11] != ele[28][11];
    ele[21][11] != ele[29][11];
    ele[21][11] != ele[30][11];
    ele[21][11] != ele[31][11];
    ele[21][11] != ele[32][11];
    ele[21][11] != ele[33][11];
    ele[21][11] != ele[34][11];
    ele[21][11] != ele[35][11];
    ele[21][12] != ele[21][13];
    ele[21][12] != ele[21][14];
    ele[21][12] != ele[21][15];
    ele[21][12] != ele[21][16];
    ele[21][12] != ele[21][17];
    ele[21][12] != ele[21][18];
    ele[21][12] != ele[21][19];
    ele[21][12] != ele[21][20];
    ele[21][12] != ele[21][21];
    ele[21][12] != ele[21][22];
    ele[21][12] != ele[21][23];
    ele[21][12] != ele[21][24];
    ele[21][12] != ele[21][25];
    ele[21][12] != ele[21][26];
    ele[21][12] != ele[21][27];
    ele[21][12] != ele[21][28];
    ele[21][12] != ele[21][29];
    ele[21][12] != ele[21][30];
    ele[21][12] != ele[21][31];
    ele[21][12] != ele[21][32];
    ele[21][12] != ele[21][33];
    ele[21][12] != ele[21][34];
    ele[21][12] != ele[21][35];
    ele[21][12] != ele[22][12];
    ele[21][12] != ele[22][13];
    ele[21][12] != ele[22][14];
    ele[21][12] != ele[22][15];
    ele[21][12] != ele[22][16];
    ele[21][12] != ele[22][17];
    ele[21][12] != ele[23][12];
    ele[21][12] != ele[23][13];
    ele[21][12] != ele[23][14];
    ele[21][12] != ele[23][15];
    ele[21][12] != ele[23][16];
    ele[21][12] != ele[23][17];
    ele[21][12] != ele[24][12];
    ele[21][12] != ele[25][12];
    ele[21][12] != ele[26][12];
    ele[21][12] != ele[27][12];
    ele[21][12] != ele[28][12];
    ele[21][12] != ele[29][12];
    ele[21][12] != ele[30][12];
    ele[21][12] != ele[31][12];
    ele[21][12] != ele[32][12];
    ele[21][12] != ele[33][12];
    ele[21][12] != ele[34][12];
    ele[21][12] != ele[35][12];
    ele[21][13] != ele[21][14];
    ele[21][13] != ele[21][15];
    ele[21][13] != ele[21][16];
    ele[21][13] != ele[21][17];
    ele[21][13] != ele[21][18];
    ele[21][13] != ele[21][19];
    ele[21][13] != ele[21][20];
    ele[21][13] != ele[21][21];
    ele[21][13] != ele[21][22];
    ele[21][13] != ele[21][23];
    ele[21][13] != ele[21][24];
    ele[21][13] != ele[21][25];
    ele[21][13] != ele[21][26];
    ele[21][13] != ele[21][27];
    ele[21][13] != ele[21][28];
    ele[21][13] != ele[21][29];
    ele[21][13] != ele[21][30];
    ele[21][13] != ele[21][31];
    ele[21][13] != ele[21][32];
    ele[21][13] != ele[21][33];
    ele[21][13] != ele[21][34];
    ele[21][13] != ele[21][35];
    ele[21][13] != ele[22][12];
    ele[21][13] != ele[22][13];
    ele[21][13] != ele[22][14];
    ele[21][13] != ele[22][15];
    ele[21][13] != ele[22][16];
    ele[21][13] != ele[22][17];
    ele[21][13] != ele[23][12];
    ele[21][13] != ele[23][13];
    ele[21][13] != ele[23][14];
    ele[21][13] != ele[23][15];
    ele[21][13] != ele[23][16];
    ele[21][13] != ele[23][17];
    ele[21][13] != ele[24][13];
    ele[21][13] != ele[25][13];
    ele[21][13] != ele[26][13];
    ele[21][13] != ele[27][13];
    ele[21][13] != ele[28][13];
    ele[21][13] != ele[29][13];
    ele[21][13] != ele[30][13];
    ele[21][13] != ele[31][13];
    ele[21][13] != ele[32][13];
    ele[21][13] != ele[33][13];
    ele[21][13] != ele[34][13];
    ele[21][13] != ele[35][13];
    ele[21][14] != ele[21][15];
    ele[21][14] != ele[21][16];
    ele[21][14] != ele[21][17];
    ele[21][14] != ele[21][18];
    ele[21][14] != ele[21][19];
    ele[21][14] != ele[21][20];
    ele[21][14] != ele[21][21];
    ele[21][14] != ele[21][22];
    ele[21][14] != ele[21][23];
    ele[21][14] != ele[21][24];
    ele[21][14] != ele[21][25];
    ele[21][14] != ele[21][26];
    ele[21][14] != ele[21][27];
    ele[21][14] != ele[21][28];
    ele[21][14] != ele[21][29];
    ele[21][14] != ele[21][30];
    ele[21][14] != ele[21][31];
    ele[21][14] != ele[21][32];
    ele[21][14] != ele[21][33];
    ele[21][14] != ele[21][34];
    ele[21][14] != ele[21][35];
    ele[21][14] != ele[22][12];
    ele[21][14] != ele[22][13];
    ele[21][14] != ele[22][14];
    ele[21][14] != ele[22][15];
    ele[21][14] != ele[22][16];
    ele[21][14] != ele[22][17];
    ele[21][14] != ele[23][12];
    ele[21][14] != ele[23][13];
    ele[21][14] != ele[23][14];
    ele[21][14] != ele[23][15];
    ele[21][14] != ele[23][16];
    ele[21][14] != ele[23][17];
    ele[21][14] != ele[24][14];
    ele[21][14] != ele[25][14];
    ele[21][14] != ele[26][14];
    ele[21][14] != ele[27][14];
    ele[21][14] != ele[28][14];
    ele[21][14] != ele[29][14];
    ele[21][14] != ele[30][14];
    ele[21][14] != ele[31][14];
    ele[21][14] != ele[32][14];
    ele[21][14] != ele[33][14];
    ele[21][14] != ele[34][14];
    ele[21][14] != ele[35][14];
    ele[21][15] != ele[21][16];
    ele[21][15] != ele[21][17];
    ele[21][15] != ele[21][18];
    ele[21][15] != ele[21][19];
    ele[21][15] != ele[21][20];
    ele[21][15] != ele[21][21];
    ele[21][15] != ele[21][22];
    ele[21][15] != ele[21][23];
    ele[21][15] != ele[21][24];
    ele[21][15] != ele[21][25];
    ele[21][15] != ele[21][26];
    ele[21][15] != ele[21][27];
    ele[21][15] != ele[21][28];
    ele[21][15] != ele[21][29];
    ele[21][15] != ele[21][30];
    ele[21][15] != ele[21][31];
    ele[21][15] != ele[21][32];
    ele[21][15] != ele[21][33];
    ele[21][15] != ele[21][34];
    ele[21][15] != ele[21][35];
    ele[21][15] != ele[22][12];
    ele[21][15] != ele[22][13];
    ele[21][15] != ele[22][14];
    ele[21][15] != ele[22][15];
    ele[21][15] != ele[22][16];
    ele[21][15] != ele[22][17];
    ele[21][15] != ele[23][12];
    ele[21][15] != ele[23][13];
    ele[21][15] != ele[23][14];
    ele[21][15] != ele[23][15];
    ele[21][15] != ele[23][16];
    ele[21][15] != ele[23][17];
    ele[21][15] != ele[24][15];
    ele[21][15] != ele[25][15];
    ele[21][15] != ele[26][15];
    ele[21][15] != ele[27][15];
    ele[21][15] != ele[28][15];
    ele[21][15] != ele[29][15];
    ele[21][15] != ele[30][15];
    ele[21][15] != ele[31][15];
    ele[21][15] != ele[32][15];
    ele[21][15] != ele[33][15];
    ele[21][15] != ele[34][15];
    ele[21][15] != ele[35][15];
    ele[21][16] != ele[21][17];
    ele[21][16] != ele[21][18];
    ele[21][16] != ele[21][19];
    ele[21][16] != ele[21][20];
    ele[21][16] != ele[21][21];
    ele[21][16] != ele[21][22];
    ele[21][16] != ele[21][23];
    ele[21][16] != ele[21][24];
    ele[21][16] != ele[21][25];
    ele[21][16] != ele[21][26];
    ele[21][16] != ele[21][27];
    ele[21][16] != ele[21][28];
    ele[21][16] != ele[21][29];
    ele[21][16] != ele[21][30];
    ele[21][16] != ele[21][31];
    ele[21][16] != ele[21][32];
    ele[21][16] != ele[21][33];
    ele[21][16] != ele[21][34];
    ele[21][16] != ele[21][35];
    ele[21][16] != ele[22][12];
    ele[21][16] != ele[22][13];
    ele[21][16] != ele[22][14];
    ele[21][16] != ele[22][15];
    ele[21][16] != ele[22][16];
    ele[21][16] != ele[22][17];
    ele[21][16] != ele[23][12];
    ele[21][16] != ele[23][13];
    ele[21][16] != ele[23][14];
    ele[21][16] != ele[23][15];
    ele[21][16] != ele[23][16];
    ele[21][16] != ele[23][17];
    ele[21][16] != ele[24][16];
    ele[21][16] != ele[25][16];
    ele[21][16] != ele[26][16];
    ele[21][16] != ele[27][16];
    ele[21][16] != ele[28][16];
    ele[21][16] != ele[29][16];
    ele[21][16] != ele[30][16];
    ele[21][16] != ele[31][16];
    ele[21][16] != ele[32][16];
    ele[21][16] != ele[33][16];
    ele[21][16] != ele[34][16];
    ele[21][16] != ele[35][16];
    ele[21][17] != ele[21][18];
    ele[21][17] != ele[21][19];
    ele[21][17] != ele[21][20];
    ele[21][17] != ele[21][21];
    ele[21][17] != ele[21][22];
    ele[21][17] != ele[21][23];
    ele[21][17] != ele[21][24];
    ele[21][17] != ele[21][25];
    ele[21][17] != ele[21][26];
    ele[21][17] != ele[21][27];
    ele[21][17] != ele[21][28];
    ele[21][17] != ele[21][29];
    ele[21][17] != ele[21][30];
    ele[21][17] != ele[21][31];
    ele[21][17] != ele[21][32];
    ele[21][17] != ele[21][33];
    ele[21][17] != ele[21][34];
    ele[21][17] != ele[21][35];
    ele[21][17] != ele[22][12];
    ele[21][17] != ele[22][13];
    ele[21][17] != ele[22][14];
    ele[21][17] != ele[22][15];
    ele[21][17] != ele[22][16];
    ele[21][17] != ele[22][17];
    ele[21][17] != ele[23][12];
    ele[21][17] != ele[23][13];
    ele[21][17] != ele[23][14];
    ele[21][17] != ele[23][15];
    ele[21][17] != ele[23][16];
    ele[21][17] != ele[23][17];
    ele[21][17] != ele[24][17];
    ele[21][17] != ele[25][17];
    ele[21][17] != ele[26][17];
    ele[21][17] != ele[27][17];
    ele[21][17] != ele[28][17];
    ele[21][17] != ele[29][17];
    ele[21][17] != ele[30][17];
    ele[21][17] != ele[31][17];
    ele[21][17] != ele[32][17];
    ele[21][17] != ele[33][17];
    ele[21][17] != ele[34][17];
    ele[21][17] != ele[35][17];
    ele[21][18] != ele[21][19];
    ele[21][18] != ele[21][20];
    ele[21][18] != ele[21][21];
    ele[21][18] != ele[21][22];
    ele[21][18] != ele[21][23];
    ele[21][18] != ele[21][24];
    ele[21][18] != ele[21][25];
    ele[21][18] != ele[21][26];
    ele[21][18] != ele[21][27];
    ele[21][18] != ele[21][28];
    ele[21][18] != ele[21][29];
    ele[21][18] != ele[21][30];
    ele[21][18] != ele[21][31];
    ele[21][18] != ele[21][32];
    ele[21][18] != ele[21][33];
    ele[21][18] != ele[21][34];
    ele[21][18] != ele[21][35];
    ele[21][18] != ele[22][18];
    ele[21][18] != ele[22][19];
    ele[21][18] != ele[22][20];
    ele[21][18] != ele[22][21];
    ele[21][18] != ele[22][22];
    ele[21][18] != ele[22][23];
    ele[21][18] != ele[23][18];
    ele[21][18] != ele[23][19];
    ele[21][18] != ele[23][20];
    ele[21][18] != ele[23][21];
    ele[21][18] != ele[23][22];
    ele[21][18] != ele[23][23];
    ele[21][18] != ele[24][18];
    ele[21][18] != ele[25][18];
    ele[21][18] != ele[26][18];
    ele[21][18] != ele[27][18];
    ele[21][18] != ele[28][18];
    ele[21][18] != ele[29][18];
    ele[21][18] != ele[30][18];
    ele[21][18] != ele[31][18];
    ele[21][18] != ele[32][18];
    ele[21][18] != ele[33][18];
    ele[21][18] != ele[34][18];
    ele[21][18] != ele[35][18];
    ele[21][19] != ele[21][20];
    ele[21][19] != ele[21][21];
    ele[21][19] != ele[21][22];
    ele[21][19] != ele[21][23];
    ele[21][19] != ele[21][24];
    ele[21][19] != ele[21][25];
    ele[21][19] != ele[21][26];
    ele[21][19] != ele[21][27];
    ele[21][19] != ele[21][28];
    ele[21][19] != ele[21][29];
    ele[21][19] != ele[21][30];
    ele[21][19] != ele[21][31];
    ele[21][19] != ele[21][32];
    ele[21][19] != ele[21][33];
    ele[21][19] != ele[21][34];
    ele[21][19] != ele[21][35];
    ele[21][19] != ele[22][18];
    ele[21][19] != ele[22][19];
    ele[21][19] != ele[22][20];
    ele[21][19] != ele[22][21];
    ele[21][19] != ele[22][22];
    ele[21][19] != ele[22][23];
    ele[21][19] != ele[23][18];
    ele[21][19] != ele[23][19];
    ele[21][19] != ele[23][20];
    ele[21][19] != ele[23][21];
    ele[21][19] != ele[23][22];
    ele[21][19] != ele[23][23];
    ele[21][19] != ele[24][19];
    ele[21][19] != ele[25][19];
    ele[21][19] != ele[26][19];
    ele[21][19] != ele[27][19];
    ele[21][19] != ele[28][19];
    ele[21][19] != ele[29][19];
    ele[21][19] != ele[30][19];
    ele[21][19] != ele[31][19];
    ele[21][19] != ele[32][19];
    ele[21][19] != ele[33][19];
    ele[21][19] != ele[34][19];
    ele[21][19] != ele[35][19];
    ele[21][2] != ele[21][10];
    ele[21][2] != ele[21][11];
    ele[21][2] != ele[21][12];
    ele[21][2] != ele[21][13];
    ele[21][2] != ele[21][14];
    ele[21][2] != ele[21][15];
    ele[21][2] != ele[21][16];
    ele[21][2] != ele[21][17];
    ele[21][2] != ele[21][18];
    ele[21][2] != ele[21][19];
    ele[21][2] != ele[21][20];
    ele[21][2] != ele[21][21];
    ele[21][2] != ele[21][22];
    ele[21][2] != ele[21][23];
    ele[21][2] != ele[21][24];
    ele[21][2] != ele[21][25];
    ele[21][2] != ele[21][26];
    ele[21][2] != ele[21][27];
    ele[21][2] != ele[21][28];
    ele[21][2] != ele[21][29];
    ele[21][2] != ele[21][3];
    ele[21][2] != ele[21][30];
    ele[21][2] != ele[21][31];
    ele[21][2] != ele[21][32];
    ele[21][2] != ele[21][33];
    ele[21][2] != ele[21][34];
    ele[21][2] != ele[21][35];
    ele[21][2] != ele[21][4];
    ele[21][2] != ele[21][5];
    ele[21][2] != ele[21][6];
    ele[21][2] != ele[21][7];
    ele[21][2] != ele[21][8];
    ele[21][2] != ele[21][9];
    ele[21][2] != ele[22][0];
    ele[21][2] != ele[22][1];
    ele[21][2] != ele[22][2];
    ele[21][2] != ele[22][3];
    ele[21][2] != ele[22][4];
    ele[21][2] != ele[22][5];
    ele[21][2] != ele[23][0];
    ele[21][2] != ele[23][1];
    ele[21][2] != ele[23][2];
    ele[21][2] != ele[23][3];
    ele[21][2] != ele[23][4];
    ele[21][2] != ele[23][5];
    ele[21][2] != ele[24][2];
    ele[21][2] != ele[25][2];
    ele[21][2] != ele[26][2];
    ele[21][2] != ele[27][2];
    ele[21][2] != ele[28][2];
    ele[21][2] != ele[29][2];
    ele[21][2] != ele[30][2];
    ele[21][2] != ele[31][2];
    ele[21][2] != ele[32][2];
    ele[21][2] != ele[33][2];
    ele[21][2] != ele[34][2];
    ele[21][2] != ele[35][2];
    ele[21][20] != ele[21][21];
    ele[21][20] != ele[21][22];
    ele[21][20] != ele[21][23];
    ele[21][20] != ele[21][24];
    ele[21][20] != ele[21][25];
    ele[21][20] != ele[21][26];
    ele[21][20] != ele[21][27];
    ele[21][20] != ele[21][28];
    ele[21][20] != ele[21][29];
    ele[21][20] != ele[21][30];
    ele[21][20] != ele[21][31];
    ele[21][20] != ele[21][32];
    ele[21][20] != ele[21][33];
    ele[21][20] != ele[21][34];
    ele[21][20] != ele[21][35];
    ele[21][20] != ele[22][18];
    ele[21][20] != ele[22][19];
    ele[21][20] != ele[22][20];
    ele[21][20] != ele[22][21];
    ele[21][20] != ele[22][22];
    ele[21][20] != ele[22][23];
    ele[21][20] != ele[23][18];
    ele[21][20] != ele[23][19];
    ele[21][20] != ele[23][20];
    ele[21][20] != ele[23][21];
    ele[21][20] != ele[23][22];
    ele[21][20] != ele[23][23];
    ele[21][20] != ele[24][20];
    ele[21][20] != ele[25][20];
    ele[21][20] != ele[26][20];
    ele[21][20] != ele[27][20];
    ele[21][20] != ele[28][20];
    ele[21][20] != ele[29][20];
    ele[21][20] != ele[30][20];
    ele[21][20] != ele[31][20];
    ele[21][20] != ele[32][20];
    ele[21][20] != ele[33][20];
    ele[21][20] != ele[34][20];
    ele[21][20] != ele[35][20];
    ele[21][21] != ele[21][22];
    ele[21][21] != ele[21][23];
    ele[21][21] != ele[21][24];
    ele[21][21] != ele[21][25];
    ele[21][21] != ele[21][26];
    ele[21][21] != ele[21][27];
    ele[21][21] != ele[21][28];
    ele[21][21] != ele[21][29];
    ele[21][21] != ele[21][30];
    ele[21][21] != ele[21][31];
    ele[21][21] != ele[21][32];
    ele[21][21] != ele[21][33];
    ele[21][21] != ele[21][34];
    ele[21][21] != ele[21][35];
    ele[21][21] != ele[22][18];
    ele[21][21] != ele[22][19];
    ele[21][21] != ele[22][20];
    ele[21][21] != ele[22][21];
    ele[21][21] != ele[22][22];
    ele[21][21] != ele[22][23];
    ele[21][21] != ele[23][18];
    ele[21][21] != ele[23][19];
    ele[21][21] != ele[23][20];
    ele[21][21] != ele[23][21];
    ele[21][21] != ele[23][22];
    ele[21][21] != ele[23][23];
    ele[21][21] != ele[24][21];
    ele[21][21] != ele[25][21];
    ele[21][21] != ele[26][21];
    ele[21][21] != ele[27][21];
    ele[21][21] != ele[28][21];
    ele[21][21] != ele[29][21];
    ele[21][21] != ele[30][21];
    ele[21][21] != ele[31][21];
    ele[21][21] != ele[32][21];
    ele[21][21] != ele[33][21];
    ele[21][21] != ele[34][21];
    ele[21][21] != ele[35][21];
    ele[21][22] != ele[21][23];
    ele[21][22] != ele[21][24];
    ele[21][22] != ele[21][25];
    ele[21][22] != ele[21][26];
    ele[21][22] != ele[21][27];
    ele[21][22] != ele[21][28];
    ele[21][22] != ele[21][29];
    ele[21][22] != ele[21][30];
    ele[21][22] != ele[21][31];
    ele[21][22] != ele[21][32];
    ele[21][22] != ele[21][33];
    ele[21][22] != ele[21][34];
    ele[21][22] != ele[21][35];
    ele[21][22] != ele[22][18];
    ele[21][22] != ele[22][19];
    ele[21][22] != ele[22][20];
    ele[21][22] != ele[22][21];
    ele[21][22] != ele[22][22];
    ele[21][22] != ele[22][23];
    ele[21][22] != ele[23][18];
    ele[21][22] != ele[23][19];
    ele[21][22] != ele[23][20];
    ele[21][22] != ele[23][21];
    ele[21][22] != ele[23][22];
    ele[21][22] != ele[23][23];
    ele[21][22] != ele[24][22];
    ele[21][22] != ele[25][22];
    ele[21][22] != ele[26][22];
    ele[21][22] != ele[27][22];
    ele[21][22] != ele[28][22];
    ele[21][22] != ele[29][22];
    ele[21][22] != ele[30][22];
    ele[21][22] != ele[31][22];
    ele[21][22] != ele[32][22];
    ele[21][22] != ele[33][22];
    ele[21][22] != ele[34][22];
    ele[21][22] != ele[35][22];
    ele[21][23] != ele[21][24];
    ele[21][23] != ele[21][25];
    ele[21][23] != ele[21][26];
    ele[21][23] != ele[21][27];
    ele[21][23] != ele[21][28];
    ele[21][23] != ele[21][29];
    ele[21][23] != ele[21][30];
    ele[21][23] != ele[21][31];
    ele[21][23] != ele[21][32];
    ele[21][23] != ele[21][33];
    ele[21][23] != ele[21][34];
    ele[21][23] != ele[21][35];
    ele[21][23] != ele[22][18];
    ele[21][23] != ele[22][19];
    ele[21][23] != ele[22][20];
    ele[21][23] != ele[22][21];
    ele[21][23] != ele[22][22];
    ele[21][23] != ele[22][23];
    ele[21][23] != ele[23][18];
    ele[21][23] != ele[23][19];
    ele[21][23] != ele[23][20];
    ele[21][23] != ele[23][21];
    ele[21][23] != ele[23][22];
    ele[21][23] != ele[23][23];
    ele[21][23] != ele[24][23];
    ele[21][23] != ele[25][23];
    ele[21][23] != ele[26][23];
    ele[21][23] != ele[27][23];
    ele[21][23] != ele[28][23];
    ele[21][23] != ele[29][23];
    ele[21][23] != ele[30][23];
    ele[21][23] != ele[31][23];
    ele[21][23] != ele[32][23];
    ele[21][23] != ele[33][23];
    ele[21][23] != ele[34][23];
    ele[21][23] != ele[35][23];
    ele[21][24] != ele[21][25];
    ele[21][24] != ele[21][26];
    ele[21][24] != ele[21][27];
    ele[21][24] != ele[21][28];
    ele[21][24] != ele[21][29];
    ele[21][24] != ele[21][30];
    ele[21][24] != ele[21][31];
    ele[21][24] != ele[21][32];
    ele[21][24] != ele[21][33];
    ele[21][24] != ele[21][34];
    ele[21][24] != ele[21][35];
    ele[21][24] != ele[22][24];
    ele[21][24] != ele[22][25];
    ele[21][24] != ele[22][26];
    ele[21][24] != ele[22][27];
    ele[21][24] != ele[22][28];
    ele[21][24] != ele[22][29];
    ele[21][24] != ele[23][24];
    ele[21][24] != ele[23][25];
    ele[21][24] != ele[23][26];
    ele[21][24] != ele[23][27];
    ele[21][24] != ele[23][28];
    ele[21][24] != ele[23][29];
    ele[21][24] != ele[24][24];
    ele[21][24] != ele[25][24];
    ele[21][24] != ele[26][24];
    ele[21][24] != ele[27][24];
    ele[21][24] != ele[28][24];
    ele[21][24] != ele[29][24];
    ele[21][24] != ele[30][24];
    ele[21][24] != ele[31][24];
    ele[21][24] != ele[32][24];
    ele[21][24] != ele[33][24];
    ele[21][24] != ele[34][24];
    ele[21][24] != ele[35][24];
    ele[21][25] != ele[21][26];
    ele[21][25] != ele[21][27];
    ele[21][25] != ele[21][28];
    ele[21][25] != ele[21][29];
    ele[21][25] != ele[21][30];
    ele[21][25] != ele[21][31];
    ele[21][25] != ele[21][32];
    ele[21][25] != ele[21][33];
    ele[21][25] != ele[21][34];
    ele[21][25] != ele[21][35];
    ele[21][25] != ele[22][24];
    ele[21][25] != ele[22][25];
    ele[21][25] != ele[22][26];
    ele[21][25] != ele[22][27];
    ele[21][25] != ele[22][28];
    ele[21][25] != ele[22][29];
    ele[21][25] != ele[23][24];
    ele[21][25] != ele[23][25];
    ele[21][25] != ele[23][26];
    ele[21][25] != ele[23][27];
    ele[21][25] != ele[23][28];
    ele[21][25] != ele[23][29];
    ele[21][25] != ele[24][25];
    ele[21][25] != ele[25][25];
    ele[21][25] != ele[26][25];
    ele[21][25] != ele[27][25];
    ele[21][25] != ele[28][25];
    ele[21][25] != ele[29][25];
    ele[21][25] != ele[30][25];
    ele[21][25] != ele[31][25];
    ele[21][25] != ele[32][25];
    ele[21][25] != ele[33][25];
    ele[21][25] != ele[34][25];
    ele[21][25] != ele[35][25];
    ele[21][26] != ele[21][27];
    ele[21][26] != ele[21][28];
    ele[21][26] != ele[21][29];
    ele[21][26] != ele[21][30];
    ele[21][26] != ele[21][31];
    ele[21][26] != ele[21][32];
    ele[21][26] != ele[21][33];
    ele[21][26] != ele[21][34];
    ele[21][26] != ele[21][35];
    ele[21][26] != ele[22][24];
    ele[21][26] != ele[22][25];
    ele[21][26] != ele[22][26];
    ele[21][26] != ele[22][27];
    ele[21][26] != ele[22][28];
    ele[21][26] != ele[22][29];
    ele[21][26] != ele[23][24];
    ele[21][26] != ele[23][25];
    ele[21][26] != ele[23][26];
    ele[21][26] != ele[23][27];
    ele[21][26] != ele[23][28];
    ele[21][26] != ele[23][29];
    ele[21][26] != ele[24][26];
    ele[21][26] != ele[25][26];
    ele[21][26] != ele[26][26];
    ele[21][26] != ele[27][26];
    ele[21][26] != ele[28][26];
    ele[21][26] != ele[29][26];
    ele[21][26] != ele[30][26];
    ele[21][26] != ele[31][26];
    ele[21][26] != ele[32][26];
    ele[21][26] != ele[33][26];
    ele[21][26] != ele[34][26];
    ele[21][26] != ele[35][26];
    ele[21][27] != ele[21][28];
    ele[21][27] != ele[21][29];
    ele[21][27] != ele[21][30];
    ele[21][27] != ele[21][31];
    ele[21][27] != ele[21][32];
    ele[21][27] != ele[21][33];
    ele[21][27] != ele[21][34];
    ele[21][27] != ele[21][35];
    ele[21][27] != ele[22][24];
    ele[21][27] != ele[22][25];
    ele[21][27] != ele[22][26];
    ele[21][27] != ele[22][27];
    ele[21][27] != ele[22][28];
    ele[21][27] != ele[22][29];
    ele[21][27] != ele[23][24];
    ele[21][27] != ele[23][25];
    ele[21][27] != ele[23][26];
    ele[21][27] != ele[23][27];
    ele[21][27] != ele[23][28];
    ele[21][27] != ele[23][29];
    ele[21][27] != ele[24][27];
    ele[21][27] != ele[25][27];
    ele[21][27] != ele[26][27];
    ele[21][27] != ele[27][27];
    ele[21][27] != ele[28][27];
    ele[21][27] != ele[29][27];
    ele[21][27] != ele[30][27];
    ele[21][27] != ele[31][27];
    ele[21][27] != ele[32][27];
    ele[21][27] != ele[33][27];
    ele[21][27] != ele[34][27];
    ele[21][27] != ele[35][27];
    ele[21][28] != ele[21][29];
    ele[21][28] != ele[21][30];
    ele[21][28] != ele[21][31];
    ele[21][28] != ele[21][32];
    ele[21][28] != ele[21][33];
    ele[21][28] != ele[21][34];
    ele[21][28] != ele[21][35];
    ele[21][28] != ele[22][24];
    ele[21][28] != ele[22][25];
    ele[21][28] != ele[22][26];
    ele[21][28] != ele[22][27];
    ele[21][28] != ele[22][28];
    ele[21][28] != ele[22][29];
    ele[21][28] != ele[23][24];
    ele[21][28] != ele[23][25];
    ele[21][28] != ele[23][26];
    ele[21][28] != ele[23][27];
    ele[21][28] != ele[23][28];
    ele[21][28] != ele[23][29];
    ele[21][28] != ele[24][28];
    ele[21][28] != ele[25][28];
    ele[21][28] != ele[26][28];
    ele[21][28] != ele[27][28];
    ele[21][28] != ele[28][28];
    ele[21][28] != ele[29][28];
    ele[21][28] != ele[30][28];
    ele[21][28] != ele[31][28];
    ele[21][28] != ele[32][28];
    ele[21][28] != ele[33][28];
    ele[21][28] != ele[34][28];
    ele[21][28] != ele[35][28];
    ele[21][29] != ele[21][30];
    ele[21][29] != ele[21][31];
    ele[21][29] != ele[21][32];
    ele[21][29] != ele[21][33];
    ele[21][29] != ele[21][34];
    ele[21][29] != ele[21][35];
    ele[21][29] != ele[22][24];
    ele[21][29] != ele[22][25];
    ele[21][29] != ele[22][26];
    ele[21][29] != ele[22][27];
    ele[21][29] != ele[22][28];
    ele[21][29] != ele[22][29];
    ele[21][29] != ele[23][24];
    ele[21][29] != ele[23][25];
    ele[21][29] != ele[23][26];
    ele[21][29] != ele[23][27];
    ele[21][29] != ele[23][28];
    ele[21][29] != ele[23][29];
    ele[21][29] != ele[24][29];
    ele[21][29] != ele[25][29];
    ele[21][29] != ele[26][29];
    ele[21][29] != ele[27][29];
    ele[21][29] != ele[28][29];
    ele[21][29] != ele[29][29];
    ele[21][29] != ele[30][29];
    ele[21][29] != ele[31][29];
    ele[21][29] != ele[32][29];
    ele[21][29] != ele[33][29];
    ele[21][29] != ele[34][29];
    ele[21][29] != ele[35][29];
    ele[21][3] != ele[21][10];
    ele[21][3] != ele[21][11];
    ele[21][3] != ele[21][12];
    ele[21][3] != ele[21][13];
    ele[21][3] != ele[21][14];
    ele[21][3] != ele[21][15];
    ele[21][3] != ele[21][16];
    ele[21][3] != ele[21][17];
    ele[21][3] != ele[21][18];
    ele[21][3] != ele[21][19];
    ele[21][3] != ele[21][20];
    ele[21][3] != ele[21][21];
    ele[21][3] != ele[21][22];
    ele[21][3] != ele[21][23];
    ele[21][3] != ele[21][24];
    ele[21][3] != ele[21][25];
    ele[21][3] != ele[21][26];
    ele[21][3] != ele[21][27];
    ele[21][3] != ele[21][28];
    ele[21][3] != ele[21][29];
    ele[21][3] != ele[21][30];
    ele[21][3] != ele[21][31];
    ele[21][3] != ele[21][32];
    ele[21][3] != ele[21][33];
    ele[21][3] != ele[21][34];
    ele[21][3] != ele[21][35];
    ele[21][3] != ele[21][4];
    ele[21][3] != ele[21][5];
    ele[21][3] != ele[21][6];
    ele[21][3] != ele[21][7];
    ele[21][3] != ele[21][8];
    ele[21][3] != ele[21][9];
    ele[21][3] != ele[22][0];
    ele[21][3] != ele[22][1];
    ele[21][3] != ele[22][2];
    ele[21][3] != ele[22][3];
    ele[21][3] != ele[22][4];
    ele[21][3] != ele[22][5];
    ele[21][3] != ele[23][0];
    ele[21][3] != ele[23][1];
    ele[21][3] != ele[23][2];
    ele[21][3] != ele[23][3];
    ele[21][3] != ele[23][4];
    ele[21][3] != ele[23][5];
    ele[21][3] != ele[24][3];
    ele[21][3] != ele[25][3];
    ele[21][3] != ele[26][3];
    ele[21][3] != ele[27][3];
    ele[21][3] != ele[28][3];
    ele[21][3] != ele[29][3];
    ele[21][3] != ele[30][3];
    ele[21][3] != ele[31][3];
    ele[21][3] != ele[32][3];
    ele[21][3] != ele[33][3];
    ele[21][3] != ele[34][3];
    ele[21][3] != ele[35][3];
    ele[21][30] != ele[21][31];
    ele[21][30] != ele[21][32];
    ele[21][30] != ele[21][33];
    ele[21][30] != ele[21][34];
    ele[21][30] != ele[21][35];
    ele[21][30] != ele[22][30];
    ele[21][30] != ele[22][31];
    ele[21][30] != ele[22][32];
    ele[21][30] != ele[22][33];
    ele[21][30] != ele[22][34];
    ele[21][30] != ele[22][35];
    ele[21][30] != ele[23][30];
    ele[21][30] != ele[23][31];
    ele[21][30] != ele[23][32];
    ele[21][30] != ele[23][33];
    ele[21][30] != ele[23][34];
    ele[21][30] != ele[23][35];
    ele[21][30] != ele[24][30];
    ele[21][30] != ele[25][30];
    ele[21][30] != ele[26][30];
    ele[21][30] != ele[27][30];
    ele[21][30] != ele[28][30];
    ele[21][30] != ele[29][30];
    ele[21][30] != ele[30][30];
    ele[21][30] != ele[31][30];
    ele[21][30] != ele[32][30];
    ele[21][30] != ele[33][30];
    ele[21][30] != ele[34][30];
    ele[21][30] != ele[35][30];
    ele[21][31] != ele[21][32];
    ele[21][31] != ele[21][33];
    ele[21][31] != ele[21][34];
    ele[21][31] != ele[21][35];
    ele[21][31] != ele[22][30];
    ele[21][31] != ele[22][31];
    ele[21][31] != ele[22][32];
    ele[21][31] != ele[22][33];
    ele[21][31] != ele[22][34];
    ele[21][31] != ele[22][35];
    ele[21][31] != ele[23][30];
    ele[21][31] != ele[23][31];
    ele[21][31] != ele[23][32];
    ele[21][31] != ele[23][33];
    ele[21][31] != ele[23][34];
    ele[21][31] != ele[23][35];
    ele[21][31] != ele[24][31];
    ele[21][31] != ele[25][31];
    ele[21][31] != ele[26][31];
    ele[21][31] != ele[27][31];
    ele[21][31] != ele[28][31];
    ele[21][31] != ele[29][31];
    ele[21][31] != ele[30][31];
    ele[21][31] != ele[31][31];
    ele[21][31] != ele[32][31];
    ele[21][31] != ele[33][31];
    ele[21][31] != ele[34][31];
    ele[21][31] != ele[35][31];
    ele[21][32] != ele[21][33];
    ele[21][32] != ele[21][34];
    ele[21][32] != ele[21][35];
    ele[21][32] != ele[22][30];
    ele[21][32] != ele[22][31];
    ele[21][32] != ele[22][32];
    ele[21][32] != ele[22][33];
    ele[21][32] != ele[22][34];
    ele[21][32] != ele[22][35];
    ele[21][32] != ele[23][30];
    ele[21][32] != ele[23][31];
    ele[21][32] != ele[23][32];
    ele[21][32] != ele[23][33];
    ele[21][32] != ele[23][34];
    ele[21][32] != ele[23][35];
    ele[21][32] != ele[24][32];
    ele[21][32] != ele[25][32];
    ele[21][32] != ele[26][32];
    ele[21][32] != ele[27][32];
    ele[21][32] != ele[28][32];
    ele[21][32] != ele[29][32];
    ele[21][32] != ele[30][32];
    ele[21][32] != ele[31][32];
    ele[21][32] != ele[32][32];
    ele[21][32] != ele[33][32];
    ele[21][32] != ele[34][32];
    ele[21][32] != ele[35][32];
    ele[21][33] != ele[21][34];
    ele[21][33] != ele[21][35];
    ele[21][33] != ele[22][30];
    ele[21][33] != ele[22][31];
    ele[21][33] != ele[22][32];
    ele[21][33] != ele[22][33];
    ele[21][33] != ele[22][34];
    ele[21][33] != ele[22][35];
    ele[21][33] != ele[23][30];
    ele[21][33] != ele[23][31];
    ele[21][33] != ele[23][32];
    ele[21][33] != ele[23][33];
    ele[21][33] != ele[23][34];
    ele[21][33] != ele[23][35];
    ele[21][33] != ele[24][33];
    ele[21][33] != ele[25][33];
    ele[21][33] != ele[26][33];
    ele[21][33] != ele[27][33];
    ele[21][33] != ele[28][33];
    ele[21][33] != ele[29][33];
    ele[21][33] != ele[30][33];
    ele[21][33] != ele[31][33];
    ele[21][33] != ele[32][33];
    ele[21][33] != ele[33][33];
    ele[21][33] != ele[34][33];
    ele[21][33] != ele[35][33];
    ele[21][34] != ele[21][35];
    ele[21][34] != ele[22][30];
    ele[21][34] != ele[22][31];
    ele[21][34] != ele[22][32];
    ele[21][34] != ele[22][33];
    ele[21][34] != ele[22][34];
    ele[21][34] != ele[22][35];
    ele[21][34] != ele[23][30];
    ele[21][34] != ele[23][31];
    ele[21][34] != ele[23][32];
    ele[21][34] != ele[23][33];
    ele[21][34] != ele[23][34];
    ele[21][34] != ele[23][35];
    ele[21][34] != ele[24][34];
    ele[21][34] != ele[25][34];
    ele[21][34] != ele[26][34];
    ele[21][34] != ele[27][34];
    ele[21][34] != ele[28][34];
    ele[21][34] != ele[29][34];
    ele[21][34] != ele[30][34];
    ele[21][34] != ele[31][34];
    ele[21][34] != ele[32][34];
    ele[21][34] != ele[33][34];
    ele[21][34] != ele[34][34];
    ele[21][34] != ele[35][34];
    ele[21][35] != ele[22][30];
    ele[21][35] != ele[22][31];
    ele[21][35] != ele[22][32];
    ele[21][35] != ele[22][33];
    ele[21][35] != ele[22][34];
    ele[21][35] != ele[22][35];
    ele[21][35] != ele[23][30];
    ele[21][35] != ele[23][31];
    ele[21][35] != ele[23][32];
    ele[21][35] != ele[23][33];
    ele[21][35] != ele[23][34];
    ele[21][35] != ele[23][35];
    ele[21][35] != ele[24][35];
    ele[21][35] != ele[25][35];
    ele[21][35] != ele[26][35];
    ele[21][35] != ele[27][35];
    ele[21][35] != ele[28][35];
    ele[21][35] != ele[29][35];
    ele[21][35] != ele[30][35];
    ele[21][35] != ele[31][35];
    ele[21][35] != ele[32][35];
    ele[21][35] != ele[33][35];
    ele[21][35] != ele[34][35];
    ele[21][35] != ele[35][35];
    ele[21][4] != ele[21][10];
    ele[21][4] != ele[21][11];
    ele[21][4] != ele[21][12];
    ele[21][4] != ele[21][13];
    ele[21][4] != ele[21][14];
    ele[21][4] != ele[21][15];
    ele[21][4] != ele[21][16];
    ele[21][4] != ele[21][17];
    ele[21][4] != ele[21][18];
    ele[21][4] != ele[21][19];
    ele[21][4] != ele[21][20];
    ele[21][4] != ele[21][21];
    ele[21][4] != ele[21][22];
    ele[21][4] != ele[21][23];
    ele[21][4] != ele[21][24];
    ele[21][4] != ele[21][25];
    ele[21][4] != ele[21][26];
    ele[21][4] != ele[21][27];
    ele[21][4] != ele[21][28];
    ele[21][4] != ele[21][29];
    ele[21][4] != ele[21][30];
    ele[21][4] != ele[21][31];
    ele[21][4] != ele[21][32];
    ele[21][4] != ele[21][33];
    ele[21][4] != ele[21][34];
    ele[21][4] != ele[21][35];
    ele[21][4] != ele[21][5];
    ele[21][4] != ele[21][6];
    ele[21][4] != ele[21][7];
    ele[21][4] != ele[21][8];
    ele[21][4] != ele[21][9];
    ele[21][4] != ele[22][0];
    ele[21][4] != ele[22][1];
    ele[21][4] != ele[22][2];
    ele[21][4] != ele[22][3];
    ele[21][4] != ele[22][4];
    ele[21][4] != ele[22][5];
    ele[21][4] != ele[23][0];
    ele[21][4] != ele[23][1];
    ele[21][4] != ele[23][2];
    ele[21][4] != ele[23][3];
    ele[21][4] != ele[23][4];
    ele[21][4] != ele[23][5];
    ele[21][4] != ele[24][4];
    ele[21][4] != ele[25][4];
    ele[21][4] != ele[26][4];
    ele[21][4] != ele[27][4];
    ele[21][4] != ele[28][4];
    ele[21][4] != ele[29][4];
    ele[21][4] != ele[30][4];
    ele[21][4] != ele[31][4];
    ele[21][4] != ele[32][4];
    ele[21][4] != ele[33][4];
    ele[21][4] != ele[34][4];
    ele[21][4] != ele[35][4];
    ele[21][5] != ele[21][10];
    ele[21][5] != ele[21][11];
    ele[21][5] != ele[21][12];
    ele[21][5] != ele[21][13];
    ele[21][5] != ele[21][14];
    ele[21][5] != ele[21][15];
    ele[21][5] != ele[21][16];
    ele[21][5] != ele[21][17];
    ele[21][5] != ele[21][18];
    ele[21][5] != ele[21][19];
    ele[21][5] != ele[21][20];
    ele[21][5] != ele[21][21];
    ele[21][5] != ele[21][22];
    ele[21][5] != ele[21][23];
    ele[21][5] != ele[21][24];
    ele[21][5] != ele[21][25];
    ele[21][5] != ele[21][26];
    ele[21][5] != ele[21][27];
    ele[21][5] != ele[21][28];
    ele[21][5] != ele[21][29];
    ele[21][5] != ele[21][30];
    ele[21][5] != ele[21][31];
    ele[21][5] != ele[21][32];
    ele[21][5] != ele[21][33];
    ele[21][5] != ele[21][34];
    ele[21][5] != ele[21][35];
    ele[21][5] != ele[21][6];
    ele[21][5] != ele[21][7];
    ele[21][5] != ele[21][8];
    ele[21][5] != ele[21][9];
    ele[21][5] != ele[22][0];
    ele[21][5] != ele[22][1];
    ele[21][5] != ele[22][2];
    ele[21][5] != ele[22][3];
    ele[21][5] != ele[22][4];
    ele[21][5] != ele[22][5];
    ele[21][5] != ele[23][0];
    ele[21][5] != ele[23][1];
    ele[21][5] != ele[23][2];
    ele[21][5] != ele[23][3];
    ele[21][5] != ele[23][4];
    ele[21][5] != ele[23][5];
    ele[21][5] != ele[24][5];
    ele[21][5] != ele[25][5];
    ele[21][5] != ele[26][5];
    ele[21][5] != ele[27][5];
    ele[21][5] != ele[28][5];
    ele[21][5] != ele[29][5];
    ele[21][5] != ele[30][5];
    ele[21][5] != ele[31][5];
    ele[21][5] != ele[32][5];
    ele[21][5] != ele[33][5];
    ele[21][5] != ele[34][5];
    ele[21][5] != ele[35][5];
    ele[21][6] != ele[21][10];
    ele[21][6] != ele[21][11];
    ele[21][6] != ele[21][12];
    ele[21][6] != ele[21][13];
    ele[21][6] != ele[21][14];
    ele[21][6] != ele[21][15];
    ele[21][6] != ele[21][16];
    ele[21][6] != ele[21][17];
    ele[21][6] != ele[21][18];
    ele[21][6] != ele[21][19];
    ele[21][6] != ele[21][20];
    ele[21][6] != ele[21][21];
    ele[21][6] != ele[21][22];
    ele[21][6] != ele[21][23];
    ele[21][6] != ele[21][24];
    ele[21][6] != ele[21][25];
    ele[21][6] != ele[21][26];
    ele[21][6] != ele[21][27];
    ele[21][6] != ele[21][28];
    ele[21][6] != ele[21][29];
    ele[21][6] != ele[21][30];
    ele[21][6] != ele[21][31];
    ele[21][6] != ele[21][32];
    ele[21][6] != ele[21][33];
    ele[21][6] != ele[21][34];
    ele[21][6] != ele[21][35];
    ele[21][6] != ele[21][7];
    ele[21][6] != ele[21][8];
    ele[21][6] != ele[21][9];
    ele[21][6] != ele[22][10];
    ele[21][6] != ele[22][11];
    ele[21][6] != ele[22][6];
    ele[21][6] != ele[22][7];
    ele[21][6] != ele[22][8];
    ele[21][6] != ele[22][9];
    ele[21][6] != ele[23][10];
    ele[21][6] != ele[23][11];
    ele[21][6] != ele[23][6];
    ele[21][6] != ele[23][7];
    ele[21][6] != ele[23][8];
    ele[21][6] != ele[23][9];
    ele[21][6] != ele[24][6];
    ele[21][6] != ele[25][6];
    ele[21][6] != ele[26][6];
    ele[21][6] != ele[27][6];
    ele[21][6] != ele[28][6];
    ele[21][6] != ele[29][6];
    ele[21][6] != ele[30][6];
    ele[21][6] != ele[31][6];
    ele[21][6] != ele[32][6];
    ele[21][6] != ele[33][6];
    ele[21][6] != ele[34][6];
    ele[21][6] != ele[35][6];
    ele[21][7] != ele[21][10];
    ele[21][7] != ele[21][11];
    ele[21][7] != ele[21][12];
    ele[21][7] != ele[21][13];
    ele[21][7] != ele[21][14];
    ele[21][7] != ele[21][15];
    ele[21][7] != ele[21][16];
    ele[21][7] != ele[21][17];
    ele[21][7] != ele[21][18];
    ele[21][7] != ele[21][19];
    ele[21][7] != ele[21][20];
    ele[21][7] != ele[21][21];
    ele[21][7] != ele[21][22];
    ele[21][7] != ele[21][23];
    ele[21][7] != ele[21][24];
    ele[21][7] != ele[21][25];
    ele[21][7] != ele[21][26];
    ele[21][7] != ele[21][27];
    ele[21][7] != ele[21][28];
    ele[21][7] != ele[21][29];
    ele[21][7] != ele[21][30];
    ele[21][7] != ele[21][31];
    ele[21][7] != ele[21][32];
    ele[21][7] != ele[21][33];
    ele[21][7] != ele[21][34];
    ele[21][7] != ele[21][35];
    ele[21][7] != ele[21][8];
    ele[21][7] != ele[21][9];
    ele[21][7] != ele[22][10];
    ele[21][7] != ele[22][11];
    ele[21][7] != ele[22][6];
    ele[21][7] != ele[22][7];
    ele[21][7] != ele[22][8];
    ele[21][7] != ele[22][9];
    ele[21][7] != ele[23][10];
    ele[21][7] != ele[23][11];
    ele[21][7] != ele[23][6];
    ele[21][7] != ele[23][7];
    ele[21][7] != ele[23][8];
    ele[21][7] != ele[23][9];
    ele[21][7] != ele[24][7];
    ele[21][7] != ele[25][7];
    ele[21][7] != ele[26][7];
    ele[21][7] != ele[27][7];
    ele[21][7] != ele[28][7];
    ele[21][7] != ele[29][7];
    ele[21][7] != ele[30][7];
    ele[21][7] != ele[31][7];
    ele[21][7] != ele[32][7];
    ele[21][7] != ele[33][7];
    ele[21][7] != ele[34][7];
    ele[21][7] != ele[35][7];
    ele[21][8] != ele[21][10];
    ele[21][8] != ele[21][11];
    ele[21][8] != ele[21][12];
    ele[21][8] != ele[21][13];
    ele[21][8] != ele[21][14];
    ele[21][8] != ele[21][15];
    ele[21][8] != ele[21][16];
    ele[21][8] != ele[21][17];
    ele[21][8] != ele[21][18];
    ele[21][8] != ele[21][19];
    ele[21][8] != ele[21][20];
    ele[21][8] != ele[21][21];
    ele[21][8] != ele[21][22];
    ele[21][8] != ele[21][23];
    ele[21][8] != ele[21][24];
    ele[21][8] != ele[21][25];
    ele[21][8] != ele[21][26];
    ele[21][8] != ele[21][27];
    ele[21][8] != ele[21][28];
    ele[21][8] != ele[21][29];
    ele[21][8] != ele[21][30];
    ele[21][8] != ele[21][31];
    ele[21][8] != ele[21][32];
    ele[21][8] != ele[21][33];
    ele[21][8] != ele[21][34];
    ele[21][8] != ele[21][35];
    ele[21][8] != ele[21][9];
    ele[21][8] != ele[22][10];
    ele[21][8] != ele[22][11];
    ele[21][8] != ele[22][6];
    ele[21][8] != ele[22][7];
    ele[21][8] != ele[22][8];
    ele[21][8] != ele[22][9];
    ele[21][8] != ele[23][10];
    ele[21][8] != ele[23][11];
    ele[21][8] != ele[23][6];
    ele[21][8] != ele[23][7];
    ele[21][8] != ele[23][8];
    ele[21][8] != ele[23][9];
    ele[21][8] != ele[24][8];
    ele[21][8] != ele[25][8];
    ele[21][8] != ele[26][8];
    ele[21][8] != ele[27][8];
    ele[21][8] != ele[28][8];
    ele[21][8] != ele[29][8];
    ele[21][8] != ele[30][8];
    ele[21][8] != ele[31][8];
    ele[21][8] != ele[32][8];
    ele[21][8] != ele[33][8];
    ele[21][8] != ele[34][8];
    ele[21][8] != ele[35][8];
    ele[21][9] != ele[21][10];
    ele[21][9] != ele[21][11];
    ele[21][9] != ele[21][12];
    ele[21][9] != ele[21][13];
    ele[21][9] != ele[21][14];
    ele[21][9] != ele[21][15];
    ele[21][9] != ele[21][16];
    ele[21][9] != ele[21][17];
    ele[21][9] != ele[21][18];
    ele[21][9] != ele[21][19];
    ele[21][9] != ele[21][20];
    ele[21][9] != ele[21][21];
    ele[21][9] != ele[21][22];
    ele[21][9] != ele[21][23];
    ele[21][9] != ele[21][24];
    ele[21][9] != ele[21][25];
    ele[21][9] != ele[21][26];
    ele[21][9] != ele[21][27];
    ele[21][9] != ele[21][28];
    ele[21][9] != ele[21][29];
    ele[21][9] != ele[21][30];
    ele[21][9] != ele[21][31];
    ele[21][9] != ele[21][32];
    ele[21][9] != ele[21][33];
    ele[21][9] != ele[21][34];
    ele[21][9] != ele[21][35];
    ele[21][9] != ele[22][10];
    ele[21][9] != ele[22][11];
    ele[21][9] != ele[22][6];
    ele[21][9] != ele[22][7];
    ele[21][9] != ele[22][8];
    ele[21][9] != ele[22][9];
    ele[21][9] != ele[23][10];
    ele[21][9] != ele[23][11];
    ele[21][9] != ele[23][6];
    ele[21][9] != ele[23][7];
    ele[21][9] != ele[23][8];
    ele[21][9] != ele[23][9];
    ele[21][9] != ele[24][9];
    ele[21][9] != ele[25][9];
    ele[21][9] != ele[26][9];
    ele[21][9] != ele[27][9];
    ele[21][9] != ele[28][9];
    ele[21][9] != ele[29][9];
    ele[21][9] != ele[30][9];
    ele[21][9] != ele[31][9];
    ele[21][9] != ele[32][9];
    ele[21][9] != ele[33][9];
    ele[21][9] != ele[34][9];
    ele[21][9] != ele[35][9];
    ele[22][0] != ele[22][1];
    ele[22][0] != ele[22][10];
    ele[22][0] != ele[22][11];
    ele[22][0] != ele[22][12];
    ele[22][0] != ele[22][13];
    ele[22][0] != ele[22][14];
    ele[22][0] != ele[22][15];
    ele[22][0] != ele[22][16];
    ele[22][0] != ele[22][17];
    ele[22][0] != ele[22][18];
    ele[22][0] != ele[22][19];
    ele[22][0] != ele[22][2];
    ele[22][0] != ele[22][20];
    ele[22][0] != ele[22][21];
    ele[22][0] != ele[22][22];
    ele[22][0] != ele[22][23];
    ele[22][0] != ele[22][24];
    ele[22][0] != ele[22][25];
    ele[22][0] != ele[22][26];
    ele[22][0] != ele[22][27];
    ele[22][0] != ele[22][28];
    ele[22][0] != ele[22][29];
    ele[22][0] != ele[22][3];
    ele[22][0] != ele[22][30];
    ele[22][0] != ele[22][31];
    ele[22][0] != ele[22][32];
    ele[22][0] != ele[22][33];
    ele[22][0] != ele[22][34];
    ele[22][0] != ele[22][35];
    ele[22][0] != ele[22][4];
    ele[22][0] != ele[22][5];
    ele[22][0] != ele[22][6];
    ele[22][0] != ele[22][7];
    ele[22][0] != ele[22][8];
    ele[22][0] != ele[22][9];
    ele[22][0] != ele[23][0];
    ele[22][0] != ele[23][1];
    ele[22][0] != ele[23][2];
    ele[22][0] != ele[23][3];
    ele[22][0] != ele[23][4];
    ele[22][0] != ele[23][5];
    ele[22][0] != ele[24][0];
    ele[22][0] != ele[25][0];
    ele[22][0] != ele[26][0];
    ele[22][0] != ele[27][0];
    ele[22][0] != ele[28][0];
    ele[22][0] != ele[29][0];
    ele[22][0] != ele[30][0];
    ele[22][0] != ele[31][0];
    ele[22][0] != ele[32][0];
    ele[22][0] != ele[33][0];
    ele[22][0] != ele[34][0];
    ele[22][0] != ele[35][0];
    ele[22][1] != ele[22][10];
    ele[22][1] != ele[22][11];
    ele[22][1] != ele[22][12];
    ele[22][1] != ele[22][13];
    ele[22][1] != ele[22][14];
    ele[22][1] != ele[22][15];
    ele[22][1] != ele[22][16];
    ele[22][1] != ele[22][17];
    ele[22][1] != ele[22][18];
    ele[22][1] != ele[22][19];
    ele[22][1] != ele[22][2];
    ele[22][1] != ele[22][20];
    ele[22][1] != ele[22][21];
    ele[22][1] != ele[22][22];
    ele[22][1] != ele[22][23];
    ele[22][1] != ele[22][24];
    ele[22][1] != ele[22][25];
    ele[22][1] != ele[22][26];
    ele[22][1] != ele[22][27];
    ele[22][1] != ele[22][28];
    ele[22][1] != ele[22][29];
    ele[22][1] != ele[22][3];
    ele[22][1] != ele[22][30];
    ele[22][1] != ele[22][31];
    ele[22][1] != ele[22][32];
    ele[22][1] != ele[22][33];
    ele[22][1] != ele[22][34];
    ele[22][1] != ele[22][35];
    ele[22][1] != ele[22][4];
    ele[22][1] != ele[22][5];
    ele[22][1] != ele[22][6];
    ele[22][1] != ele[22][7];
    ele[22][1] != ele[22][8];
    ele[22][1] != ele[22][9];
    ele[22][1] != ele[23][0];
    ele[22][1] != ele[23][1];
    ele[22][1] != ele[23][2];
    ele[22][1] != ele[23][3];
    ele[22][1] != ele[23][4];
    ele[22][1] != ele[23][5];
    ele[22][1] != ele[24][1];
    ele[22][1] != ele[25][1];
    ele[22][1] != ele[26][1];
    ele[22][1] != ele[27][1];
    ele[22][1] != ele[28][1];
    ele[22][1] != ele[29][1];
    ele[22][1] != ele[30][1];
    ele[22][1] != ele[31][1];
    ele[22][1] != ele[32][1];
    ele[22][1] != ele[33][1];
    ele[22][1] != ele[34][1];
    ele[22][1] != ele[35][1];
    ele[22][10] != ele[22][11];
    ele[22][10] != ele[22][12];
    ele[22][10] != ele[22][13];
    ele[22][10] != ele[22][14];
    ele[22][10] != ele[22][15];
    ele[22][10] != ele[22][16];
    ele[22][10] != ele[22][17];
    ele[22][10] != ele[22][18];
    ele[22][10] != ele[22][19];
    ele[22][10] != ele[22][20];
    ele[22][10] != ele[22][21];
    ele[22][10] != ele[22][22];
    ele[22][10] != ele[22][23];
    ele[22][10] != ele[22][24];
    ele[22][10] != ele[22][25];
    ele[22][10] != ele[22][26];
    ele[22][10] != ele[22][27];
    ele[22][10] != ele[22][28];
    ele[22][10] != ele[22][29];
    ele[22][10] != ele[22][30];
    ele[22][10] != ele[22][31];
    ele[22][10] != ele[22][32];
    ele[22][10] != ele[22][33];
    ele[22][10] != ele[22][34];
    ele[22][10] != ele[22][35];
    ele[22][10] != ele[23][10];
    ele[22][10] != ele[23][11];
    ele[22][10] != ele[23][6];
    ele[22][10] != ele[23][7];
    ele[22][10] != ele[23][8];
    ele[22][10] != ele[23][9];
    ele[22][10] != ele[24][10];
    ele[22][10] != ele[25][10];
    ele[22][10] != ele[26][10];
    ele[22][10] != ele[27][10];
    ele[22][10] != ele[28][10];
    ele[22][10] != ele[29][10];
    ele[22][10] != ele[30][10];
    ele[22][10] != ele[31][10];
    ele[22][10] != ele[32][10];
    ele[22][10] != ele[33][10];
    ele[22][10] != ele[34][10];
    ele[22][10] != ele[35][10];
    ele[22][11] != ele[22][12];
    ele[22][11] != ele[22][13];
    ele[22][11] != ele[22][14];
    ele[22][11] != ele[22][15];
    ele[22][11] != ele[22][16];
    ele[22][11] != ele[22][17];
    ele[22][11] != ele[22][18];
    ele[22][11] != ele[22][19];
    ele[22][11] != ele[22][20];
    ele[22][11] != ele[22][21];
    ele[22][11] != ele[22][22];
    ele[22][11] != ele[22][23];
    ele[22][11] != ele[22][24];
    ele[22][11] != ele[22][25];
    ele[22][11] != ele[22][26];
    ele[22][11] != ele[22][27];
    ele[22][11] != ele[22][28];
    ele[22][11] != ele[22][29];
    ele[22][11] != ele[22][30];
    ele[22][11] != ele[22][31];
    ele[22][11] != ele[22][32];
    ele[22][11] != ele[22][33];
    ele[22][11] != ele[22][34];
    ele[22][11] != ele[22][35];
    ele[22][11] != ele[23][10];
    ele[22][11] != ele[23][11];
    ele[22][11] != ele[23][6];
    ele[22][11] != ele[23][7];
    ele[22][11] != ele[23][8];
    ele[22][11] != ele[23][9];
    ele[22][11] != ele[24][11];
    ele[22][11] != ele[25][11];
    ele[22][11] != ele[26][11];
    ele[22][11] != ele[27][11];
    ele[22][11] != ele[28][11];
    ele[22][11] != ele[29][11];
    ele[22][11] != ele[30][11];
    ele[22][11] != ele[31][11];
    ele[22][11] != ele[32][11];
    ele[22][11] != ele[33][11];
    ele[22][11] != ele[34][11];
    ele[22][11] != ele[35][11];
    ele[22][12] != ele[22][13];
    ele[22][12] != ele[22][14];
    ele[22][12] != ele[22][15];
    ele[22][12] != ele[22][16];
    ele[22][12] != ele[22][17];
    ele[22][12] != ele[22][18];
    ele[22][12] != ele[22][19];
    ele[22][12] != ele[22][20];
    ele[22][12] != ele[22][21];
    ele[22][12] != ele[22][22];
    ele[22][12] != ele[22][23];
    ele[22][12] != ele[22][24];
    ele[22][12] != ele[22][25];
    ele[22][12] != ele[22][26];
    ele[22][12] != ele[22][27];
    ele[22][12] != ele[22][28];
    ele[22][12] != ele[22][29];
    ele[22][12] != ele[22][30];
    ele[22][12] != ele[22][31];
    ele[22][12] != ele[22][32];
    ele[22][12] != ele[22][33];
    ele[22][12] != ele[22][34];
    ele[22][12] != ele[22][35];
    ele[22][12] != ele[23][12];
    ele[22][12] != ele[23][13];
    ele[22][12] != ele[23][14];
    ele[22][12] != ele[23][15];
    ele[22][12] != ele[23][16];
    ele[22][12] != ele[23][17];
    ele[22][12] != ele[24][12];
    ele[22][12] != ele[25][12];
    ele[22][12] != ele[26][12];
    ele[22][12] != ele[27][12];
    ele[22][12] != ele[28][12];
    ele[22][12] != ele[29][12];
    ele[22][12] != ele[30][12];
    ele[22][12] != ele[31][12];
    ele[22][12] != ele[32][12];
    ele[22][12] != ele[33][12];
    ele[22][12] != ele[34][12];
    ele[22][12] != ele[35][12];
    ele[22][13] != ele[22][14];
    ele[22][13] != ele[22][15];
    ele[22][13] != ele[22][16];
    ele[22][13] != ele[22][17];
    ele[22][13] != ele[22][18];
    ele[22][13] != ele[22][19];
    ele[22][13] != ele[22][20];
    ele[22][13] != ele[22][21];
    ele[22][13] != ele[22][22];
    ele[22][13] != ele[22][23];
    ele[22][13] != ele[22][24];
    ele[22][13] != ele[22][25];
    ele[22][13] != ele[22][26];
    ele[22][13] != ele[22][27];
    ele[22][13] != ele[22][28];
    ele[22][13] != ele[22][29];
    ele[22][13] != ele[22][30];
    ele[22][13] != ele[22][31];
    ele[22][13] != ele[22][32];
    ele[22][13] != ele[22][33];
    ele[22][13] != ele[22][34];
    ele[22][13] != ele[22][35];
    ele[22][13] != ele[23][12];
    ele[22][13] != ele[23][13];
    ele[22][13] != ele[23][14];
    ele[22][13] != ele[23][15];
    ele[22][13] != ele[23][16];
    ele[22][13] != ele[23][17];
    ele[22][13] != ele[24][13];
    ele[22][13] != ele[25][13];
    ele[22][13] != ele[26][13];
    ele[22][13] != ele[27][13];
    ele[22][13] != ele[28][13];
    ele[22][13] != ele[29][13];
    ele[22][13] != ele[30][13];
    ele[22][13] != ele[31][13];
    ele[22][13] != ele[32][13];
    ele[22][13] != ele[33][13];
    ele[22][13] != ele[34][13];
    ele[22][13] != ele[35][13];
    ele[22][14] != ele[22][15];
    ele[22][14] != ele[22][16];
    ele[22][14] != ele[22][17];
    ele[22][14] != ele[22][18];
    ele[22][14] != ele[22][19];
    ele[22][14] != ele[22][20];
    ele[22][14] != ele[22][21];
    ele[22][14] != ele[22][22];
    ele[22][14] != ele[22][23];
    ele[22][14] != ele[22][24];
    ele[22][14] != ele[22][25];
    ele[22][14] != ele[22][26];
    ele[22][14] != ele[22][27];
    ele[22][14] != ele[22][28];
    ele[22][14] != ele[22][29];
    ele[22][14] != ele[22][30];
    ele[22][14] != ele[22][31];
    ele[22][14] != ele[22][32];
    ele[22][14] != ele[22][33];
    ele[22][14] != ele[22][34];
    ele[22][14] != ele[22][35];
    ele[22][14] != ele[23][12];
    ele[22][14] != ele[23][13];
    ele[22][14] != ele[23][14];
    ele[22][14] != ele[23][15];
    ele[22][14] != ele[23][16];
    ele[22][14] != ele[23][17];
    ele[22][14] != ele[24][14];
    ele[22][14] != ele[25][14];
    ele[22][14] != ele[26][14];
    ele[22][14] != ele[27][14];
    ele[22][14] != ele[28][14];
    ele[22][14] != ele[29][14];
    ele[22][14] != ele[30][14];
    ele[22][14] != ele[31][14];
    ele[22][14] != ele[32][14];
    ele[22][14] != ele[33][14];
    ele[22][14] != ele[34][14];
    ele[22][14] != ele[35][14];
    ele[22][15] != ele[22][16];
    ele[22][15] != ele[22][17];
    ele[22][15] != ele[22][18];
    ele[22][15] != ele[22][19];
    ele[22][15] != ele[22][20];
    ele[22][15] != ele[22][21];
    ele[22][15] != ele[22][22];
    ele[22][15] != ele[22][23];
    ele[22][15] != ele[22][24];
    ele[22][15] != ele[22][25];
    ele[22][15] != ele[22][26];
    ele[22][15] != ele[22][27];
    ele[22][15] != ele[22][28];
    ele[22][15] != ele[22][29];
    ele[22][15] != ele[22][30];
    ele[22][15] != ele[22][31];
    ele[22][15] != ele[22][32];
    ele[22][15] != ele[22][33];
    ele[22][15] != ele[22][34];
    ele[22][15] != ele[22][35];
    ele[22][15] != ele[23][12];
    ele[22][15] != ele[23][13];
    ele[22][15] != ele[23][14];
    ele[22][15] != ele[23][15];
    ele[22][15] != ele[23][16];
    ele[22][15] != ele[23][17];
    ele[22][15] != ele[24][15];
    ele[22][15] != ele[25][15];
    ele[22][15] != ele[26][15];
    ele[22][15] != ele[27][15];
    ele[22][15] != ele[28][15];
    ele[22][15] != ele[29][15];
    ele[22][15] != ele[30][15];
    ele[22][15] != ele[31][15];
    ele[22][15] != ele[32][15];
    ele[22][15] != ele[33][15];
    ele[22][15] != ele[34][15];
    ele[22][15] != ele[35][15];
    ele[22][16] != ele[22][17];
    ele[22][16] != ele[22][18];
    ele[22][16] != ele[22][19];
    ele[22][16] != ele[22][20];
    ele[22][16] != ele[22][21];
    ele[22][16] != ele[22][22];
    ele[22][16] != ele[22][23];
    ele[22][16] != ele[22][24];
    ele[22][16] != ele[22][25];
    ele[22][16] != ele[22][26];
    ele[22][16] != ele[22][27];
    ele[22][16] != ele[22][28];
    ele[22][16] != ele[22][29];
    ele[22][16] != ele[22][30];
    ele[22][16] != ele[22][31];
    ele[22][16] != ele[22][32];
    ele[22][16] != ele[22][33];
    ele[22][16] != ele[22][34];
    ele[22][16] != ele[22][35];
    ele[22][16] != ele[23][12];
    ele[22][16] != ele[23][13];
    ele[22][16] != ele[23][14];
    ele[22][16] != ele[23][15];
    ele[22][16] != ele[23][16];
    ele[22][16] != ele[23][17];
    ele[22][16] != ele[24][16];
    ele[22][16] != ele[25][16];
    ele[22][16] != ele[26][16];
    ele[22][16] != ele[27][16];
    ele[22][16] != ele[28][16];
    ele[22][16] != ele[29][16];
    ele[22][16] != ele[30][16];
    ele[22][16] != ele[31][16];
    ele[22][16] != ele[32][16];
    ele[22][16] != ele[33][16];
    ele[22][16] != ele[34][16];
    ele[22][16] != ele[35][16];
    ele[22][17] != ele[22][18];
    ele[22][17] != ele[22][19];
    ele[22][17] != ele[22][20];
    ele[22][17] != ele[22][21];
    ele[22][17] != ele[22][22];
    ele[22][17] != ele[22][23];
    ele[22][17] != ele[22][24];
    ele[22][17] != ele[22][25];
    ele[22][17] != ele[22][26];
    ele[22][17] != ele[22][27];
    ele[22][17] != ele[22][28];
    ele[22][17] != ele[22][29];
    ele[22][17] != ele[22][30];
    ele[22][17] != ele[22][31];
    ele[22][17] != ele[22][32];
    ele[22][17] != ele[22][33];
    ele[22][17] != ele[22][34];
    ele[22][17] != ele[22][35];
    ele[22][17] != ele[23][12];
    ele[22][17] != ele[23][13];
    ele[22][17] != ele[23][14];
    ele[22][17] != ele[23][15];
    ele[22][17] != ele[23][16];
    ele[22][17] != ele[23][17];
    ele[22][17] != ele[24][17];
    ele[22][17] != ele[25][17];
    ele[22][17] != ele[26][17];
    ele[22][17] != ele[27][17];
    ele[22][17] != ele[28][17];
    ele[22][17] != ele[29][17];
    ele[22][17] != ele[30][17];
    ele[22][17] != ele[31][17];
    ele[22][17] != ele[32][17];
    ele[22][17] != ele[33][17];
    ele[22][17] != ele[34][17];
    ele[22][17] != ele[35][17];
    ele[22][18] != ele[22][19];
    ele[22][18] != ele[22][20];
    ele[22][18] != ele[22][21];
    ele[22][18] != ele[22][22];
    ele[22][18] != ele[22][23];
    ele[22][18] != ele[22][24];
    ele[22][18] != ele[22][25];
    ele[22][18] != ele[22][26];
    ele[22][18] != ele[22][27];
    ele[22][18] != ele[22][28];
    ele[22][18] != ele[22][29];
    ele[22][18] != ele[22][30];
    ele[22][18] != ele[22][31];
    ele[22][18] != ele[22][32];
    ele[22][18] != ele[22][33];
    ele[22][18] != ele[22][34];
    ele[22][18] != ele[22][35];
    ele[22][18] != ele[23][18];
    ele[22][18] != ele[23][19];
    ele[22][18] != ele[23][20];
    ele[22][18] != ele[23][21];
    ele[22][18] != ele[23][22];
    ele[22][18] != ele[23][23];
    ele[22][18] != ele[24][18];
    ele[22][18] != ele[25][18];
    ele[22][18] != ele[26][18];
    ele[22][18] != ele[27][18];
    ele[22][18] != ele[28][18];
    ele[22][18] != ele[29][18];
    ele[22][18] != ele[30][18];
    ele[22][18] != ele[31][18];
    ele[22][18] != ele[32][18];
    ele[22][18] != ele[33][18];
    ele[22][18] != ele[34][18];
    ele[22][18] != ele[35][18];
    ele[22][19] != ele[22][20];
    ele[22][19] != ele[22][21];
    ele[22][19] != ele[22][22];
    ele[22][19] != ele[22][23];
    ele[22][19] != ele[22][24];
    ele[22][19] != ele[22][25];
    ele[22][19] != ele[22][26];
    ele[22][19] != ele[22][27];
    ele[22][19] != ele[22][28];
    ele[22][19] != ele[22][29];
    ele[22][19] != ele[22][30];
    ele[22][19] != ele[22][31];
    ele[22][19] != ele[22][32];
    ele[22][19] != ele[22][33];
    ele[22][19] != ele[22][34];
    ele[22][19] != ele[22][35];
    ele[22][19] != ele[23][18];
    ele[22][19] != ele[23][19];
    ele[22][19] != ele[23][20];
    ele[22][19] != ele[23][21];
    ele[22][19] != ele[23][22];
    ele[22][19] != ele[23][23];
    ele[22][19] != ele[24][19];
    ele[22][19] != ele[25][19];
    ele[22][19] != ele[26][19];
    ele[22][19] != ele[27][19];
    ele[22][19] != ele[28][19];
    ele[22][19] != ele[29][19];
    ele[22][19] != ele[30][19];
    ele[22][19] != ele[31][19];
    ele[22][19] != ele[32][19];
    ele[22][19] != ele[33][19];
    ele[22][19] != ele[34][19];
    ele[22][19] != ele[35][19];
    ele[22][2] != ele[22][10];
    ele[22][2] != ele[22][11];
    ele[22][2] != ele[22][12];
    ele[22][2] != ele[22][13];
    ele[22][2] != ele[22][14];
    ele[22][2] != ele[22][15];
    ele[22][2] != ele[22][16];
    ele[22][2] != ele[22][17];
    ele[22][2] != ele[22][18];
    ele[22][2] != ele[22][19];
    ele[22][2] != ele[22][20];
    ele[22][2] != ele[22][21];
    ele[22][2] != ele[22][22];
    ele[22][2] != ele[22][23];
    ele[22][2] != ele[22][24];
    ele[22][2] != ele[22][25];
    ele[22][2] != ele[22][26];
    ele[22][2] != ele[22][27];
    ele[22][2] != ele[22][28];
    ele[22][2] != ele[22][29];
    ele[22][2] != ele[22][3];
    ele[22][2] != ele[22][30];
    ele[22][2] != ele[22][31];
    ele[22][2] != ele[22][32];
    ele[22][2] != ele[22][33];
    ele[22][2] != ele[22][34];
    ele[22][2] != ele[22][35];
    ele[22][2] != ele[22][4];
    ele[22][2] != ele[22][5];
    ele[22][2] != ele[22][6];
    ele[22][2] != ele[22][7];
    ele[22][2] != ele[22][8];
    ele[22][2] != ele[22][9];
    ele[22][2] != ele[23][0];
    ele[22][2] != ele[23][1];
    ele[22][2] != ele[23][2];
    ele[22][2] != ele[23][3];
    ele[22][2] != ele[23][4];
    ele[22][2] != ele[23][5];
    ele[22][2] != ele[24][2];
    ele[22][2] != ele[25][2];
    ele[22][2] != ele[26][2];
    ele[22][2] != ele[27][2];
    ele[22][2] != ele[28][2];
    ele[22][2] != ele[29][2];
    ele[22][2] != ele[30][2];
    ele[22][2] != ele[31][2];
    ele[22][2] != ele[32][2];
    ele[22][2] != ele[33][2];
    ele[22][2] != ele[34][2];
    ele[22][2] != ele[35][2];
    ele[22][20] != ele[22][21];
    ele[22][20] != ele[22][22];
    ele[22][20] != ele[22][23];
    ele[22][20] != ele[22][24];
    ele[22][20] != ele[22][25];
    ele[22][20] != ele[22][26];
    ele[22][20] != ele[22][27];
    ele[22][20] != ele[22][28];
    ele[22][20] != ele[22][29];
    ele[22][20] != ele[22][30];
    ele[22][20] != ele[22][31];
    ele[22][20] != ele[22][32];
    ele[22][20] != ele[22][33];
    ele[22][20] != ele[22][34];
    ele[22][20] != ele[22][35];
    ele[22][20] != ele[23][18];
    ele[22][20] != ele[23][19];
    ele[22][20] != ele[23][20];
    ele[22][20] != ele[23][21];
    ele[22][20] != ele[23][22];
    ele[22][20] != ele[23][23];
    ele[22][20] != ele[24][20];
    ele[22][20] != ele[25][20];
    ele[22][20] != ele[26][20];
    ele[22][20] != ele[27][20];
    ele[22][20] != ele[28][20];
    ele[22][20] != ele[29][20];
    ele[22][20] != ele[30][20];
    ele[22][20] != ele[31][20];
    ele[22][20] != ele[32][20];
    ele[22][20] != ele[33][20];
    ele[22][20] != ele[34][20];
    ele[22][20] != ele[35][20];
    ele[22][21] != ele[22][22];
    ele[22][21] != ele[22][23];
    ele[22][21] != ele[22][24];
    ele[22][21] != ele[22][25];
    ele[22][21] != ele[22][26];
    ele[22][21] != ele[22][27];
    ele[22][21] != ele[22][28];
    ele[22][21] != ele[22][29];
    ele[22][21] != ele[22][30];
    ele[22][21] != ele[22][31];
    ele[22][21] != ele[22][32];
    ele[22][21] != ele[22][33];
    ele[22][21] != ele[22][34];
    ele[22][21] != ele[22][35];
    ele[22][21] != ele[23][18];
    ele[22][21] != ele[23][19];
    ele[22][21] != ele[23][20];
    ele[22][21] != ele[23][21];
    ele[22][21] != ele[23][22];
    ele[22][21] != ele[23][23];
    ele[22][21] != ele[24][21];
    ele[22][21] != ele[25][21];
    ele[22][21] != ele[26][21];
    ele[22][21] != ele[27][21];
    ele[22][21] != ele[28][21];
    ele[22][21] != ele[29][21];
    ele[22][21] != ele[30][21];
    ele[22][21] != ele[31][21];
    ele[22][21] != ele[32][21];
    ele[22][21] != ele[33][21];
    ele[22][21] != ele[34][21];
    ele[22][21] != ele[35][21];
    ele[22][22] != ele[22][23];
    ele[22][22] != ele[22][24];
    ele[22][22] != ele[22][25];
    ele[22][22] != ele[22][26];
    ele[22][22] != ele[22][27];
    ele[22][22] != ele[22][28];
    ele[22][22] != ele[22][29];
    ele[22][22] != ele[22][30];
    ele[22][22] != ele[22][31];
    ele[22][22] != ele[22][32];
    ele[22][22] != ele[22][33];
    ele[22][22] != ele[22][34];
    ele[22][22] != ele[22][35];
    ele[22][22] != ele[23][18];
    ele[22][22] != ele[23][19];
    ele[22][22] != ele[23][20];
    ele[22][22] != ele[23][21];
    ele[22][22] != ele[23][22];
    ele[22][22] != ele[23][23];
    ele[22][22] != ele[24][22];
    ele[22][22] != ele[25][22];
    ele[22][22] != ele[26][22];
    ele[22][22] != ele[27][22];
    ele[22][22] != ele[28][22];
    ele[22][22] != ele[29][22];
    ele[22][22] != ele[30][22];
    ele[22][22] != ele[31][22];
    ele[22][22] != ele[32][22];
    ele[22][22] != ele[33][22];
    ele[22][22] != ele[34][22];
    ele[22][22] != ele[35][22];
    ele[22][23] != ele[22][24];
    ele[22][23] != ele[22][25];
    ele[22][23] != ele[22][26];
    ele[22][23] != ele[22][27];
    ele[22][23] != ele[22][28];
    ele[22][23] != ele[22][29];
    ele[22][23] != ele[22][30];
    ele[22][23] != ele[22][31];
    ele[22][23] != ele[22][32];
    ele[22][23] != ele[22][33];
    ele[22][23] != ele[22][34];
    ele[22][23] != ele[22][35];
    ele[22][23] != ele[23][18];
    ele[22][23] != ele[23][19];
    ele[22][23] != ele[23][20];
    ele[22][23] != ele[23][21];
    ele[22][23] != ele[23][22];
    ele[22][23] != ele[23][23];
    ele[22][23] != ele[24][23];
    ele[22][23] != ele[25][23];
    ele[22][23] != ele[26][23];
    ele[22][23] != ele[27][23];
    ele[22][23] != ele[28][23];
    ele[22][23] != ele[29][23];
    ele[22][23] != ele[30][23];
    ele[22][23] != ele[31][23];
    ele[22][23] != ele[32][23];
    ele[22][23] != ele[33][23];
    ele[22][23] != ele[34][23];
    ele[22][23] != ele[35][23];
    ele[22][24] != ele[22][25];
    ele[22][24] != ele[22][26];
    ele[22][24] != ele[22][27];
    ele[22][24] != ele[22][28];
    ele[22][24] != ele[22][29];
    ele[22][24] != ele[22][30];
    ele[22][24] != ele[22][31];
    ele[22][24] != ele[22][32];
    ele[22][24] != ele[22][33];
    ele[22][24] != ele[22][34];
    ele[22][24] != ele[22][35];
    ele[22][24] != ele[23][24];
    ele[22][24] != ele[23][25];
    ele[22][24] != ele[23][26];
    ele[22][24] != ele[23][27];
    ele[22][24] != ele[23][28];
    ele[22][24] != ele[23][29];
    ele[22][24] != ele[24][24];
    ele[22][24] != ele[25][24];
    ele[22][24] != ele[26][24];
    ele[22][24] != ele[27][24];
    ele[22][24] != ele[28][24];
    ele[22][24] != ele[29][24];
    ele[22][24] != ele[30][24];
    ele[22][24] != ele[31][24];
    ele[22][24] != ele[32][24];
    ele[22][24] != ele[33][24];
    ele[22][24] != ele[34][24];
    ele[22][24] != ele[35][24];
    ele[22][25] != ele[22][26];
    ele[22][25] != ele[22][27];
    ele[22][25] != ele[22][28];
    ele[22][25] != ele[22][29];
    ele[22][25] != ele[22][30];
    ele[22][25] != ele[22][31];
    ele[22][25] != ele[22][32];
    ele[22][25] != ele[22][33];
    ele[22][25] != ele[22][34];
    ele[22][25] != ele[22][35];
    ele[22][25] != ele[23][24];
    ele[22][25] != ele[23][25];
    ele[22][25] != ele[23][26];
    ele[22][25] != ele[23][27];
    ele[22][25] != ele[23][28];
    ele[22][25] != ele[23][29];
    ele[22][25] != ele[24][25];
    ele[22][25] != ele[25][25];
    ele[22][25] != ele[26][25];
    ele[22][25] != ele[27][25];
    ele[22][25] != ele[28][25];
    ele[22][25] != ele[29][25];
    ele[22][25] != ele[30][25];
    ele[22][25] != ele[31][25];
    ele[22][25] != ele[32][25];
    ele[22][25] != ele[33][25];
    ele[22][25] != ele[34][25];
    ele[22][25] != ele[35][25];
    ele[22][26] != ele[22][27];
    ele[22][26] != ele[22][28];
    ele[22][26] != ele[22][29];
    ele[22][26] != ele[22][30];
    ele[22][26] != ele[22][31];
    ele[22][26] != ele[22][32];
    ele[22][26] != ele[22][33];
    ele[22][26] != ele[22][34];
    ele[22][26] != ele[22][35];
    ele[22][26] != ele[23][24];
    ele[22][26] != ele[23][25];
    ele[22][26] != ele[23][26];
    ele[22][26] != ele[23][27];
    ele[22][26] != ele[23][28];
    ele[22][26] != ele[23][29];
    ele[22][26] != ele[24][26];
    ele[22][26] != ele[25][26];
    ele[22][26] != ele[26][26];
    ele[22][26] != ele[27][26];
    ele[22][26] != ele[28][26];
    ele[22][26] != ele[29][26];
    ele[22][26] != ele[30][26];
    ele[22][26] != ele[31][26];
    ele[22][26] != ele[32][26];
    ele[22][26] != ele[33][26];
    ele[22][26] != ele[34][26];
    ele[22][26] != ele[35][26];
    ele[22][27] != ele[22][28];
    ele[22][27] != ele[22][29];
    ele[22][27] != ele[22][30];
    ele[22][27] != ele[22][31];
    ele[22][27] != ele[22][32];
    ele[22][27] != ele[22][33];
    ele[22][27] != ele[22][34];
    ele[22][27] != ele[22][35];
    ele[22][27] != ele[23][24];
    ele[22][27] != ele[23][25];
    ele[22][27] != ele[23][26];
    ele[22][27] != ele[23][27];
    ele[22][27] != ele[23][28];
    ele[22][27] != ele[23][29];
    ele[22][27] != ele[24][27];
    ele[22][27] != ele[25][27];
    ele[22][27] != ele[26][27];
    ele[22][27] != ele[27][27];
    ele[22][27] != ele[28][27];
    ele[22][27] != ele[29][27];
    ele[22][27] != ele[30][27];
    ele[22][27] != ele[31][27];
    ele[22][27] != ele[32][27];
    ele[22][27] != ele[33][27];
    ele[22][27] != ele[34][27];
    ele[22][27] != ele[35][27];
    ele[22][28] != ele[22][29];
    ele[22][28] != ele[22][30];
    ele[22][28] != ele[22][31];
    ele[22][28] != ele[22][32];
    ele[22][28] != ele[22][33];
    ele[22][28] != ele[22][34];
    ele[22][28] != ele[22][35];
    ele[22][28] != ele[23][24];
    ele[22][28] != ele[23][25];
    ele[22][28] != ele[23][26];
    ele[22][28] != ele[23][27];
    ele[22][28] != ele[23][28];
    ele[22][28] != ele[23][29];
    ele[22][28] != ele[24][28];
    ele[22][28] != ele[25][28];
    ele[22][28] != ele[26][28];
    ele[22][28] != ele[27][28];
    ele[22][28] != ele[28][28];
    ele[22][28] != ele[29][28];
    ele[22][28] != ele[30][28];
    ele[22][28] != ele[31][28];
    ele[22][28] != ele[32][28];
    ele[22][28] != ele[33][28];
    ele[22][28] != ele[34][28];
    ele[22][28] != ele[35][28];
    ele[22][29] != ele[22][30];
    ele[22][29] != ele[22][31];
    ele[22][29] != ele[22][32];
    ele[22][29] != ele[22][33];
    ele[22][29] != ele[22][34];
    ele[22][29] != ele[22][35];
    ele[22][29] != ele[23][24];
    ele[22][29] != ele[23][25];
    ele[22][29] != ele[23][26];
    ele[22][29] != ele[23][27];
    ele[22][29] != ele[23][28];
    ele[22][29] != ele[23][29];
    ele[22][29] != ele[24][29];
    ele[22][29] != ele[25][29];
    ele[22][29] != ele[26][29];
    ele[22][29] != ele[27][29];
    ele[22][29] != ele[28][29];
    ele[22][29] != ele[29][29];
    ele[22][29] != ele[30][29];
    ele[22][29] != ele[31][29];
    ele[22][29] != ele[32][29];
    ele[22][29] != ele[33][29];
    ele[22][29] != ele[34][29];
    ele[22][29] != ele[35][29];
    ele[22][3] != ele[22][10];
    ele[22][3] != ele[22][11];
    ele[22][3] != ele[22][12];
    ele[22][3] != ele[22][13];
    ele[22][3] != ele[22][14];
    ele[22][3] != ele[22][15];
    ele[22][3] != ele[22][16];
    ele[22][3] != ele[22][17];
    ele[22][3] != ele[22][18];
    ele[22][3] != ele[22][19];
    ele[22][3] != ele[22][20];
    ele[22][3] != ele[22][21];
    ele[22][3] != ele[22][22];
    ele[22][3] != ele[22][23];
    ele[22][3] != ele[22][24];
    ele[22][3] != ele[22][25];
    ele[22][3] != ele[22][26];
    ele[22][3] != ele[22][27];
    ele[22][3] != ele[22][28];
    ele[22][3] != ele[22][29];
    ele[22][3] != ele[22][30];
    ele[22][3] != ele[22][31];
    ele[22][3] != ele[22][32];
    ele[22][3] != ele[22][33];
    ele[22][3] != ele[22][34];
    ele[22][3] != ele[22][35];
    ele[22][3] != ele[22][4];
    ele[22][3] != ele[22][5];
    ele[22][3] != ele[22][6];
    ele[22][3] != ele[22][7];
    ele[22][3] != ele[22][8];
    ele[22][3] != ele[22][9];
    ele[22][3] != ele[23][0];
    ele[22][3] != ele[23][1];
    ele[22][3] != ele[23][2];
    ele[22][3] != ele[23][3];
    ele[22][3] != ele[23][4];
    ele[22][3] != ele[23][5];
    ele[22][3] != ele[24][3];
    ele[22][3] != ele[25][3];
    ele[22][3] != ele[26][3];
    ele[22][3] != ele[27][3];
    ele[22][3] != ele[28][3];
    ele[22][3] != ele[29][3];
    ele[22][3] != ele[30][3];
    ele[22][3] != ele[31][3];
    ele[22][3] != ele[32][3];
    ele[22][3] != ele[33][3];
    ele[22][3] != ele[34][3];
    ele[22][3] != ele[35][3];
    ele[22][30] != ele[22][31];
    ele[22][30] != ele[22][32];
    ele[22][30] != ele[22][33];
    ele[22][30] != ele[22][34];
    ele[22][30] != ele[22][35];
    ele[22][30] != ele[23][30];
    ele[22][30] != ele[23][31];
    ele[22][30] != ele[23][32];
    ele[22][30] != ele[23][33];
    ele[22][30] != ele[23][34];
    ele[22][30] != ele[23][35];
    ele[22][30] != ele[24][30];
    ele[22][30] != ele[25][30];
    ele[22][30] != ele[26][30];
    ele[22][30] != ele[27][30];
    ele[22][30] != ele[28][30];
    ele[22][30] != ele[29][30];
    ele[22][30] != ele[30][30];
    ele[22][30] != ele[31][30];
    ele[22][30] != ele[32][30];
    ele[22][30] != ele[33][30];
    ele[22][30] != ele[34][30];
    ele[22][30] != ele[35][30];
    ele[22][31] != ele[22][32];
    ele[22][31] != ele[22][33];
    ele[22][31] != ele[22][34];
    ele[22][31] != ele[22][35];
    ele[22][31] != ele[23][30];
    ele[22][31] != ele[23][31];
    ele[22][31] != ele[23][32];
    ele[22][31] != ele[23][33];
    ele[22][31] != ele[23][34];
    ele[22][31] != ele[23][35];
    ele[22][31] != ele[24][31];
    ele[22][31] != ele[25][31];
    ele[22][31] != ele[26][31];
    ele[22][31] != ele[27][31];
    ele[22][31] != ele[28][31];
    ele[22][31] != ele[29][31];
    ele[22][31] != ele[30][31];
    ele[22][31] != ele[31][31];
    ele[22][31] != ele[32][31];
    ele[22][31] != ele[33][31];
    ele[22][31] != ele[34][31];
    ele[22][31] != ele[35][31];
    ele[22][32] != ele[22][33];
    ele[22][32] != ele[22][34];
    ele[22][32] != ele[22][35];
    ele[22][32] != ele[23][30];
    ele[22][32] != ele[23][31];
    ele[22][32] != ele[23][32];
    ele[22][32] != ele[23][33];
    ele[22][32] != ele[23][34];
    ele[22][32] != ele[23][35];
    ele[22][32] != ele[24][32];
    ele[22][32] != ele[25][32];
    ele[22][32] != ele[26][32];
    ele[22][32] != ele[27][32];
    ele[22][32] != ele[28][32];
    ele[22][32] != ele[29][32];
    ele[22][32] != ele[30][32];
    ele[22][32] != ele[31][32];
    ele[22][32] != ele[32][32];
    ele[22][32] != ele[33][32];
    ele[22][32] != ele[34][32];
    ele[22][32] != ele[35][32];
    ele[22][33] != ele[22][34];
    ele[22][33] != ele[22][35];
    ele[22][33] != ele[23][30];
    ele[22][33] != ele[23][31];
    ele[22][33] != ele[23][32];
    ele[22][33] != ele[23][33];
    ele[22][33] != ele[23][34];
    ele[22][33] != ele[23][35];
    ele[22][33] != ele[24][33];
    ele[22][33] != ele[25][33];
    ele[22][33] != ele[26][33];
    ele[22][33] != ele[27][33];
    ele[22][33] != ele[28][33];
    ele[22][33] != ele[29][33];
    ele[22][33] != ele[30][33];
    ele[22][33] != ele[31][33];
    ele[22][33] != ele[32][33];
    ele[22][33] != ele[33][33];
    ele[22][33] != ele[34][33];
    ele[22][33] != ele[35][33];
    ele[22][34] != ele[22][35];
    ele[22][34] != ele[23][30];
    ele[22][34] != ele[23][31];
    ele[22][34] != ele[23][32];
    ele[22][34] != ele[23][33];
    ele[22][34] != ele[23][34];
    ele[22][34] != ele[23][35];
    ele[22][34] != ele[24][34];
    ele[22][34] != ele[25][34];
    ele[22][34] != ele[26][34];
    ele[22][34] != ele[27][34];
    ele[22][34] != ele[28][34];
    ele[22][34] != ele[29][34];
    ele[22][34] != ele[30][34];
    ele[22][34] != ele[31][34];
    ele[22][34] != ele[32][34];
    ele[22][34] != ele[33][34];
    ele[22][34] != ele[34][34];
    ele[22][34] != ele[35][34];
    ele[22][35] != ele[23][30];
    ele[22][35] != ele[23][31];
    ele[22][35] != ele[23][32];
    ele[22][35] != ele[23][33];
    ele[22][35] != ele[23][34];
    ele[22][35] != ele[23][35];
    ele[22][35] != ele[24][35];
    ele[22][35] != ele[25][35];
    ele[22][35] != ele[26][35];
    ele[22][35] != ele[27][35];
    ele[22][35] != ele[28][35];
    ele[22][35] != ele[29][35];
    ele[22][35] != ele[30][35];
    ele[22][35] != ele[31][35];
    ele[22][35] != ele[32][35];
    ele[22][35] != ele[33][35];
    ele[22][35] != ele[34][35];
    ele[22][35] != ele[35][35];
    ele[22][4] != ele[22][10];
    ele[22][4] != ele[22][11];
    ele[22][4] != ele[22][12];
    ele[22][4] != ele[22][13];
    ele[22][4] != ele[22][14];
    ele[22][4] != ele[22][15];
    ele[22][4] != ele[22][16];
    ele[22][4] != ele[22][17];
    ele[22][4] != ele[22][18];
    ele[22][4] != ele[22][19];
    ele[22][4] != ele[22][20];
    ele[22][4] != ele[22][21];
    ele[22][4] != ele[22][22];
    ele[22][4] != ele[22][23];
    ele[22][4] != ele[22][24];
    ele[22][4] != ele[22][25];
    ele[22][4] != ele[22][26];
    ele[22][4] != ele[22][27];
    ele[22][4] != ele[22][28];
    ele[22][4] != ele[22][29];
    ele[22][4] != ele[22][30];
    ele[22][4] != ele[22][31];
    ele[22][4] != ele[22][32];
    ele[22][4] != ele[22][33];
    ele[22][4] != ele[22][34];
    ele[22][4] != ele[22][35];
    ele[22][4] != ele[22][5];
    ele[22][4] != ele[22][6];
    ele[22][4] != ele[22][7];
    ele[22][4] != ele[22][8];
    ele[22][4] != ele[22][9];
    ele[22][4] != ele[23][0];
    ele[22][4] != ele[23][1];
    ele[22][4] != ele[23][2];
    ele[22][4] != ele[23][3];
    ele[22][4] != ele[23][4];
    ele[22][4] != ele[23][5];
    ele[22][4] != ele[24][4];
    ele[22][4] != ele[25][4];
    ele[22][4] != ele[26][4];
    ele[22][4] != ele[27][4];
    ele[22][4] != ele[28][4];
    ele[22][4] != ele[29][4];
    ele[22][4] != ele[30][4];
    ele[22][4] != ele[31][4];
    ele[22][4] != ele[32][4];
    ele[22][4] != ele[33][4];
    ele[22][4] != ele[34][4];
    ele[22][4] != ele[35][4];
    ele[22][5] != ele[22][10];
    ele[22][5] != ele[22][11];
    ele[22][5] != ele[22][12];
    ele[22][5] != ele[22][13];
    ele[22][5] != ele[22][14];
    ele[22][5] != ele[22][15];
    ele[22][5] != ele[22][16];
    ele[22][5] != ele[22][17];
    ele[22][5] != ele[22][18];
    ele[22][5] != ele[22][19];
    ele[22][5] != ele[22][20];
    ele[22][5] != ele[22][21];
    ele[22][5] != ele[22][22];
    ele[22][5] != ele[22][23];
    ele[22][5] != ele[22][24];
    ele[22][5] != ele[22][25];
    ele[22][5] != ele[22][26];
    ele[22][5] != ele[22][27];
    ele[22][5] != ele[22][28];
    ele[22][5] != ele[22][29];
    ele[22][5] != ele[22][30];
    ele[22][5] != ele[22][31];
    ele[22][5] != ele[22][32];
    ele[22][5] != ele[22][33];
    ele[22][5] != ele[22][34];
    ele[22][5] != ele[22][35];
    ele[22][5] != ele[22][6];
    ele[22][5] != ele[22][7];
    ele[22][5] != ele[22][8];
    ele[22][5] != ele[22][9];
    ele[22][5] != ele[23][0];
    ele[22][5] != ele[23][1];
    ele[22][5] != ele[23][2];
    ele[22][5] != ele[23][3];
    ele[22][5] != ele[23][4];
    ele[22][5] != ele[23][5];
    ele[22][5] != ele[24][5];
    ele[22][5] != ele[25][5];
    ele[22][5] != ele[26][5];
    ele[22][5] != ele[27][5];
    ele[22][5] != ele[28][5];
    ele[22][5] != ele[29][5];
    ele[22][5] != ele[30][5];
    ele[22][5] != ele[31][5];
    ele[22][5] != ele[32][5];
    ele[22][5] != ele[33][5];
    ele[22][5] != ele[34][5];
    ele[22][5] != ele[35][5];
    ele[22][6] != ele[22][10];
    ele[22][6] != ele[22][11];
    ele[22][6] != ele[22][12];
    ele[22][6] != ele[22][13];
    ele[22][6] != ele[22][14];
    ele[22][6] != ele[22][15];
    ele[22][6] != ele[22][16];
    ele[22][6] != ele[22][17];
    ele[22][6] != ele[22][18];
    ele[22][6] != ele[22][19];
    ele[22][6] != ele[22][20];
    ele[22][6] != ele[22][21];
    ele[22][6] != ele[22][22];
    ele[22][6] != ele[22][23];
    ele[22][6] != ele[22][24];
    ele[22][6] != ele[22][25];
    ele[22][6] != ele[22][26];
    ele[22][6] != ele[22][27];
    ele[22][6] != ele[22][28];
    ele[22][6] != ele[22][29];
    ele[22][6] != ele[22][30];
    ele[22][6] != ele[22][31];
    ele[22][6] != ele[22][32];
    ele[22][6] != ele[22][33];
    ele[22][6] != ele[22][34];
    ele[22][6] != ele[22][35];
    ele[22][6] != ele[22][7];
    ele[22][6] != ele[22][8];
    ele[22][6] != ele[22][9];
    ele[22][6] != ele[23][10];
    ele[22][6] != ele[23][11];
    ele[22][6] != ele[23][6];
    ele[22][6] != ele[23][7];
    ele[22][6] != ele[23][8];
    ele[22][6] != ele[23][9];
    ele[22][6] != ele[24][6];
    ele[22][6] != ele[25][6];
    ele[22][6] != ele[26][6];
    ele[22][6] != ele[27][6];
    ele[22][6] != ele[28][6];
    ele[22][6] != ele[29][6];
    ele[22][6] != ele[30][6];
    ele[22][6] != ele[31][6];
    ele[22][6] != ele[32][6];
    ele[22][6] != ele[33][6];
    ele[22][6] != ele[34][6];
    ele[22][6] != ele[35][6];
    ele[22][7] != ele[22][10];
    ele[22][7] != ele[22][11];
    ele[22][7] != ele[22][12];
    ele[22][7] != ele[22][13];
    ele[22][7] != ele[22][14];
    ele[22][7] != ele[22][15];
    ele[22][7] != ele[22][16];
    ele[22][7] != ele[22][17];
    ele[22][7] != ele[22][18];
    ele[22][7] != ele[22][19];
    ele[22][7] != ele[22][20];
    ele[22][7] != ele[22][21];
    ele[22][7] != ele[22][22];
    ele[22][7] != ele[22][23];
    ele[22][7] != ele[22][24];
    ele[22][7] != ele[22][25];
    ele[22][7] != ele[22][26];
    ele[22][7] != ele[22][27];
    ele[22][7] != ele[22][28];
    ele[22][7] != ele[22][29];
    ele[22][7] != ele[22][30];
    ele[22][7] != ele[22][31];
    ele[22][7] != ele[22][32];
    ele[22][7] != ele[22][33];
    ele[22][7] != ele[22][34];
    ele[22][7] != ele[22][35];
    ele[22][7] != ele[22][8];
    ele[22][7] != ele[22][9];
    ele[22][7] != ele[23][10];
    ele[22][7] != ele[23][11];
    ele[22][7] != ele[23][6];
    ele[22][7] != ele[23][7];
    ele[22][7] != ele[23][8];
    ele[22][7] != ele[23][9];
    ele[22][7] != ele[24][7];
    ele[22][7] != ele[25][7];
    ele[22][7] != ele[26][7];
    ele[22][7] != ele[27][7];
    ele[22][7] != ele[28][7];
    ele[22][7] != ele[29][7];
    ele[22][7] != ele[30][7];
    ele[22][7] != ele[31][7];
    ele[22][7] != ele[32][7];
    ele[22][7] != ele[33][7];
    ele[22][7] != ele[34][7];
    ele[22][7] != ele[35][7];
    ele[22][8] != ele[22][10];
    ele[22][8] != ele[22][11];
    ele[22][8] != ele[22][12];
    ele[22][8] != ele[22][13];
    ele[22][8] != ele[22][14];
    ele[22][8] != ele[22][15];
    ele[22][8] != ele[22][16];
    ele[22][8] != ele[22][17];
    ele[22][8] != ele[22][18];
    ele[22][8] != ele[22][19];
    ele[22][8] != ele[22][20];
    ele[22][8] != ele[22][21];
    ele[22][8] != ele[22][22];
    ele[22][8] != ele[22][23];
    ele[22][8] != ele[22][24];
    ele[22][8] != ele[22][25];
    ele[22][8] != ele[22][26];
    ele[22][8] != ele[22][27];
    ele[22][8] != ele[22][28];
    ele[22][8] != ele[22][29];
    ele[22][8] != ele[22][30];
    ele[22][8] != ele[22][31];
    ele[22][8] != ele[22][32];
    ele[22][8] != ele[22][33];
    ele[22][8] != ele[22][34];
    ele[22][8] != ele[22][35];
    ele[22][8] != ele[22][9];
    ele[22][8] != ele[23][10];
    ele[22][8] != ele[23][11];
    ele[22][8] != ele[23][6];
    ele[22][8] != ele[23][7];
    ele[22][8] != ele[23][8];
    ele[22][8] != ele[23][9];
    ele[22][8] != ele[24][8];
    ele[22][8] != ele[25][8];
    ele[22][8] != ele[26][8];
    ele[22][8] != ele[27][8];
    ele[22][8] != ele[28][8];
    ele[22][8] != ele[29][8];
    ele[22][8] != ele[30][8];
    ele[22][8] != ele[31][8];
    ele[22][8] != ele[32][8];
    ele[22][8] != ele[33][8];
    ele[22][8] != ele[34][8];
    ele[22][8] != ele[35][8];
    ele[22][9] != ele[22][10];
    ele[22][9] != ele[22][11];
    ele[22][9] != ele[22][12];
    ele[22][9] != ele[22][13];
    ele[22][9] != ele[22][14];
    ele[22][9] != ele[22][15];
    ele[22][9] != ele[22][16];
    ele[22][9] != ele[22][17];
    ele[22][9] != ele[22][18];
    ele[22][9] != ele[22][19];
    ele[22][9] != ele[22][20];
    ele[22][9] != ele[22][21];
    ele[22][9] != ele[22][22];
    ele[22][9] != ele[22][23];
    ele[22][9] != ele[22][24];
    ele[22][9] != ele[22][25];
    ele[22][9] != ele[22][26];
    ele[22][9] != ele[22][27];
    ele[22][9] != ele[22][28];
    ele[22][9] != ele[22][29];
    ele[22][9] != ele[22][30];
    ele[22][9] != ele[22][31];
    ele[22][9] != ele[22][32];
    ele[22][9] != ele[22][33];
    ele[22][9] != ele[22][34];
    ele[22][9] != ele[22][35];
    ele[22][9] != ele[23][10];
    ele[22][9] != ele[23][11];
    ele[22][9] != ele[23][6];
    ele[22][9] != ele[23][7];
    ele[22][9] != ele[23][8];
    ele[22][9] != ele[23][9];
    ele[22][9] != ele[24][9];
    ele[22][9] != ele[25][9];
    ele[22][9] != ele[26][9];
    ele[22][9] != ele[27][9];
    ele[22][9] != ele[28][9];
    ele[22][9] != ele[29][9];
    ele[22][9] != ele[30][9];
    ele[22][9] != ele[31][9];
    ele[22][9] != ele[32][9];
    ele[22][9] != ele[33][9];
    ele[22][9] != ele[34][9];
    ele[22][9] != ele[35][9];
    ele[23][0] != ele[23][1];
    ele[23][0] != ele[23][10];
    ele[23][0] != ele[23][11];
    ele[23][0] != ele[23][12];
    ele[23][0] != ele[23][13];
    ele[23][0] != ele[23][14];
    ele[23][0] != ele[23][15];
    ele[23][0] != ele[23][16];
    ele[23][0] != ele[23][17];
    ele[23][0] != ele[23][18];
    ele[23][0] != ele[23][19];
    ele[23][0] != ele[23][2];
    ele[23][0] != ele[23][20];
    ele[23][0] != ele[23][21];
    ele[23][0] != ele[23][22];
    ele[23][0] != ele[23][23];
    ele[23][0] != ele[23][24];
    ele[23][0] != ele[23][25];
    ele[23][0] != ele[23][26];
    ele[23][0] != ele[23][27];
    ele[23][0] != ele[23][28];
    ele[23][0] != ele[23][29];
    ele[23][0] != ele[23][3];
    ele[23][0] != ele[23][30];
    ele[23][0] != ele[23][31];
    ele[23][0] != ele[23][32];
    ele[23][0] != ele[23][33];
    ele[23][0] != ele[23][34];
    ele[23][0] != ele[23][35];
    ele[23][0] != ele[23][4];
    ele[23][0] != ele[23][5];
    ele[23][0] != ele[23][6];
    ele[23][0] != ele[23][7];
    ele[23][0] != ele[23][8];
    ele[23][0] != ele[23][9];
    ele[23][0] != ele[24][0];
    ele[23][0] != ele[25][0];
    ele[23][0] != ele[26][0];
    ele[23][0] != ele[27][0];
    ele[23][0] != ele[28][0];
    ele[23][0] != ele[29][0];
    ele[23][0] != ele[30][0];
    ele[23][0] != ele[31][0];
    ele[23][0] != ele[32][0];
    ele[23][0] != ele[33][0];
    ele[23][0] != ele[34][0];
    ele[23][0] != ele[35][0];
    ele[23][1] != ele[23][10];
    ele[23][1] != ele[23][11];
    ele[23][1] != ele[23][12];
    ele[23][1] != ele[23][13];
    ele[23][1] != ele[23][14];
    ele[23][1] != ele[23][15];
    ele[23][1] != ele[23][16];
    ele[23][1] != ele[23][17];
    ele[23][1] != ele[23][18];
    ele[23][1] != ele[23][19];
    ele[23][1] != ele[23][2];
    ele[23][1] != ele[23][20];
    ele[23][1] != ele[23][21];
    ele[23][1] != ele[23][22];
    ele[23][1] != ele[23][23];
    ele[23][1] != ele[23][24];
    ele[23][1] != ele[23][25];
    ele[23][1] != ele[23][26];
    ele[23][1] != ele[23][27];
    ele[23][1] != ele[23][28];
    ele[23][1] != ele[23][29];
    ele[23][1] != ele[23][3];
    ele[23][1] != ele[23][30];
    ele[23][1] != ele[23][31];
    ele[23][1] != ele[23][32];
    ele[23][1] != ele[23][33];
    ele[23][1] != ele[23][34];
    ele[23][1] != ele[23][35];
    ele[23][1] != ele[23][4];
    ele[23][1] != ele[23][5];
    ele[23][1] != ele[23][6];
    ele[23][1] != ele[23][7];
    ele[23][1] != ele[23][8];
    ele[23][1] != ele[23][9];
    ele[23][1] != ele[24][1];
    ele[23][1] != ele[25][1];
    ele[23][1] != ele[26][1];
    ele[23][1] != ele[27][1];
    ele[23][1] != ele[28][1];
    ele[23][1] != ele[29][1];
    ele[23][1] != ele[30][1];
    ele[23][1] != ele[31][1];
    ele[23][1] != ele[32][1];
    ele[23][1] != ele[33][1];
    ele[23][1] != ele[34][1];
    ele[23][1] != ele[35][1];
    ele[23][10] != ele[23][11];
    ele[23][10] != ele[23][12];
    ele[23][10] != ele[23][13];
    ele[23][10] != ele[23][14];
    ele[23][10] != ele[23][15];
    ele[23][10] != ele[23][16];
    ele[23][10] != ele[23][17];
    ele[23][10] != ele[23][18];
    ele[23][10] != ele[23][19];
    ele[23][10] != ele[23][20];
    ele[23][10] != ele[23][21];
    ele[23][10] != ele[23][22];
    ele[23][10] != ele[23][23];
    ele[23][10] != ele[23][24];
    ele[23][10] != ele[23][25];
    ele[23][10] != ele[23][26];
    ele[23][10] != ele[23][27];
    ele[23][10] != ele[23][28];
    ele[23][10] != ele[23][29];
    ele[23][10] != ele[23][30];
    ele[23][10] != ele[23][31];
    ele[23][10] != ele[23][32];
    ele[23][10] != ele[23][33];
    ele[23][10] != ele[23][34];
    ele[23][10] != ele[23][35];
    ele[23][10] != ele[24][10];
    ele[23][10] != ele[25][10];
    ele[23][10] != ele[26][10];
    ele[23][10] != ele[27][10];
    ele[23][10] != ele[28][10];
    ele[23][10] != ele[29][10];
    ele[23][10] != ele[30][10];
    ele[23][10] != ele[31][10];
    ele[23][10] != ele[32][10];
    ele[23][10] != ele[33][10];
    ele[23][10] != ele[34][10];
    ele[23][10] != ele[35][10];
    ele[23][11] != ele[23][12];
    ele[23][11] != ele[23][13];
    ele[23][11] != ele[23][14];
    ele[23][11] != ele[23][15];
    ele[23][11] != ele[23][16];
    ele[23][11] != ele[23][17];
    ele[23][11] != ele[23][18];
    ele[23][11] != ele[23][19];
    ele[23][11] != ele[23][20];
    ele[23][11] != ele[23][21];
    ele[23][11] != ele[23][22];
    ele[23][11] != ele[23][23];
    ele[23][11] != ele[23][24];
    ele[23][11] != ele[23][25];
    ele[23][11] != ele[23][26];
    ele[23][11] != ele[23][27];
    ele[23][11] != ele[23][28];
    ele[23][11] != ele[23][29];
    ele[23][11] != ele[23][30];
    ele[23][11] != ele[23][31];
    ele[23][11] != ele[23][32];
    ele[23][11] != ele[23][33];
    ele[23][11] != ele[23][34];
    ele[23][11] != ele[23][35];
    ele[23][11] != ele[24][11];
    ele[23][11] != ele[25][11];
    ele[23][11] != ele[26][11];
    ele[23][11] != ele[27][11];
    ele[23][11] != ele[28][11];
    ele[23][11] != ele[29][11];
    ele[23][11] != ele[30][11];
    ele[23][11] != ele[31][11];
    ele[23][11] != ele[32][11];
    ele[23][11] != ele[33][11];
    ele[23][11] != ele[34][11];
    ele[23][11] != ele[35][11];
    ele[23][12] != ele[23][13];
    ele[23][12] != ele[23][14];
    ele[23][12] != ele[23][15];
    ele[23][12] != ele[23][16];
    ele[23][12] != ele[23][17];
    ele[23][12] != ele[23][18];
    ele[23][12] != ele[23][19];
    ele[23][12] != ele[23][20];
    ele[23][12] != ele[23][21];
    ele[23][12] != ele[23][22];
    ele[23][12] != ele[23][23];
    ele[23][12] != ele[23][24];
    ele[23][12] != ele[23][25];
    ele[23][12] != ele[23][26];
    ele[23][12] != ele[23][27];
    ele[23][12] != ele[23][28];
    ele[23][12] != ele[23][29];
    ele[23][12] != ele[23][30];
    ele[23][12] != ele[23][31];
    ele[23][12] != ele[23][32];
    ele[23][12] != ele[23][33];
    ele[23][12] != ele[23][34];
    ele[23][12] != ele[23][35];
    ele[23][12] != ele[24][12];
    ele[23][12] != ele[25][12];
    ele[23][12] != ele[26][12];
    ele[23][12] != ele[27][12];
    ele[23][12] != ele[28][12];
    ele[23][12] != ele[29][12];
    ele[23][12] != ele[30][12];
    ele[23][12] != ele[31][12];
    ele[23][12] != ele[32][12];
    ele[23][12] != ele[33][12];
    ele[23][12] != ele[34][12];
    ele[23][12] != ele[35][12];
    ele[23][13] != ele[23][14];
    ele[23][13] != ele[23][15];
    ele[23][13] != ele[23][16];
    ele[23][13] != ele[23][17];
    ele[23][13] != ele[23][18];
    ele[23][13] != ele[23][19];
    ele[23][13] != ele[23][20];
    ele[23][13] != ele[23][21];
    ele[23][13] != ele[23][22];
    ele[23][13] != ele[23][23];
    ele[23][13] != ele[23][24];
    ele[23][13] != ele[23][25];
    ele[23][13] != ele[23][26];
    ele[23][13] != ele[23][27];
    ele[23][13] != ele[23][28];
    ele[23][13] != ele[23][29];
    ele[23][13] != ele[23][30];
    ele[23][13] != ele[23][31];
    ele[23][13] != ele[23][32];
    ele[23][13] != ele[23][33];
    ele[23][13] != ele[23][34];
    ele[23][13] != ele[23][35];
    ele[23][13] != ele[24][13];
    ele[23][13] != ele[25][13];
    ele[23][13] != ele[26][13];
    ele[23][13] != ele[27][13];
    ele[23][13] != ele[28][13];
    ele[23][13] != ele[29][13];
    ele[23][13] != ele[30][13];
    ele[23][13] != ele[31][13];
    ele[23][13] != ele[32][13];
    ele[23][13] != ele[33][13];
    ele[23][13] != ele[34][13];
    ele[23][13] != ele[35][13];
    ele[23][14] != ele[23][15];
    ele[23][14] != ele[23][16];
    ele[23][14] != ele[23][17];
    ele[23][14] != ele[23][18];
    ele[23][14] != ele[23][19];
    ele[23][14] != ele[23][20];
    ele[23][14] != ele[23][21];
    ele[23][14] != ele[23][22];
    ele[23][14] != ele[23][23];
    ele[23][14] != ele[23][24];
    ele[23][14] != ele[23][25];
    ele[23][14] != ele[23][26];
    ele[23][14] != ele[23][27];
    ele[23][14] != ele[23][28];
    ele[23][14] != ele[23][29];
    ele[23][14] != ele[23][30];
    ele[23][14] != ele[23][31];
    ele[23][14] != ele[23][32];
    ele[23][14] != ele[23][33];
    ele[23][14] != ele[23][34];
    ele[23][14] != ele[23][35];
    ele[23][14] != ele[24][14];
    ele[23][14] != ele[25][14];
    ele[23][14] != ele[26][14];
    ele[23][14] != ele[27][14];
    ele[23][14] != ele[28][14];
    ele[23][14] != ele[29][14];
    ele[23][14] != ele[30][14];
    ele[23][14] != ele[31][14];
    ele[23][14] != ele[32][14];
    ele[23][14] != ele[33][14];
    ele[23][14] != ele[34][14];
    ele[23][14] != ele[35][14];
    ele[23][15] != ele[23][16];
    ele[23][15] != ele[23][17];
    ele[23][15] != ele[23][18];
    ele[23][15] != ele[23][19];
    ele[23][15] != ele[23][20];
    ele[23][15] != ele[23][21];
    ele[23][15] != ele[23][22];
    ele[23][15] != ele[23][23];
    ele[23][15] != ele[23][24];
    ele[23][15] != ele[23][25];
    ele[23][15] != ele[23][26];
    ele[23][15] != ele[23][27];
    ele[23][15] != ele[23][28];
    ele[23][15] != ele[23][29];
    ele[23][15] != ele[23][30];
    ele[23][15] != ele[23][31];
    ele[23][15] != ele[23][32];
    ele[23][15] != ele[23][33];
    ele[23][15] != ele[23][34];
    ele[23][15] != ele[23][35];
    ele[23][15] != ele[24][15];
    ele[23][15] != ele[25][15];
    ele[23][15] != ele[26][15];
    ele[23][15] != ele[27][15];
    ele[23][15] != ele[28][15];
    ele[23][15] != ele[29][15];
    ele[23][15] != ele[30][15];
    ele[23][15] != ele[31][15];
    ele[23][15] != ele[32][15];
    ele[23][15] != ele[33][15];
    ele[23][15] != ele[34][15];
    ele[23][15] != ele[35][15];
    ele[23][16] != ele[23][17];
    ele[23][16] != ele[23][18];
    ele[23][16] != ele[23][19];
    ele[23][16] != ele[23][20];
    ele[23][16] != ele[23][21];
    ele[23][16] != ele[23][22];
    ele[23][16] != ele[23][23];
    ele[23][16] != ele[23][24];
    ele[23][16] != ele[23][25];
    ele[23][16] != ele[23][26];
    ele[23][16] != ele[23][27];
    ele[23][16] != ele[23][28];
    ele[23][16] != ele[23][29];
    ele[23][16] != ele[23][30];
    ele[23][16] != ele[23][31];
    ele[23][16] != ele[23][32];
    ele[23][16] != ele[23][33];
    ele[23][16] != ele[23][34];
    ele[23][16] != ele[23][35];
    ele[23][16] != ele[24][16];
    ele[23][16] != ele[25][16];
    ele[23][16] != ele[26][16];
    ele[23][16] != ele[27][16];
    ele[23][16] != ele[28][16];
    ele[23][16] != ele[29][16];
    ele[23][16] != ele[30][16];
    ele[23][16] != ele[31][16];
    ele[23][16] != ele[32][16];
    ele[23][16] != ele[33][16];
    ele[23][16] != ele[34][16];
    ele[23][16] != ele[35][16];
    ele[23][17] != ele[23][18];
    ele[23][17] != ele[23][19];
    ele[23][17] != ele[23][20];
    ele[23][17] != ele[23][21];
    ele[23][17] != ele[23][22];
    ele[23][17] != ele[23][23];
    ele[23][17] != ele[23][24];
    ele[23][17] != ele[23][25];
    ele[23][17] != ele[23][26];
    ele[23][17] != ele[23][27];
    ele[23][17] != ele[23][28];
    ele[23][17] != ele[23][29];
    ele[23][17] != ele[23][30];
    ele[23][17] != ele[23][31];
    ele[23][17] != ele[23][32];
    ele[23][17] != ele[23][33];
    ele[23][17] != ele[23][34];
    ele[23][17] != ele[23][35];
    ele[23][17] != ele[24][17];
    ele[23][17] != ele[25][17];
    ele[23][17] != ele[26][17];
    ele[23][17] != ele[27][17];
    ele[23][17] != ele[28][17];
    ele[23][17] != ele[29][17];
    ele[23][17] != ele[30][17];
    ele[23][17] != ele[31][17];
    ele[23][17] != ele[32][17];
    ele[23][17] != ele[33][17];
    ele[23][17] != ele[34][17];
    ele[23][17] != ele[35][17];
    ele[23][18] != ele[23][19];
    ele[23][18] != ele[23][20];
    ele[23][18] != ele[23][21];
    ele[23][18] != ele[23][22];
    ele[23][18] != ele[23][23];
    ele[23][18] != ele[23][24];
    ele[23][18] != ele[23][25];
    ele[23][18] != ele[23][26];
    ele[23][18] != ele[23][27];
    ele[23][18] != ele[23][28];
    ele[23][18] != ele[23][29];
    ele[23][18] != ele[23][30];
    ele[23][18] != ele[23][31];
    ele[23][18] != ele[23][32];
    ele[23][18] != ele[23][33];
    ele[23][18] != ele[23][34];
    ele[23][18] != ele[23][35];
    ele[23][18] != ele[24][18];
    ele[23][18] != ele[25][18];
    ele[23][18] != ele[26][18];
    ele[23][18] != ele[27][18];
    ele[23][18] != ele[28][18];
    ele[23][18] != ele[29][18];
    ele[23][18] != ele[30][18];
    ele[23][18] != ele[31][18];
    ele[23][18] != ele[32][18];
    ele[23][18] != ele[33][18];
    ele[23][18] != ele[34][18];
    ele[23][18] != ele[35][18];
    ele[23][19] != ele[23][20];
    ele[23][19] != ele[23][21];
    ele[23][19] != ele[23][22];
    ele[23][19] != ele[23][23];
    ele[23][19] != ele[23][24];
    ele[23][19] != ele[23][25];
    ele[23][19] != ele[23][26];
    ele[23][19] != ele[23][27];
    ele[23][19] != ele[23][28];
    ele[23][19] != ele[23][29];
    ele[23][19] != ele[23][30];
    ele[23][19] != ele[23][31];
    ele[23][19] != ele[23][32];
    ele[23][19] != ele[23][33];
    ele[23][19] != ele[23][34];
    ele[23][19] != ele[23][35];
    ele[23][19] != ele[24][19];
    ele[23][19] != ele[25][19];
    ele[23][19] != ele[26][19];
    ele[23][19] != ele[27][19];
    ele[23][19] != ele[28][19];
    ele[23][19] != ele[29][19];
    ele[23][19] != ele[30][19];
    ele[23][19] != ele[31][19];
    ele[23][19] != ele[32][19];
    ele[23][19] != ele[33][19];
    ele[23][19] != ele[34][19];
    ele[23][19] != ele[35][19];
    ele[23][2] != ele[23][10];
    ele[23][2] != ele[23][11];
    ele[23][2] != ele[23][12];
    ele[23][2] != ele[23][13];
    ele[23][2] != ele[23][14];
    ele[23][2] != ele[23][15];
    ele[23][2] != ele[23][16];
    ele[23][2] != ele[23][17];
    ele[23][2] != ele[23][18];
    ele[23][2] != ele[23][19];
    ele[23][2] != ele[23][20];
    ele[23][2] != ele[23][21];
    ele[23][2] != ele[23][22];
    ele[23][2] != ele[23][23];
    ele[23][2] != ele[23][24];
    ele[23][2] != ele[23][25];
    ele[23][2] != ele[23][26];
    ele[23][2] != ele[23][27];
    ele[23][2] != ele[23][28];
    ele[23][2] != ele[23][29];
    ele[23][2] != ele[23][3];
    ele[23][2] != ele[23][30];
    ele[23][2] != ele[23][31];
    ele[23][2] != ele[23][32];
    ele[23][2] != ele[23][33];
    ele[23][2] != ele[23][34];
    ele[23][2] != ele[23][35];
    ele[23][2] != ele[23][4];
    ele[23][2] != ele[23][5];
    ele[23][2] != ele[23][6];
    ele[23][2] != ele[23][7];
    ele[23][2] != ele[23][8];
    ele[23][2] != ele[23][9];
    ele[23][2] != ele[24][2];
    ele[23][2] != ele[25][2];
    ele[23][2] != ele[26][2];
    ele[23][2] != ele[27][2];
    ele[23][2] != ele[28][2];
    ele[23][2] != ele[29][2];
    ele[23][2] != ele[30][2];
    ele[23][2] != ele[31][2];
    ele[23][2] != ele[32][2];
    ele[23][2] != ele[33][2];
    ele[23][2] != ele[34][2];
    ele[23][2] != ele[35][2];
    ele[23][20] != ele[23][21];
    ele[23][20] != ele[23][22];
    ele[23][20] != ele[23][23];
    ele[23][20] != ele[23][24];
    ele[23][20] != ele[23][25];
    ele[23][20] != ele[23][26];
    ele[23][20] != ele[23][27];
    ele[23][20] != ele[23][28];
    ele[23][20] != ele[23][29];
    ele[23][20] != ele[23][30];
    ele[23][20] != ele[23][31];
    ele[23][20] != ele[23][32];
    ele[23][20] != ele[23][33];
    ele[23][20] != ele[23][34];
    ele[23][20] != ele[23][35];
    ele[23][20] != ele[24][20];
    ele[23][20] != ele[25][20];
    ele[23][20] != ele[26][20];
    ele[23][20] != ele[27][20];
    ele[23][20] != ele[28][20];
    ele[23][20] != ele[29][20];
    ele[23][20] != ele[30][20];
    ele[23][20] != ele[31][20];
    ele[23][20] != ele[32][20];
    ele[23][20] != ele[33][20];
    ele[23][20] != ele[34][20];
    ele[23][20] != ele[35][20];
    ele[23][21] != ele[23][22];
    ele[23][21] != ele[23][23];
    ele[23][21] != ele[23][24];
    ele[23][21] != ele[23][25];
    ele[23][21] != ele[23][26];
    ele[23][21] != ele[23][27];
    ele[23][21] != ele[23][28];
    ele[23][21] != ele[23][29];
    ele[23][21] != ele[23][30];
    ele[23][21] != ele[23][31];
    ele[23][21] != ele[23][32];
    ele[23][21] != ele[23][33];
    ele[23][21] != ele[23][34];
    ele[23][21] != ele[23][35];
    ele[23][21] != ele[24][21];
    ele[23][21] != ele[25][21];
    ele[23][21] != ele[26][21];
    ele[23][21] != ele[27][21];
    ele[23][21] != ele[28][21];
    ele[23][21] != ele[29][21];
    ele[23][21] != ele[30][21];
    ele[23][21] != ele[31][21];
    ele[23][21] != ele[32][21];
    ele[23][21] != ele[33][21];
    ele[23][21] != ele[34][21];
    ele[23][21] != ele[35][21];
    ele[23][22] != ele[23][23];
    ele[23][22] != ele[23][24];
    ele[23][22] != ele[23][25];
    ele[23][22] != ele[23][26];
    ele[23][22] != ele[23][27];
    ele[23][22] != ele[23][28];
    ele[23][22] != ele[23][29];
    ele[23][22] != ele[23][30];
    ele[23][22] != ele[23][31];
    ele[23][22] != ele[23][32];
    ele[23][22] != ele[23][33];
    ele[23][22] != ele[23][34];
    ele[23][22] != ele[23][35];
    ele[23][22] != ele[24][22];
    ele[23][22] != ele[25][22];
    ele[23][22] != ele[26][22];
    ele[23][22] != ele[27][22];
    ele[23][22] != ele[28][22];
    ele[23][22] != ele[29][22];
    ele[23][22] != ele[30][22];
    ele[23][22] != ele[31][22];
    ele[23][22] != ele[32][22];
    ele[23][22] != ele[33][22];
    ele[23][22] != ele[34][22];
    ele[23][22] != ele[35][22];
    ele[23][23] != ele[23][24];
    ele[23][23] != ele[23][25];
    ele[23][23] != ele[23][26];
    ele[23][23] != ele[23][27];
    ele[23][23] != ele[23][28];
    ele[23][23] != ele[23][29];
    ele[23][23] != ele[23][30];
    ele[23][23] != ele[23][31];
    ele[23][23] != ele[23][32];
    ele[23][23] != ele[23][33];
    ele[23][23] != ele[23][34];
    ele[23][23] != ele[23][35];
    ele[23][23] != ele[24][23];
    ele[23][23] != ele[25][23];
    ele[23][23] != ele[26][23];
    ele[23][23] != ele[27][23];
    ele[23][23] != ele[28][23];
    ele[23][23] != ele[29][23];
    ele[23][23] != ele[30][23];
    ele[23][23] != ele[31][23];
    ele[23][23] != ele[32][23];
    ele[23][23] != ele[33][23];
    ele[23][23] != ele[34][23];
    ele[23][23] != ele[35][23];
    ele[23][24] != ele[23][25];
    ele[23][24] != ele[23][26];
    ele[23][24] != ele[23][27];
    ele[23][24] != ele[23][28];
    ele[23][24] != ele[23][29];
    ele[23][24] != ele[23][30];
    ele[23][24] != ele[23][31];
    ele[23][24] != ele[23][32];
    ele[23][24] != ele[23][33];
    ele[23][24] != ele[23][34];
    ele[23][24] != ele[23][35];
    ele[23][24] != ele[24][24];
    ele[23][24] != ele[25][24];
    ele[23][24] != ele[26][24];
    ele[23][24] != ele[27][24];
    ele[23][24] != ele[28][24];
    ele[23][24] != ele[29][24];
    ele[23][24] != ele[30][24];
    ele[23][24] != ele[31][24];
    ele[23][24] != ele[32][24];
    ele[23][24] != ele[33][24];
    ele[23][24] != ele[34][24];
    ele[23][24] != ele[35][24];
    ele[23][25] != ele[23][26];
    ele[23][25] != ele[23][27];
    ele[23][25] != ele[23][28];
    ele[23][25] != ele[23][29];
    ele[23][25] != ele[23][30];
    ele[23][25] != ele[23][31];
    ele[23][25] != ele[23][32];
    ele[23][25] != ele[23][33];
    ele[23][25] != ele[23][34];
    ele[23][25] != ele[23][35];
    ele[23][25] != ele[24][25];
    ele[23][25] != ele[25][25];
    ele[23][25] != ele[26][25];
    ele[23][25] != ele[27][25];
    ele[23][25] != ele[28][25];
    ele[23][25] != ele[29][25];
    ele[23][25] != ele[30][25];
    ele[23][25] != ele[31][25];
    ele[23][25] != ele[32][25];
    ele[23][25] != ele[33][25];
    ele[23][25] != ele[34][25];
    ele[23][25] != ele[35][25];
    ele[23][26] != ele[23][27];
    ele[23][26] != ele[23][28];
    ele[23][26] != ele[23][29];
    ele[23][26] != ele[23][30];
    ele[23][26] != ele[23][31];
    ele[23][26] != ele[23][32];
    ele[23][26] != ele[23][33];
    ele[23][26] != ele[23][34];
    ele[23][26] != ele[23][35];
    ele[23][26] != ele[24][26];
    ele[23][26] != ele[25][26];
    ele[23][26] != ele[26][26];
    ele[23][26] != ele[27][26];
    ele[23][26] != ele[28][26];
    ele[23][26] != ele[29][26];
    ele[23][26] != ele[30][26];
    ele[23][26] != ele[31][26];
    ele[23][26] != ele[32][26];
    ele[23][26] != ele[33][26];
    ele[23][26] != ele[34][26];
    ele[23][26] != ele[35][26];
    ele[23][27] != ele[23][28];
    ele[23][27] != ele[23][29];
    ele[23][27] != ele[23][30];
    ele[23][27] != ele[23][31];
    ele[23][27] != ele[23][32];
    ele[23][27] != ele[23][33];
    ele[23][27] != ele[23][34];
    ele[23][27] != ele[23][35];
    ele[23][27] != ele[24][27];
    ele[23][27] != ele[25][27];
    ele[23][27] != ele[26][27];
    ele[23][27] != ele[27][27];
    ele[23][27] != ele[28][27];
    ele[23][27] != ele[29][27];
    ele[23][27] != ele[30][27];
    ele[23][27] != ele[31][27];
    ele[23][27] != ele[32][27];
    ele[23][27] != ele[33][27];
    ele[23][27] != ele[34][27];
    ele[23][27] != ele[35][27];
    ele[23][28] != ele[23][29];
    ele[23][28] != ele[23][30];
    ele[23][28] != ele[23][31];
    ele[23][28] != ele[23][32];
    ele[23][28] != ele[23][33];
    ele[23][28] != ele[23][34];
    ele[23][28] != ele[23][35];
    ele[23][28] != ele[24][28];
    ele[23][28] != ele[25][28];
    ele[23][28] != ele[26][28];
    ele[23][28] != ele[27][28];
    ele[23][28] != ele[28][28];
    ele[23][28] != ele[29][28];
    ele[23][28] != ele[30][28];
    ele[23][28] != ele[31][28];
    ele[23][28] != ele[32][28];
    ele[23][28] != ele[33][28];
    ele[23][28] != ele[34][28];
    ele[23][28] != ele[35][28];
    ele[23][29] != ele[23][30];
    ele[23][29] != ele[23][31];
    ele[23][29] != ele[23][32];
    ele[23][29] != ele[23][33];
    ele[23][29] != ele[23][34];
    ele[23][29] != ele[23][35];
    ele[23][29] != ele[24][29];
    ele[23][29] != ele[25][29];
    ele[23][29] != ele[26][29];
    ele[23][29] != ele[27][29];
    ele[23][29] != ele[28][29];
    ele[23][29] != ele[29][29];
    ele[23][29] != ele[30][29];
    ele[23][29] != ele[31][29];
    ele[23][29] != ele[32][29];
    ele[23][29] != ele[33][29];
    ele[23][29] != ele[34][29];
    ele[23][29] != ele[35][29];
    ele[23][3] != ele[23][10];
    ele[23][3] != ele[23][11];
    ele[23][3] != ele[23][12];
    ele[23][3] != ele[23][13];
    ele[23][3] != ele[23][14];
    ele[23][3] != ele[23][15];
    ele[23][3] != ele[23][16];
    ele[23][3] != ele[23][17];
    ele[23][3] != ele[23][18];
    ele[23][3] != ele[23][19];
    ele[23][3] != ele[23][20];
    ele[23][3] != ele[23][21];
    ele[23][3] != ele[23][22];
    ele[23][3] != ele[23][23];
    ele[23][3] != ele[23][24];
    ele[23][3] != ele[23][25];
    ele[23][3] != ele[23][26];
    ele[23][3] != ele[23][27];
    ele[23][3] != ele[23][28];
    ele[23][3] != ele[23][29];
    ele[23][3] != ele[23][30];
    ele[23][3] != ele[23][31];
    ele[23][3] != ele[23][32];
    ele[23][3] != ele[23][33];
    ele[23][3] != ele[23][34];
    ele[23][3] != ele[23][35];
    ele[23][3] != ele[23][4];
    ele[23][3] != ele[23][5];
    ele[23][3] != ele[23][6];
    ele[23][3] != ele[23][7];
    ele[23][3] != ele[23][8];
    ele[23][3] != ele[23][9];
    ele[23][3] != ele[24][3];
    ele[23][3] != ele[25][3];
    ele[23][3] != ele[26][3];
    ele[23][3] != ele[27][3];
    ele[23][3] != ele[28][3];
    ele[23][3] != ele[29][3];
    ele[23][3] != ele[30][3];
    ele[23][3] != ele[31][3];
    ele[23][3] != ele[32][3];
    ele[23][3] != ele[33][3];
    ele[23][3] != ele[34][3];
    ele[23][3] != ele[35][3];
    ele[23][30] != ele[23][31];
    ele[23][30] != ele[23][32];
    ele[23][30] != ele[23][33];
    ele[23][30] != ele[23][34];
    ele[23][30] != ele[23][35];
    ele[23][30] != ele[24][30];
    ele[23][30] != ele[25][30];
    ele[23][30] != ele[26][30];
    ele[23][30] != ele[27][30];
    ele[23][30] != ele[28][30];
    ele[23][30] != ele[29][30];
    ele[23][30] != ele[30][30];
    ele[23][30] != ele[31][30];
    ele[23][30] != ele[32][30];
    ele[23][30] != ele[33][30];
    ele[23][30] != ele[34][30];
    ele[23][30] != ele[35][30];
    ele[23][31] != ele[23][32];
    ele[23][31] != ele[23][33];
    ele[23][31] != ele[23][34];
    ele[23][31] != ele[23][35];
    ele[23][31] != ele[24][31];
    ele[23][31] != ele[25][31];
    ele[23][31] != ele[26][31];
    ele[23][31] != ele[27][31];
    ele[23][31] != ele[28][31];
    ele[23][31] != ele[29][31];
    ele[23][31] != ele[30][31];
    ele[23][31] != ele[31][31];
    ele[23][31] != ele[32][31];
    ele[23][31] != ele[33][31];
    ele[23][31] != ele[34][31];
    ele[23][31] != ele[35][31];
    ele[23][32] != ele[23][33];
    ele[23][32] != ele[23][34];
    ele[23][32] != ele[23][35];
    ele[23][32] != ele[24][32];
    ele[23][32] != ele[25][32];
    ele[23][32] != ele[26][32];
    ele[23][32] != ele[27][32];
    ele[23][32] != ele[28][32];
    ele[23][32] != ele[29][32];
    ele[23][32] != ele[30][32];
    ele[23][32] != ele[31][32];
    ele[23][32] != ele[32][32];
    ele[23][32] != ele[33][32];
    ele[23][32] != ele[34][32];
    ele[23][32] != ele[35][32];
    ele[23][33] != ele[23][34];
    ele[23][33] != ele[23][35];
    ele[23][33] != ele[24][33];
    ele[23][33] != ele[25][33];
    ele[23][33] != ele[26][33];
    ele[23][33] != ele[27][33];
    ele[23][33] != ele[28][33];
    ele[23][33] != ele[29][33];
    ele[23][33] != ele[30][33];
    ele[23][33] != ele[31][33];
    ele[23][33] != ele[32][33];
    ele[23][33] != ele[33][33];
    ele[23][33] != ele[34][33];
    ele[23][33] != ele[35][33];
    ele[23][34] != ele[23][35];
    ele[23][34] != ele[24][34];
    ele[23][34] != ele[25][34];
    ele[23][34] != ele[26][34];
    ele[23][34] != ele[27][34];
    ele[23][34] != ele[28][34];
    ele[23][34] != ele[29][34];
    ele[23][34] != ele[30][34];
    ele[23][34] != ele[31][34];
    ele[23][34] != ele[32][34];
    ele[23][34] != ele[33][34];
    ele[23][34] != ele[34][34];
    ele[23][34] != ele[35][34];
    ele[23][35] != ele[24][35];
    ele[23][35] != ele[25][35];
    ele[23][35] != ele[26][35];
    ele[23][35] != ele[27][35];
    ele[23][35] != ele[28][35];
    ele[23][35] != ele[29][35];
    ele[23][35] != ele[30][35];
    ele[23][35] != ele[31][35];
    ele[23][35] != ele[32][35];
    ele[23][35] != ele[33][35];
    ele[23][35] != ele[34][35];
    ele[23][35] != ele[35][35];
    ele[23][4] != ele[23][10];
    ele[23][4] != ele[23][11];
    ele[23][4] != ele[23][12];
    ele[23][4] != ele[23][13];
    ele[23][4] != ele[23][14];
    ele[23][4] != ele[23][15];
    ele[23][4] != ele[23][16];
    ele[23][4] != ele[23][17];
    ele[23][4] != ele[23][18];
    ele[23][4] != ele[23][19];
    ele[23][4] != ele[23][20];
    ele[23][4] != ele[23][21];
    ele[23][4] != ele[23][22];
    ele[23][4] != ele[23][23];
    ele[23][4] != ele[23][24];
    ele[23][4] != ele[23][25];
    ele[23][4] != ele[23][26];
    ele[23][4] != ele[23][27];
    ele[23][4] != ele[23][28];
    ele[23][4] != ele[23][29];
    ele[23][4] != ele[23][30];
    ele[23][4] != ele[23][31];
    ele[23][4] != ele[23][32];
    ele[23][4] != ele[23][33];
    ele[23][4] != ele[23][34];
    ele[23][4] != ele[23][35];
    ele[23][4] != ele[23][5];
    ele[23][4] != ele[23][6];
    ele[23][4] != ele[23][7];
    ele[23][4] != ele[23][8];
    ele[23][4] != ele[23][9];
    ele[23][4] != ele[24][4];
    ele[23][4] != ele[25][4];
    ele[23][4] != ele[26][4];
    ele[23][4] != ele[27][4];
    ele[23][4] != ele[28][4];
    ele[23][4] != ele[29][4];
    ele[23][4] != ele[30][4];
    ele[23][4] != ele[31][4];
    ele[23][4] != ele[32][4];
    ele[23][4] != ele[33][4];
    ele[23][4] != ele[34][4];
    ele[23][4] != ele[35][4];
    ele[23][5] != ele[23][10];
    ele[23][5] != ele[23][11];
    ele[23][5] != ele[23][12];
    ele[23][5] != ele[23][13];
    ele[23][5] != ele[23][14];
    ele[23][5] != ele[23][15];
    ele[23][5] != ele[23][16];
    ele[23][5] != ele[23][17];
    ele[23][5] != ele[23][18];
    ele[23][5] != ele[23][19];
    ele[23][5] != ele[23][20];
    ele[23][5] != ele[23][21];
    ele[23][5] != ele[23][22];
    ele[23][5] != ele[23][23];
    ele[23][5] != ele[23][24];
    ele[23][5] != ele[23][25];
    ele[23][5] != ele[23][26];
    ele[23][5] != ele[23][27];
    ele[23][5] != ele[23][28];
    ele[23][5] != ele[23][29];
    ele[23][5] != ele[23][30];
    ele[23][5] != ele[23][31];
    ele[23][5] != ele[23][32];
    ele[23][5] != ele[23][33];
    ele[23][5] != ele[23][34];
    ele[23][5] != ele[23][35];
    ele[23][5] != ele[23][6];
    ele[23][5] != ele[23][7];
    ele[23][5] != ele[23][8];
    ele[23][5] != ele[23][9];
    ele[23][5] != ele[24][5];
    ele[23][5] != ele[25][5];
    ele[23][5] != ele[26][5];
    ele[23][5] != ele[27][5];
    ele[23][5] != ele[28][5];
    ele[23][5] != ele[29][5];
    ele[23][5] != ele[30][5];
    ele[23][5] != ele[31][5];
    ele[23][5] != ele[32][5];
    ele[23][5] != ele[33][5];
    ele[23][5] != ele[34][5];
    ele[23][5] != ele[35][5];
    ele[23][6] != ele[23][10];
    ele[23][6] != ele[23][11];
    ele[23][6] != ele[23][12];
    ele[23][6] != ele[23][13];
    ele[23][6] != ele[23][14];
    ele[23][6] != ele[23][15];
    ele[23][6] != ele[23][16];
    ele[23][6] != ele[23][17];
    ele[23][6] != ele[23][18];
    ele[23][6] != ele[23][19];
    ele[23][6] != ele[23][20];
    ele[23][6] != ele[23][21];
    ele[23][6] != ele[23][22];
    ele[23][6] != ele[23][23];
    ele[23][6] != ele[23][24];
    ele[23][6] != ele[23][25];
    ele[23][6] != ele[23][26];
    ele[23][6] != ele[23][27];
    ele[23][6] != ele[23][28];
    ele[23][6] != ele[23][29];
    ele[23][6] != ele[23][30];
    ele[23][6] != ele[23][31];
    ele[23][6] != ele[23][32];
    ele[23][6] != ele[23][33];
    ele[23][6] != ele[23][34];
    ele[23][6] != ele[23][35];
    ele[23][6] != ele[23][7];
    ele[23][6] != ele[23][8];
    ele[23][6] != ele[23][9];
    ele[23][6] != ele[24][6];
    ele[23][6] != ele[25][6];
    ele[23][6] != ele[26][6];
    ele[23][6] != ele[27][6];
    ele[23][6] != ele[28][6];
    ele[23][6] != ele[29][6];
    ele[23][6] != ele[30][6];
    ele[23][6] != ele[31][6];
    ele[23][6] != ele[32][6];
    ele[23][6] != ele[33][6];
    ele[23][6] != ele[34][6];
    ele[23][6] != ele[35][6];
    ele[23][7] != ele[23][10];
    ele[23][7] != ele[23][11];
    ele[23][7] != ele[23][12];
    ele[23][7] != ele[23][13];
    ele[23][7] != ele[23][14];
    ele[23][7] != ele[23][15];
    ele[23][7] != ele[23][16];
    ele[23][7] != ele[23][17];
    ele[23][7] != ele[23][18];
    ele[23][7] != ele[23][19];
    ele[23][7] != ele[23][20];
    ele[23][7] != ele[23][21];
    ele[23][7] != ele[23][22];
    ele[23][7] != ele[23][23];
    ele[23][7] != ele[23][24];
    ele[23][7] != ele[23][25];
    ele[23][7] != ele[23][26];
    ele[23][7] != ele[23][27];
    ele[23][7] != ele[23][28];
    ele[23][7] != ele[23][29];
    ele[23][7] != ele[23][30];
    ele[23][7] != ele[23][31];
    ele[23][7] != ele[23][32];
    ele[23][7] != ele[23][33];
    ele[23][7] != ele[23][34];
    ele[23][7] != ele[23][35];
    ele[23][7] != ele[23][8];
    ele[23][7] != ele[23][9];
    ele[23][7] != ele[24][7];
    ele[23][7] != ele[25][7];
    ele[23][7] != ele[26][7];
    ele[23][7] != ele[27][7];
    ele[23][7] != ele[28][7];
    ele[23][7] != ele[29][7];
    ele[23][7] != ele[30][7];
    ele[23][7] != ele[31][7];
    ele[23][7] != ele[32][7];
    ele[23][7] != ele[33][7];
    ele[23][7] != ele[34][7];
    ele[23][7] != ele[35][7];
    ele[23][8] != ele[23][10];
    ele[23][8] != ele[23][11];
    ele[23][8] != ele[23][12];
    ele[23][8] != ele[23][13];
    ele[23][8] != ele[23][14];
    ele[23][8] != ele[23][15];
    ele[23][8] != ele[23][16];
    ele[23][8] != ele[23][17];
    ele[23][8] != ele[23][18];
    ele[23][8] != ele[23][19];
    ele[23][8] != ele[23][20];
    ele[23][8] != ele[23][21];
    ele[23][8] != ele[23][22];
    ele[23][8] != ele[23][23];
    ele[23][8] != ele[23][24];
    ele[23][8] != ele[23][25];
    ele[23][8] != ele[23][26];
    ele[23][8] != ele[23][27];
    ele[23][8] != ele[23][28];
    ele[23][8] != ele[23][29];
    ele[23][8] != ele[23][30];
    ele[23][8] != ele[23][31];
    ele[23][8] != ele[23][32];
    ele[23][8] != ele[23][33];
    ele[23][8] != ele[23][34];
    ele[23][8] != ele[23][35];
    ele[23][8] != ele[23][9];
    ele[23][8] != ele[24][8];
    ele[23][8] != ele[25][8];
    ele[23][8] != ele[26][8];
    ele[23][8] != ele[27][8];
    ele[23][8] != ele[28][8];
    ele[23][8] != ele[29][8];
    ele[23][8] != ele[30][8];
    ele[23][8] != ele[31][8];
    ele[23][8] != ele[32][8];
    ele[23][8] != ele[33][8];
    ele[23][8] != ele[34][8];
    ele[23][8] != ele[35][8];
    ele[23][9] != ele[23][10];
    ele[23][9] != ele[23][11];
    ele[23][9] != ele[23][12];
    ele[23][9] != ele[23][13];
    ele[23][9] != ele[23][14];
    ele[23][9] != ele[23][15];
    ele[23][9] != ele[23][16];
    ele[23][9] != ele[23][17];
    ele[23][9] != ele[23][18];
    ele[23][9] != ele[23][19];
    ele[23][9] != ele[23][20];
    ele[23][9] != ele[23][21];
    ele[23][9] != ele[23][22];
    ele[23][9] != ele[23][23];
    ele[23][9] != ele[23][24];
    ele[23][9] != ele[23][25];
    ele[23][9] != ele[23][26];
    ele[23][9] != ele[23][27];
    ele[23][9] != ele[23][28];
    ele[23][9] != ele[23][29];
    ele[23][9] != ele[23][30];
    ele[23][9] != ele[23][31];
    ele[23][9] != ele[23][32];
    ele[23][9] != ele[23][33];
    ele[23][9] != ele[23][34];
    ele[23][9] != ele[23][35];
    ele[23][9] != ele[24][9];
    ele[23][9] != ele[25][9];
    ele[23][9] != ele[26][9];
    ele[23][9] != ele[27][9];
    ele[23][9] != ele[28][9];
    ele[23][9] != ele[29][9];
    ele[23][9] != ele[30][9];
    ele[23][9] != ele[31][9];
    ele[23][9] != ele[32][9];
    ele[23][9] != ele[33][9];
    ele[23][9] != ele[34][9];
    ele[23][9] != ele[35][9];
    ele[24][0] != ele[24][1];
    ele[24][0] != ele[24][10];
    ele[24][0] != ele[24][11];
    ele[24][0] != ele[24][12];
    ele[24][0] != ele[24][13];
    ele[24][0] != ele[24][14];
    ele[24][0] != ele[24][15];
    ele[24][0] != ele[24][16];
    ele[24][0] != ele[24][17];
    ele[24][0] != ele[24][18];
    ele[24][0] != ele[24][19];
    ele[24][0] != ele[24][2];
    ele[24][0] != ele[24][20];
    ele[24][0] != ele[24][21];
    ele[24][0] != ele[24][22];
    ele[24][0] != ele[24][23];
    ele[24][0] != ele[24][24];
    ele[24][0] != ele[24][25];
    ele[24][0] != ele[24][26];
    ele[24][0] != ele[24][27];
    ele[24][0] != ele[24][28];
    ele[24][0] != ele[24][29];
    ele[24][0] != ele[24][3];
    ele[24][0] != ele[24][30];
    ele[24][0] != ele[24][31];
    ele[24][0] != ele[24][32];
    ele[24][0] != ele[24][33];
    ele[24][0] != ele[24][34];
    ele[24][0] != ele[24][35];
    ele[24][0] != ele[24][4];
    ele[24][0] != ele[24][5];
    ele[24][0] != ele[24][6];
    ele[24][0] != ele[24][7];
    ele[24][0] != ele[24][8];
    ele[24][0] != ele[24][9];
    ele[24][0] != ele[25][0];
    ele[24][0] != ele[25][1];
    ele[24][0] != ele[25][2];
    ele[24][0] != ele[25][3];
    ele[24][0] != ele[25][4];
    ele[24][0] != ele[25][5];
    ele[24][0] != ele[26][0];
    ele[24][0] != ele[26][1];
    ele[24][0] != ele[26][2];
    ele[24][0] != ele[26][3];
    ele[24][0] != ele[26][4];
    ele[24][0] != ele[26][5];
    ele[24][0] != ele[27][0];
    ele[24][0] != ele[27][1];
    ele[24][0] != ele[27][2];
    ele[24][0] != ele[27][3];
    ele[24][0] != ele[27][4];
    ele[24][0] != ele[27][5];
    ele[24][0] != ele[28][0];
    ele[24][0] != ele[28][1];
    ele[24][0] != ele[28][2];
    ele[24][0] != ele[28][3];
    ele[24][0] != ele[28][4];
    ele[24][0] != ele[28][5];
    ele[24][0] != ele[29][0];
    ele[24][0] != ele[29][1];
    ele[24][0] != ele[29][2];
    ele[24][0] != ele[29][3];
    ele[24][0] != ele[29][4];
    ele[24][0] != ele[29][5];
    ele[24][0] != ele[30][0];
    ele[24][0] != ele[31][0];
    ele[24][0] != ele[32][0];
    ele[24][0] != ele[33][0];
    ele[24][0] != ele[34][0];
    ele[24][0] != ele[35][0];
    ele[24][1] != ele[24][10];
    ele[24][1] != ele[24][11];
    ele[24][1] != ele[24][12];
    ele[24][1] != ele[24][13];
    ele[24][1] != ele[24][14];
    ele[24][1] != ele[24][15];
    ele[24][1] != ele[24][16];
    ele[24][1] != ele[24][17];
    ele[24][1] != ele[24][18];
    ele[24][1] != ele[24][19];
    ele[24][1] != ele[24][2];
    ele[24][1] != ele[24][20];
    ele[24][1] != ele[24][21];
    ele[24][1] != ele[24][22];
    ele[24][1] != ele[24][23];
    ele[24][1] != ele[24][24];
    ele[24][1] != ele[24][25];
    ele[24][1] != ele[24][26];
    ele[24][1] != ele[24][27];
    ele[24][1] != ele[24][28];
    ele[24][1] != ele[24][29];
    ele[24][1] != ele[24][3];
    ele[24][1] != ele[24][30];
    ele[24][1] != ele[24][31];
    ele[24][1] != ele[24][32];
    ele[24][1] != ele[24][33];
    ele[24][1] != ele[24][34];
    ele[24][1] != ele[24][35];
    ele[24][1] != ele[24][4];
    ele[24][1] != ele[24][5];
    ele[24][1] != ele[24][6];
    ele[24][1] != ele[24][7];
    ele[24][1] != ele[24][8];
    ele[24][1] != ele[24][9];
    ele[24][1] != ele[25][0];
    ele[24][1] != ele[25][1];
    ele[24][1] != ele[25][2];
    ele[24][1] != ele[25][3];
    ele[24][1] != ele[25][4];
    ele[24][1] != ele[25][5];
    ele[24][1] != ele[26][0];
    ele[24][1] != ele[26][1];
    ele[24][1] != ele[26][2];
    ele[24][1] != ele[26][3];
    ele[24][1] != ele[26][4];
    ele[24][1] != ele[26][5];
    ele[24][1] != ele[27][0];
    ele[24][1] != ele[27][1];
    ele[24][1] != ele[27][2];
    ele[24][1] != ele[27][3];
    ele[24][1] != ele[27][4];
    ele[24][1] != ele[27][5];
    ele[24][1] != ele[28][0];
    ele[24][1] != ele[28][1];
    ele[24][1] != ele[28][2];
    ele[24][1] != ele[28][3];
    ele[24][1] != ele[28][4];
    ele[24][1] != ele[28][5];
    ele[24][1] != ele[29][0];
    ele[24][1] != ele[29][1];
    ele[24][1] != ele[29][2];
    ele[24][1] != ele[29][3];
    ele[24][1] != ele[29][4];
    ele[24][1] != ele[29][5];
    ele[24][1] != ele[30][1];
    ele[24][1] != ele[31][1];
    ele[24][1] != ele[32][1];
    ele[24][1] != ele[33][1];
    ele[24][1] != ele[34][1];
    ele[24][1] != ele[35][1];
    ele[24][10] != ele[24][11];
    ele[24][10] != ele[24][12];
    ele[24][10] != ele[24][13];
    ele[24][10] != ele[24][14];
    ele[24][10] != ele[24][15];
    ele[24][10] != ele[24][16];
    ele[24][10] != ele[24][17];
    ele[24][10] != ele[24][18];
    ele[24][10] != ele[24][19];
    ele[24][10] != ele[24][20];
    ele[24][10] != ele[24][21];
    ele[24][10] != ele[24][22];
    ele[24][10] != ele[24][23];
    ele[24][10] != ele[24][24];
    ele[24][10] != ele[24][25];
    ele[24][10] != ele[24][26];
    ele[24][10] != ele[24][27];
    ele[24][10] != ele[24][28];
    ele[24][10] != ele[24][29];
    ele[24][10] != ele[24][30];
    ele[24][10] != ele[24][31];
    ele[24][10] != ele[24][32];
    ele[24][10] != ele[24][33];
    ele[24][10] != ele[24][34];
    ele[24][10] != ele[24][35];
    ele[24][10] != ele[25][10];
    ele[24][10] != ele[25][11];
    ele[24][10] != ele[25][6];
    ele[24][10] != ele[25][7];
    ele[24][10] != ele[25][8];
    ele[24][10] != ele[25][9];
    ele[24][10] != ele[26][10];
    ele[24][10] != ele[26][11];
    ele[24][10] != ele[26][6];
    ele[24][10] != ele[26][7];
    ele[24][10] != ele[26][8];
    ele[24][10] != ele[26][9];
    ele[24][10] != ele[27][10];
    ele[24][10] != ele[27][11];
    ele[24][10] != ele[27][6];
    ele[24][10] != ele[27][7];
    ele[24][10] != ele[27][8];
    ele[24][10] != ele[27][9];
    ele[24][10] != ele[28][10];
    ele[24][10] != ele[28][11];
    ele[24][10] != ele[28][6];
    ele[24][10] != ele[28][7];
    ele[24][10] != ele[28][8];
    ele[24][10] != ele[28][9];
    ele[24][10] != ele[29][10];
    ele[24][10] != ele[29][11];
    ele[24][10] != ele[29][6];
    ele[24][10] != ele[29][7];
    ele[24][10] != ele[29][8];
    ele[24][10] != ele[29][9];
    ele[24][10] != ele[30][10];
    ele[24][10] != ele[31][10];
    ele[24][10] != ele[32][10];
    ele[24][10] != ele[33][10];
    ele[24][10] != ele[34][10];
    ele[24][10] != ele[35][10];
    ele[24][11] != ele[24][12];
    ele[24][11] != ele[24][13];
    ele[24][11] != ele[24][14];
    ele[24][11] != ele[24][15];
    ele[24][11] != ele[24][16];
    ele[24][11] != ele[24][17];
    ele[24][11] != ele[24][18];
    ele[24][11] != ele[24][19];
    ele[24][11] != ele[24][20];
    ele[24][11] != ele[24][21];
    ele[24][11] != ele[24][22];
    ele[24][11] != ele[24][23];
    ele[24][11] != ele[24][24];
    ele[24][11] != ele[24][25];
    ele[24][11] != ele[24][26];
    ele[24][11] != ele[24][27];
    ele[24][11] != ele[24][28];
    ele[24][11] != ele[24][29];
    ele[24][11] != ele[24][30];
    ele[24][11] != ele[24][31];
    ele[24][11] != ele[24][32];
    ele[24][11] != ele[24][33];
    ele[24][11] != ele[24][34];
    ele[24][11] != ele[24][35];
    ele[24][11] != ele[25][10];
    ele[24][11] != ele[25][11];
    ele[24][11] != ele[25][6];
    ele[24][11] != ele[25][7];
    ele[24][11] != ele[25][8];
    ele[24][11] != ele[25][9];
    ele[24][11] != ele[26][10];
    ele[24][11] != ele[26][11];
    ele[24][11] != ele[26][6];
    ele[24][11] != ele[26][7];
    ele[24][11] != ele[26][8];
    ele[24][11] != ele[26][9];
    ele[24][11] != ele[27][10];
    ele[24][11] != ele[27][11];
    ele[24][11] != ele[27][6];
    ele[24][11] != ele[27][7];
    ele[24][11] != ele[27][8];
    ele[24][11] != ele[27][9];
    ele[24][11] != ele[28][10];
    ele[24][11] != ele[28][11];
    ele[24][11] != ele[28][6];
    ele[24][11] != ele[28][7];
    ele[24][11] != ele[28][8];
    ele[24][11] != ele[28][9];
    ele[24][11] != ele[29][10];
    ele[24][11] != ele[29][11];
    ele[24][11] != ele[29][6];
    ele[24][11] != ele[29][7];
    ele[24][11] != ele[29][8];
    ele[24][11] != ele[29][9];
    ele[24][11] != ele[30][11];
    ele[24][11] != ele[31][11];
    ele[24][11] != ele[32][11];
    ele[24][11] != ele[33][11];
    ele[24][11] != ele[34][11];
    ele[24][11] != ele[35][11];
    ele[24][12] != ele[24][13];
    ele[24][12] != ele[24][14];
    ele[24][12] != ele[24][15];
    ele[24][12] != ele[24][16];
    ele[24][12] != ele[24][17];
    ele[24][12] != ele[24][18];
    ele[24][12] != ele[24][19];
    ele[24][12] != ele[24][20];
    ele[24][12] != ele[24][21];
    ele[24][12] != ele[24][22];
    ele[24][12] != ele[24][23];
    ele[24][12] != ele[24][24];
    ele[24][12] != ele[24][25];
    ele[24][12] != ele[24][26];
    ele[24][12] != ele[24][27];
    ele[24][12] != ele[24][28];
    ele[24][12] != ele[24][29];
    ele[24][12] != ele[24][30];
    ele[24][12] != ele[24][31];
    ele[24][12] != ele[24][32];
    ele[24][12] != ele[24][33];
    ele[24][12] != ele[24][34];
    ele[24][12] != ele[24][35];
    ele[24][12] != ele[25][12];
    ele[24][12] != ele[25][13];
    ele[24][12] != ele[25][14];
    ele[24][12] != ele[25][15];
    ele[24][12] != ele[25][16];
    ele[24][12] != ele[25][17];
    ele[24][12] != ele[26][12];
    ele[24][12] != ele[26][13];
    ele[24][12] != ele[26][14];
    ele[24][12] != ele[26][15];
    ele[24][12] != ele[26][16];
    ele[24][12] != ele[26][17];
    ele[24][12] != ele[27][12];
    ele[24][12] != ele[27][13];
    ele[24][12] != ele[27][14];
    ele[24][12] != ele[27][15];
    ele[24][12] != ele[27][16];
    ele[24][12] != ele[27][17];
    ele[24][12] != ele[28][12];
    ele[24][12] != ele[28][13];
    ele[24][12] != ele[28][14];
    ele[24][12] != ele[28][15];
    ele[24][12] != ele[28][16];
    ele[24][12] != ele[28][17];
    ele[24][12] != ele[29][12];
    ele[24][12] != ele[29][13];
    ele[24][12] != ele[29][14];
    ele[24][12] != ele[29][15];
    ele[24][12] != ele[29][16];
    ele[24][12] != ele[29][17];
    ele[24][12] != ele[30][12];
    ele[24][12] != ele[31][12];
    ele[24][12] != ele[32][12];
    ele[24][12] != ele[33][12];
    ele[24][12] != ele[34][12];
    ele[24][12] != ele[35][12];
    ele[24][13] != ele[24][14];
    ele[24][13] != ele[24][15];
    ele[24][13] != ele[24][16];
    ele[24][13] != ele[24][17];
    ele[24][13] != ele[24][18];
    ele[24][13] != ele[24][19];
    ele[24][13] != ele[24][20];
    ele[24][13] != ele[24][21];
    ele[24][13] != ele[24][22];
    ele[24][13] != ele[24][23];
    ele[24][13] != ele[24][24];
    ele[24][13] != ele[24][25];
    ele[24][13] != ele[24][26];
    ele[24][13] != ele[24][27];
    ele[24][13] != ele[24][28];
    ele[24][13] != ele[24][29];
    ele[24][13] != ele[24][30];
    ele[24][13] != ele[24][31];
    ele[24][13] != ele[24][32];
    ele[24][13] != ele[24][33];
    ele[24][13] != ele[24][34];
    ele[24][13] != ele[24][35];
    ele[24][13] != ele[25][12];
    ele[24][13] != ele[25][13];
    ele[24][13] != ele[25][14];
    ele[24][13] != ele[25][15];
    ele[24][13] != ele[25][16];
    ele[24][13] != ele[25][17];
    ele[24][13] != ele[26][12];
    ele[24][13] != ele[26][13];
    ele[24][13] != ele[26][14];
    ele[24][13] != ele[26][15];
    ele[24][13] != ele[26][16];
    ele[24][13] != ele[26][17];
    ele[24][13] != ele[27][12];
    ele[24][13] != ele[27][13];
    ele[24][13] != ele[27][14];
    ele[24][13] != ele[27][15];
    ele[24][13] != ele[27][16];
    ele[24][13] != ele[27][17];
    ele[24][13] != ele[28][12];
    ele[24][13] != ele[28][13];
    ele[24][13] != ele[28][14];
    ele[24][13] != ele[28][15];
    ele[24][13] != ele[28][16];
    ele[24][13] != ele[28][17];
    ele[24][13] != ele[29][12];
    ele[24][13] != ele[29][13];
    ele[24][13] != ele[29][14];
    ele[24][13] != ele[29][15];
    ele[24][13] != ele[29][16];
    ele[24][13] != ele[29][17];
    ele[24][13] != ele[30][13];
    ele[24][13] != ele[31][13];
    ele[24][13] != ele[32][13];
    ele[24][13] != ele[33][13];
    ele[24][13] != ele[34][13];
    ele[24][13] != ele[35][13];
    ele[24][14] != ele[24][15];
    ele[24][14] != ele[24][16];
    ele[24][14] != ele[24][17];
    ele[24][14] != ele[24][18];
    ele[24][14] != ele[24][19];
    ele[24][14] != ele[24][20];
    ele[24][14] != ele[24][21];
    ele[24][14] != ele[24][22];
    ele[24][14] != ele[24][23];
    ele[24][14] != ele[24][24];
    ele[24][14] != ele[24][25];
    ele[24][14] != ele[24][26];
    ele[24][14] != ele[24][27];
    ele[24][14] != ele[24][28];
    ele[24][14] != ele[24][29];
    ele[24][14] != ele[24][30];
    ele[24][14] != ele[24][31];
    ele[24][14] != ele[24][32];
    ele[24][14] != ele[24][33];
    ele[24][14] != ele[24][34];
    ele[24][14] != ele[24][35];
    ele[24][14] != ele[25][12];
    ele[24][14] != ele[25][13];
    ele[24][14] != ele[25][14];
    ele[24][14] != ele[25][15];
    ele[24][14] != ele[25][16];
    ele[24][14] != ele[25][17];
    ele[24][14] != ele[26][12];
    ele[24][14] != ele[26][13];
    ele[24][14] != ele[26][14];
    ele[24][14] != ele[26][15];
    ele[24][14] != ele[26][16];
    ele[24][14] != ele[26][17];
    ele[24][14] != ele[27][12];
    ele[24][14] != ele[27][13];
    ele[24][14] != ele[27][14];
    ele[24][14] != ele[27][15];
    ele[24][14] != ele[27][16];
    ele[24][14] != ele[27][17];
    ele[24][14] != ele[28][12];
    ele[24][14] != ele[28][13];
    ele[24][14] != ele[28][14];
    ele[24][14] != ele[28][15];
    ele[24][14] != ele[28][16];
    ele[24][14] != ele[28][17];
    ele[24][14] != ele[29][12];
    ele[24][14] != ele[29][13];
    ele[24][14] != ele[29][14];
    ele[24][14] != ele[29][15];
    ele[24][14] != ele[29][16];
    ele[24][14] != ele[29][17];
    ele[24][14] != ele[30][14];
    ele[24][14] != ele[31][14];
    ele[24][14] != ele[32][14];
    ele[24][14] != ele[33][14];
    ele[24][14] != ele[34][14];
    ele[24][14] != ele[35][14];
    ele[24][15] != ele[24][16];
    ele[24][15] != ele[24][17];
    ele[24][15] != ele[24][18];
    ele[24][15] != ele[24][19];
    ele[24][15] != ele[24][20];
    ele[24][15] != ele[24][21];
    ele[24][15] != ele[24][22];
    ele[24][15] != ele[24][23];
    ele[24][15] != ele[24][24];
    ele[24][15] != ele[24][25];
    ele[24][15] != ele[24][26];
    ele[24][15] != ele[24][27];
    ele[24][15] != ele[24][28];
    ele[24][15] != ele[24][29];
    ele[24][15] != ele[24][30];
    ele[24][15] != ele[24][31];
    ele[24][15] != ele[24][32];
    ele[24][15] != ele[24][33];
    ele[24][15] != ele[24][34];
    ele[24][15] != ele[24][35];
    ele[24][15] != ele[25][12];
    ele[24][15] != ele[25][13];
    ele[24][15] != ele[25][14];
    ele[24][15] != ele[25][15];
    ele[24][15] != ele[25][16];
    ele[24][15] != ele[25][17];
    ele[24][15] != ele[26][12];
    ele[24][15] != ele[26][13];
    ele[24][15] != ele[26][14];
    ele[24][15] != ele[26][15];
    ele[24][15] != ele[26][16];
    ele[24][15] != ele[26][17];
    ele[24][15] != ele[27][12];
    ele[24][15] != ele[27][13];
    ele[24][15] != ele[27][14];
    ele[24][15] != ele[27][15];
    ele[24][15] != ele[27][16];
    ele[24][15] != ele[27][17];
    ele[24][15] != ele[28][12];
    ele[24][15] != ele[28][13];
    ele[24][15] != ele[28][14];
    ele[24][15] != ele[28][15];
    ele[24][15] != ele[28][16];
    ele[24][15] != ele[28][17];
    ele[24][15] != ele[29][12];
    ele[24][15] != ele[29][13];
    ele[24][15] != ele[29][14];
    ele[24][15] != ele[29][15];
    ele[24][15] != ele[29][16];
    ele[24][15] != ele[29][17];
    ele[24][15] != ele[30][15];
    ele[24][15] != ele[31][15];
    ele[24][15] != ele[32][15];
    ele[24][15] != ele[33][15];
    ele[24][15] != ele[34][15];
    ele[24][15] != ele[35][15];
    ele[24][16] != ele[24][17];
    ele[24][16] != ele[24][18];
    ele[24][16] != ele[24][19];
    ele[24][16] != ele[24][20];
    ele[24][16] != ele[24][21];
    ele[24][16] != ele[24][22];
    ele[24][16] != ele[24][23];
    ele[24][16] != ele[24][24];
    ele[24][16] != ele[24][25];
    ele[24][16] != ele[24][26];
    ele[24][16] != ele[24][27];
    ele[24][16] != ele[24][28];
    ele[24][16] != ele[24][29];
    ele[24][16] != ele[24][30];
    ele[24][16] != ele[24][31];
    ele[24][16] != ele[24][32];
    ele[24][16] != ele[24][33];
    ele[24][16] != ele[24][34];
    ele[24][16] != ele[24][35];
    ele[24][16] != ele[25][12];
    ele[24][16] != ele[25][13];
    ele[24][16] != ele[25][14];
    ele[24][16] != ele[25][15];
    ele[24][16] != ele[25][16];
    ele[24][16] != ele[25][17];
    ele[24][16] != ele[26][12];
    ele[24][16] != ele[26][13];
    ele[24][16] != ele[26][14];
    ele[24][16] != ele[26][15];
    ele[24][16] != ele[26][16];
    ele[24][16] != ele[26][17];
    ele[24][16] != ele[27][12];
    ele[24][16] != ele[27][13];
    ele[24][16] != ele[27][14];
    ele[24][16] != ele[27][15];
    ele[24][16] != ele[27][16];
    ele[24][16] != ele[27][17];
    ele[24][16] != ele[28][12];
    ele[24][16] != ele[28][13];
    ele[24][16] != ele[28][14];
    ele[24][16] != ele[28][15];
    ele[24][16] != ele[28][16];
    ele[24][16] != ele[28][17];
    ele[24][16] != ele[29][12];
    ele[24][16] != ele[29][13];
    ele[24][16] != ele[29][14];
    ele[24][16] != ele[29][15];
    ele[24][16] != ele[29][16];
    ele[24][16] != ele[29][17];
    ele[24][16] != ele[30][16];
    ele[24][16] != ele[31][16];
    ele[24][16] != ele[32][16];
    ele[24][16] != ele[33][16];
    ele[24][16] != ele[34][16];
    ele[24][16] != ele[35][16];
    ele[24][17] != ele[24][18];
    ele[24][17] != ele[24][19];
    ele[24][17] != ele[24][20];
    ele[24][17] != ele[24][21];
    ele[24][17] != ele[24][22];
    ele[24][17] != ele[24][23];
    ele[24][17] != ele[24][24];
    ele[24][17] != ele[24][25];
    ele[24][17] != ele[24][26];
    ele[24][17] != ele[24][27];
    ele[24][17] != ele[24][28];
    ele[24][17] != ele[24][29];
    ele[24][17] != ele[24][30];
    ele[24][17] != ele[24][31];
    ele[24][17] != ele[24][32];
    ele[24][17] != ele[24][33];
    ele[24][17] != ele[24][34];
    ele[24][17] != ele[24][35];
    ele[24][17] != ele[25][12];
    ele[24][17] != ele[25][13];
    ele[24][17] != ele[25][14];
    ele[24][17] != ele[25][15];
    ele[24][17] != ele[25][16];
    ele[24][17] != ele[25][17];
    ele[24][17] != ele[26][12];
    ele[24][17] != ele[26][13];
    ele[24][17] != ele[26][14];
    ele[24][17] != ele[26][15];
    ele[24][17] != ele[26][16];
    ele[24][17] != ele[26][17];
    ele[24][17] != ele[27][12];
    ele[24][17] != ele[27][13];
    ele[24][17] != ele[27][14];
    ele[24][17] != ele[27][15];
    ele[24][17] != ele[27][16];
    ele[24][17] != ele[27][17];
    ele[24][17] != ele[28][12];
    ele[24][17] != ele[28][13];
    ele[24][17] != ele[28][14];
    ele[24][17] != ele[28][15];
    ele[24][17] != ele[28][16];
    ele[24][17] != ele[28][17];
    ele[24][17] != ele[29][12];
    ele[24][17] != ele[29][13];
    ele[24][17] != ele[29][14];
    ele[24][17] != ele[29][15];
    ele[24][17] != ele[29][16];
    ele[24][17] != ele[29][17];
    ele[24][17] != ele[30][17];
    ele[24][17] != ele[31][17];
    ele[24][17] != ele[32][17];
    ele[24][17] != ele[33][17];
    ele[24][17] != ele[34][17];
    ele[24][17] != ele[35][17];
    ele[24][18] != ele[24][19];
    ele[24][18] != ele[24][20];
    ele[24][18] != ele[24][21];
    ele[24][18] != ele[24][22];
    ele[24][18] != ele[24][23];
    ele[24][18] != ele[24][24];
    ele[24][18] != ele[24][25];
    ele[24][18] != ele[24][26];
    ele[24][18] != ele[24][27];
    ele[24][18] != ele[24][28];
    ele[24][18] != ele[24][29];
    ele[24][18] != ele[24][30];
    ele[24][18] != ele[24][31];
    ele[24][18] != ele[24][32];
    ele[24][18] != ele[24][33];
    ele[24][18] != ele[24][34];
    ele[24][18] != ele[24][35];
    ele[24][18] != ele[25][18];
    ele[24][18] != ele[25][19];
    ele[24][18] != ele[25][20];
    ele[24][18] != ele[25][21];
    ele[24][18] != ele[25][22];
    ele[24][18] != ele[25][23];
    ele[24][18] != ele[26][18];
    ele[24][18] != ele[26][19];
    ele[24][18] != ele[26][20];
    ele[24][18] != ele[26][21];
    ele[24][18] != ele[26][22];
    ele[24][18] != ele[26][23];
    ele[24][18] != ele[27][18];
    ele[24][18] != ele[27][19];
    ele[24][18] != ele[27][20];
    ele[24][18] != ele[27][21];
    ele[24][18] != ele[27][22];
    ele[24][18] != ele[27][23];
    ele[24][18] != ele[28][18];
    ele[24][18] != ele[28][19];
    ele[24][18] != ele[28][20];
    ele[24][18] != ele[28][21];
    ele[24][18] != ele[28][22];
    ele[24][18] != ele[28][23];
    ele[24][18] != ele[29][18];
    ele[24][18] != ele[29][19];
    ele[24][18] != ele[29][20];
    ele[24][18] != ele[29][21];
    ele[24][18] != ele[29][22];
    ele[24][18] != ele[29][23];
    ele[24][18] != ele[30][18];
    ele[24][18] != ele[31][18];
    ele[24][18] != ele[32][18];
    ele[24][18] != ele[33][18];
    ele[24][18] != ele[34][18];
    ele[24][18] != ele[35][18];
    ele[24][19] != ele[24][20];
    ele[24][19] != ele[24][21];
    ele[24][19] != ele[24][22];
    ele[24][19] != ele[24][23];
    ele[24][19] != ele[24][24];
    ele[24][19] != ele[24][25];
    ele[24][19] != ele[24][26];
    ele[24][19] != ele[24][27];
    ele[24][19] != ele[24][28];
    ele[24][19] != ele[24][29];
    ele[24][19] != ele[24][30];
    ele[24][19] != ele[24][31];
    ele[24][19] != ele[24][32];
    ele[24][19] != ele[24][33];
    ele[24][19] != ele[24][34];
    ele[24][19] != ele[24][35];
    ele[24][19] != ele[25][18];
    ele[24][19] != ele[25][19];
    ele[24][19] != ele[25][20];
    ele[24][19] != ele[25][21];
    ele[24][19] != ele[25][22];
    ele[24][19] != ele[25][23];
    ele[24][19] != ele[26][18];
    ele[24][19] != ele[26][19];
    ele[24][19] != ele[26][20];
    ele[24][19] != ele[26][21];
    ele[24][19] != ele[26][22];
    ele[24][19] != ele[26][23];
    ele[24][19] != ele[27][18];
    ele[24][19] != ele[27][19];
    ele[24][19] != ele[27][20];
    ele[24][19] != ele[27][21];
    ele[24][19] != ele[27][22];
    ele[24][19] != ele[27][23];
    ele[24][19] != ele[28][18];
    ele[24][19] != ele[28][19];
    ele[24][19] != ele[28][20];
    ele[24][19] != ele[28][21];
    ele[24][19] != ele[28][22];
    ele[24][19] != ele[28][23];
    ele[24][19] != ele[29][18];
    ele[24][19] != ele[29][19];
    ele[24][19] != ele[29][20];
    ele[24][19] != ele[29][21];
    ele[24][19] != ele[29][22];
    ele[24][19] != ele[29][23];
    ele[24][19] != ele[30][19];
    ele[24][19] != ele[31][19];
    ele[24][19] != ele[32][19];
    ele[24][19] != ele[33][19];
    ele[24][19] != ele[34][19];
    ele[24][19] != ele[35][19];
    ele[24][2] != ele[24][10];
    ele[24][2] != ele[24][11];
    ele[24][2] != ele[24][12];
    ele[24][2] != ele[24][13];
    ele[24][2] != ele[24][14];
    ele[24][2] != ele[24][15];
    ele[24][2] != ele[24][16];
    ele[24][2] != ele[24][17];
    ele[24][2] != ele[24][18];
    ele[24][2] != ele[24][19];
    ele[24][2] != ele[24][20];
    ele[24][2] != ele[24][21];
    ele[24][2] != ele[24][22];
    ele[24][2] != ele[24][23];
    ele[24][2] != ele[24][24];
    ele[24][2] != ele[24][25];
    ele[24][2] != ele[24][26];
    ele[24][2] != ele[24][27];
    ele[24][2] != ele[24][28];
    ele[24][2] != ele[24][29];
    ele[24][2] != ele[24][3];
    ele[24][2] != ele[24][30];
    ele[24][2] != ele[24][31];
    ele[24][2] != ele[24][32];
    ele[24][2] != ele[24][33];
    ele[24][2] != ele[24][34];
    ele[24][2] != ele[24][35];
    ele[24][2] != ele[24][4];
    ele[24][2] != ele[24][5];
    ele[24][2] != ele[24][6];
    ele[24][2] != ele[24][7];
    ele[24][2] != ele[24][8];
    ele[24][2] != ele[24][9];
    ele[24][2] != ele[25][0];
    ele[24][2] != ele[25][1];
    ele[24][2] != ele[25][2];
    ele[24][2] != ele[25][3];
    ele[24][2] != ele[25][4];
    ele[24][2] != ele[25][5];
    ele[24][2] != ele[26][0];
    ele[24][2] != ele[26][1];
    ele[24][2] != ele[26][2];
    ele[24][2] != ele[26][3];
    ele[24][2] != ele[26][4];
    ele[24][2] != ele[26][5];
    ele[24][2] != ele[27][0];
    ele[24][2] != ele[27][1];
    ele[24][2] != ele[27][2];
    ele[24][2] != ele[27][3];
    ele[24][2] != ele[27][4];
    ele[24][2] != ele[27][5];
    ele[24][2] != ele[28][0];
    ele[24][2] != ele[28][1];
    ele[24][2] != ele[28][2];
    ele[24][2] != ele[28][3];
    ele[24][2] != ele[28][4];
    ele[24][2] != ele[28][5];
    ele[24][2] != ele[29][0];
    ele[24][2] != ele[29][1];
    ele[24][2] != ele[29][2];
    ele[24][2] != ele[29][3];
    ele[24][2] != ele[29][4];
    ele[24][2] != ele[29][5];
    ele[24][2] != ele[30][2];
    ele[24][2] != ele[31][2];
    ele[24][2] != ele[32][2];
    ele[24][2] != ele[33][2];
    ele[24][2] != ele[34][2];
    ele[24][2] != ele[35][2];
    ele[24][20] != ele[24][21];
    ele[24][20] != ele[24][22];
    ele[24][20] != ele[24][23];
    ele[24][20] != ele[24][24];
    ele[24][20] != ele[24][25];
    ele[24][20] != ele[24][26];
    ele[24][20] != ele[24][27];
    ele[24][20] != ele[24][28];
    ele[24][20] != ele[24][29];
    ele[24][20] != ele[24][30];
    ele[24][20] != ele[24][31];
    ele[24][20] != ele[24][32];
    ele[24][20] != ele[24][33];
    ele[24][20] != ele[24][34];
    ele[24][20] != ele[24][35];
    ele[24][20] != ele[25][18];
    ele[24][20] != ele[25][19];
    ele[24][20] != ele[25][20];
    ele[24][20] != ele[25][21];
    ele[24][20] != ele[25][22];
    ele[24][20] != ele[25][23];
    ele[24][20] != ele[26][18];
    ele[24][20] != ele[26][19];
    ele[24][20] != ele[26][20];
    ele[24][20] != ele[26][21];
    ele[24][20] != ele[26][22];
    ele[24][20] != ele[26][23];
    ele[24][20] != ele[27][18];
    ele[24][20] != ele[27][19];
    ele[24][20] != ele[27][20];
    ele[24][20] != ele[27][21];
    ele[24][20] != ele[27][22];
    ele[24][20] != ele[27][23];
    ele[24][20] != ele[28][18];
    ele[24][20] != ele[28][19];
    ele[24][20] != ele[28][20];
    ele[24][20] != ele[28][21];
    ele[24][20] != ele[28][22];
    ele[24][20] != ele[28][23];
    ele[24][20] != ele[29][18];
    ele[24][20] != ele[29][19];
    ele[24][20] != ele[29][20];
    ele[24][20] != ele[29][21];
    ele[24][20] != ele[29][22];
    ele[24][20] != ele[29][23];
    ele[24][20] != ele[30][20];
    ele[24][20] != ele[31][20];
    ele[24][20] != ele[32][20];
    ele[24][20] != ele[33][20];
    ele[24][20] != ele[34][20];
    ele[24][20] != ele[35][20];
    ele[24][21] != ele[24][22];
    ele[24][21] != ele[24][23];
    ele[24][21] != ele[24][24];
    ele[24][21] != ele[24][25];
    ele[24][21] != ele[24][26];
    ele[24][21] != ele[24][27];
    ele[24][21] != ele[24][28];
    ele[24][21] != ele[24][29];
    ele[24][21] != ele[24][30];
    ele[24][21] != ele[24][31];
    ele[24][21] != ele[24][32];
    ele[24][21] != ele[24][33];
    ele[24][21] != ele[24][34];
    ele[24][21] != ele[24][35];
    ele[24][21] != ele[25][18];
    ele[24][21] != ele[25][19];
    ele[24][21] != ele[25][20];
    ele[24][21] != ele[25][21];
    ele[24][21] != ele[25][22];
    ele[24][21] != ele[25][23];
    ele[24][21] != ele[26][18];
    ele[24][21] != ele[26][19];
    ele[24][21] != ele[26][20];
    ele[24][21] != ele[26][21];
    ele[24][21] != ele[26][22];
    ele[24][21] != ele[26][23];
    ele[24][21] != ele[27][18];
    ele[24][21] != ele[27][19];
    ele[24][21] != ele[27][20];
    ele[24][21] != ele[27][21];
    ele[24][21] != ele[27][22];
    ele[24][21] != ele[27][23];
    ele[24][21] != ele[28][18];
    ele[24][21] != ele[28][19];
    ele[24][21] != ele[28][20];
    ele[24][21] != ele[28][21];
    ele[24][21] != ele[28][22];
    ele[24][21] != ele[28][23];
    ele[24][21] != ele[29][18];
    ele[24][21] != ele[29][19];
    ele[24][21] != ele[29][20];
    ele[24][21] != ele[29][21];
    ele[24][21] != ele[29][22];
    ele[24][21] != ele[29][23];
    ele[24][21] != ele[30][21];
    ele[24][21] != ele[31][21];
    ele[24][21] != ele[32][21];
    ele[24][21] != ele[33][21];
    ele[24][21] != ele[34][21];
    ele[24][21] != ele[35][21];
    ele[24][22] != ele[24][23];
    ele[24][22] != ele[24][24];
    ele[24][22] != ele[24][25];
    ele[24][22] != ele[24][26];
    ele[24][22] != ele[24][27];
    ele[24][22] != ele[24][28];
    ele[24][22] != ele[24][29];
    ele[24][22] != ele[24][30];
    ele[24][22] != ele[24][31];
    ele[24][22] != ele[24][32];
    ele[24][22] != ele[24][33];
    ele[24][22] != ele[24][34];
    ele[24][22] != ele[24][35];
    ele[24][22] != ele[25][18];
    ele[24][22] != ele[25][19];
    ele[24][22] != ele[25][20];
    ele[24][22] != ele[25][21];
    ele[24][22] != ele[25][22];
    ele[24][22] != ele[25][23];
    ele[24][22] != ele[26][18];
    ele[24][22] != ele[26][19];
    ele[24][22] != ele[26][20];
    ele[24][22] != ele[26][21];
    ele[24][22] != ele[26][22];
    ele[24][22] != ele[26][23];
    ele[24][22] != ele[27][18];
    ele[24][22] != ele[27][19];
    ele[24][22] != ele[27][20];
    ele[24][22] != ele[27][21];
    ele[24][22] != ele[27][22];
    ele[24][22] != ele[27][23];
    ele[24][22] != ele[28][18];
    ele[24][22] != ele[28][19];
    ele[24][22] != ele[28][20];
    ele[24][22] != ele[28][21];
    ele[24][22] != ele[28][22];
    ele[24][22] != ele[28][23];
    ele[24][22] != ele[29][18];
    ele[24][22] != ele[29][19];
    ele[24][22] != ele[29][20];
    ele[24][22] != ele[29][21];
    ele[24][22] != ele[29][22];
    ele[24][22] != ele[29][23];
    ele[24][22] != ele[30][22];
    ele[24][22] != ele[31][22];
    ele[24][22] != ele[32][22];
    ele[24][22] != ele[33][22];
    ele[24][22] != ele[34][22];
    ele[24][22] != ele[35][22];
    ele[24][23] != ele[24][24];
    ele[24][23] != ele[24][25];
    ele[24][23] != ele[24][26];
    ele[24][23] != ele[24][27];
    ele[24][23] != ele[24][28];
    ele[24][23] != ele[24][29];
    ele[24][23] != ele[24][30];
    ele[24][23] != ele[24][31];
    ele[24][23] != ele[24][32];
    ele[24][23] != ele[24][33];
    ele[24][23] != ele[24][34];
    ele[24][23] != ele[24][35];
    ele[24][23] != ele[25][18];
    ele[24][23] != ele[25][19];
    ele[24][23] != ele[25][20];
    ele[24][23] != ele[25][21];
    ele[24][23] != ele[25][22];
    ele[24][23] != ele[25][23];
    ele[24][23] != ele[26][18];
    ele[24][23] != ele[26][19];
    ele[24][23] != ele[26][20];
    ele[24][23] != ele[26][21];
    ele[24][23] != ele[26][22];
    ele[24][23] != ele[26][23];
    ele[24][23] != ele[27][18];
    ele[24][23] != ele[27][19];
    ele[24][23] != ele[27][20];
    ele[24][23] != ele[27][21];
    ele[24][23] != ele[27][22];
    ele[24][23] != ele[27][23];
    ele[24][23] != ele[28][18];
    ele[24][23] != ele[28][19];
    ele[24][23] != ele[28][20];
    ele[24][23] != ele[28][21];
    ele[24][23] != ele[28][22];
    ele[24][23] != ele[28][23];
    ele[24][23] != ele[29][18];
    ele[24][23] != ele[29][19];
    ele[24][23] != ele[29][20];
    ele[24][23] != ele[29][21];
    ele[24][23] != ele[29][22];
    ele[24][23] != ele[29][23];
    ele[24][23] != ele[30][23];
    ele[24][23] != ele[31][23];
    ele[24][23] != ele[32][23];
    ele[24][23] != ele[33][23];
    ele[24][23] != ele[34][23];
    ele[24][23] != ele[35][23];
    ele[24][24] != ele[24][25];
    ele[24][24] != ele[24][26];
    ele[24][24] != ele[24][27];
    ele[24][24] != ele[24][28];
    ele[24][24] != ele[24][29];
    ele[24][24] != ele[24][30];
    ele[24][24] != ele[24][31];
    ele[24][24] != ele[24][32];
    ele[24][24] != ele[24][33];
    ele[24][24] != ele[24][34];
    ele[24][24] != ele[24][35];
    ele[24][24] != ele[25][24];
    ele[24][24] != ele[25][25];
    ele[24][24] != ele[25][26];
    ele[24][24] != ele[25][27];
    ele[24][24] != ele[25][28];
    ele[24][24] != ele[25][29];
    ele[24][24] != ele[26][24];
    ele[24][24] != ele[26][25];
    ele[24][24] != ele[26][26];
    ele[24][24] != ele[26][27];
    ele[24][24] != ele[26][28];
    ele[24][24] != ele[26][29];
    ele[24][24] != ele[27][24];
    ele[24][24] != ele[27][25];
    ele[24][24] != ele[27][26];
    ele[24][24] != ele[27][27];
    ele[24][24] != ele[27][28];
    ele[24][24] != ele[27][29];
    ele[24][24] != ele[28][24];
    ele[24][24] != ele[28][25];
    ele[24][24] != ele[28][26];
    ele[24][24] != ele[28][27];
    ele[24][24] != ele[28][28];
    ele[24][24] != ele[28][29];
    ele[24][24] != ele[29][24];
    ele[24][24] != ele[29][25];
    ele[24][24] != ele[29][26];
    ele[24][24] != ele[29][27];
    ele[24][24] != ele[29][28];
    ele[24][24] != ele[29][29];
    ele[24][24] != ele[30][24];
    ele[24][24] != ele[31][24];
    ele[24][24] != ele[32][24];
    ele[24][24] != ele[33][24];
    ele[24][24] != ele[34][24];
    ele[24][24] != ele[35][24];
    ele[24][25] != ele[24][26];
    ele[24][25] != ele[24][27];
    ele[24][25] != ele[24][28];
    ele[24][25] != ele[24][29];
    ele[24][25] != ele[24][30];
    ele[24][25] != ele[24][31];
    ele[24][25] != ele[24][32];
    ele[24][25] != ele[24][33];
    ele[24][25] != ele[24][34];
    ele[24][25] != ele[24][35];
    ele[24][25] != ele[25][24];
    ele[24][25] != ele[25][25];
    ele[24][25] != ele[25][26];
    ele[24][25] != ele[25][27];
    ele[24][25] != ele[25][28];
    ele[24][25] != ele[25][29];
    ele[24][25] != ele[26][24];
    ele[24][25] != ele[26][25];
    ele[24][25] != ele[26][26];
    ele[24][25] != ele[26][27];
    ele[24][25] != ele[26][28];
    ele[24][25] != ele[26][29];
    ele[24][25] != ele[27][24];
    ele[24][25] != ele[27][25];
    ele[24][25] != ele[27][26];
    ele[24][25] != ele[27][27];
    ele[24][25] != ele[27][28];
    ele[24][25] != ele[27][29];
    ele[24][25] != ele[28][24];
    ele[24][25] != ele[28][25];
    ele[24][25] != ele[28][26];
    ele[24][25] != ele[28][27];
    ele[24][25] != ele[28][28];
    ele[24][25] != ele[28][29];
    ele[24][25] != ele[29][24];
    ele[24][25] != ele[29][25];
    ele[24][25] != ele[29][26];
    ele[24][25] != ele[29][27];
    ele[24][25] != ele[29][28];
    ele[24][25] != ele[29][29];
    ele[24][25] != ele[30][25];
    ele[24][25] != ele[31][25];
    ele[24][25] != ele[32][25];
    ele[24][25] != ele[33][25];
    ele[24][25] != ele[34][25];
    ele[24][25] != ele[35][25];
    ele[24][26] != ele[24][27];
    ele[24][26] != ele[24][28];
    ele[24][26] != ele[24][29];
    ele[24][26] != ele[24][30];
    ele[24][26] != ele[24][31];
    ele[24][26] != ele[24][32];
    ele[24][26] != ele[24][33];
    ele[24][26] != ele[24][34];
    ele[24][26] != ele[24][35];
    ele[24][26] != ele[25][24];
    ele[24][26] != ele[25][25];
    ele[24][26] != ele[25][26];
    ele[24][26] != ele[25][27];
    ele[24][26] != ele[25][28];
    ele[24][26] != ele[25][29];
    ele[24][26] != ele[26][24];
    ele[24][26] != ele[26][25];
    ele[24][26] != ele[26][26];
    ele[24][26] != ele[26][27];
    ele[24][26] != ele[26][28];
    ele[24][26] != ele[26][29];
    ele[24][26] != ele[27][24];
    ele[24][26] != ele[27][25];
    ele[24][26] != ele[27][26];
    ele[24][26] != ele[27][27];
    ele[24][26] != ele[27][28];
    ele[24][26] != ele[27][29];
    ele[24][26] != ele[28][24];
    ele[24][26] != ele[28][25];
    ele[24][26] != ele[28][26];
    ele[24][26] != ele[28][27];
    ele[24][26] != ele[28][28];
    ele[24][26] != ele[28][29];
    ele[24][26] != ele[29][24];
    ele[24][26] != ele[29][25];
    ele[24][26] != ele[29][26];
    ele[24][26] != ele[29][27];
    ele[24][26] != ele[29][28];
    ele[24][26] != ele[29][29];
    ele[24][26] != ele[30][26];
    ele[24][26] != ele[31][26];
    ele[24][26] != ele[32][26];
    ele[24][26] != ele[33][26];
    ele[24][26] != ele[34][26];
    ele[24][26] != ele[35][26];
    ele[24][27] != ele[24][28];
    ele[24][27] != ele[24][29];
    ele[24][27] != ele[24][30];
    ele[24][27] != ele[24][31];
    ele[24][27] != ele[24][32];
    ele[24][27] != ele[24][33];
    ele[24][27] != ele[24][34];
    ele[24][27] != ele[24][35];
    ele[24][27] != ele[25][24];
    ele[24][27] != ele[25][25];
    ele[24][27] != ele[25][26];
    ele[24][27] != ele[25][27];
    ele[24][27] != ele[25][28];
    ele[24][27] != ele[25][29];
    ele[24][27] != ele[26][24];
    ele[24][27] != ele[26][25];
    ele[24][27] != ele[26][26];
    ele[24][27] != ele[26][27];
    ele[24][27] != ele[26][28];
    ele[24][27] != ele[26][29];
    ele[24][27] != ele[27][24];
    ele[24][27] != ele[27][25];
    ele[24][27] != ele[27][26];
    ele[24][27] != ele[27][27];
    ele[24][27] != ele[27][28];
    ele[24][27] != ele[27][29];
    ele[24][27] != ele[28][24];
    ele[24][27] != ele[28][25];
    ele[24][27] != ele[28][26];
    ele[24][27] != ele[28][27];
    ele[24][27] != ele[28][28];
    ele[24][27] != ele[28][29];
    ele[24][27] != ele[29][24];
    ele[24][27] != ele[29][25];
    ele[24][27] != ele[29][26];
    ele[24][27] != ele[29][27];
    ele[24][27] != ele[29][28];
    ele[24][27] != ele[29][29];
    ele[24][27] != ele[30][27];
    ele[24][27] != ele[31][27];
    ele[24][27] != ele[32][27];
    ele[24][27] != ele[33][27];
    ele[24][27] != ele[34][27];
    ele[24][27] != ele[35][27];
    ele[24][28] != ele[24][29];
    ele[24][28] != ele[24][30];
    ele[24][28] != ele[24][31];
    ele[24][28] != ele[24][32];
    ele[24][28] != ele[24][33];
    ele[24][28] != ele[24][34];
    ele[24][28] != ele[24][35];
    ele[24][28] != ele[25][24];
    ele[24][28] != ele[25][25];
    ele[24][28] != ele[25][26];
    ele[24][28] != ele[25][27];
    ele[24][28] != ele[25][28];
    ele[24][28] != ele[25][29];
    ele[24][28] != ele[26][24];
    ele[24][28] != ele[26][25];
    ele[24][28] != ele[26][26];
    ele[24][28] != ele[26][27];
    ele[24][28] != ele[26][28];
    ele[24][28] != ele[26][29];
    ele[24][28] != ele[27][24];
    ele[24][28] != ele[27][25];
    ele[24][28] != ele[27][26];
    ele[24][28] != ele[27][27];
    ele[24][28] != ele[27][28];
    ele[24][28] != ele[27][29];
    ele[24][28] != ele[28][24];
    ele[24][28] != ele[28][25];
    ele[24][28] != ele[28][26];
    ele[24][28] != ele[28][27];
    ele[24][28] != ele[28][28];
    ele[24][28] != ele[28][29];
    ele[24][28] != ele[29][24];
    ele[24][28] != ele[29][25];
    ele[24][28] != ele[29][26];
    ele[24][28] != ele[29][27];
    ele[24][28] != ele[29][28];
    ele[24][28] != ele[29][29];
    ele[24][28] != ele[30][28];
    ele[24][28] != ele[31][28];
    ele[24][28] != ele[32][28];
    ele[24][28] != ele[33][28];
    ele[24][28] != ele[34][28];
    ele[24][28] != ele[35][28];
    ele[24][29] != ele[24][30];
    ele[24][29] != ele[24][31];
    ele[24][29] != ele[24][32];
    ele[24][29] != ele[24][33];
    ele[24][29] != ele[24][34];
    ele[24][29] != ele[24][35];
    ele[24][29] != ele[25][24];
    ele[24][29] != ele[25][25];
    ele[24][29] != ele[25][26];
    ele[24][29] != ele[25][27];
    ele[24][29] != ele[25][28];
    ele[24][29] != ele[25][29];
    ele[24][29] != ele[26][24];
    ele[24][29] != ele[26][25];
    ele[24][29] != ele[26][26];
    ele[24][29] != ele[26][27];
    ele[24][29] != ele[26][28];
    ele[24][29] != ele[26][29];
    ele[24][29] != ele[27][24];
    ele[24][29] != ele[27][25];
    ele[24][29] != ele[27][26];
    ele[24][29] != ele[27][27];
    ele[24][29] != ele[27][28];
    ele[24][29] != ele[27][29];
    ele[24][29] != ele[28][24];
    ele[24][29] != ele[28][25];
    ele[24][29] != ele[28][26];
    ele[24][29] != ele[28][27];
    ele[24][29] != ele[28][28];
    ele[24][29] != ele[28][29];
    ele[24][29] != ele[29][24];
    ele[24][29] != ele[29][25];
    ele[24][29] != ele[29][26];
    ele[24][29] != ele[29][27];
    ele[24][29] != ele[29][28];
    ele[24][29] != ele[29][29];
    ele[24][29] != ele[30][29];
    ele[24][29] != ele[31][29];
    ele[24][29] != ele[32][29];
    ele[24][29] != ele[33][29];
    ele[24][29] != ele[34][29];
    ele[24][29] != ele[35][29];
    ele[24][3] != ele[24][10];
    ele[24][3] != ele[24][11];
    ele[24][3] != ele[24][12];
    ele[24][3] != ele[24][13];
    ele[24][3] != ele[24][14];
    ele[24][3] != ele[24][15];
    ele[24][3] != ele[24][16];
    ele[24][3] != ele[24][17];
    ele[24][3] != ele[24][18];
    ele[24][3] != ele[24][19];
    ele[24][3] != ele[24][20];
    ele[24][3] != ele[24][21];
    ele[24][3] != ele[24][22];
    ele[24][3] != ele[24][23];
    ele[24][3] != ele[24][24];
    ele[24][3] != ele[24][25];
    ele[24][3] != ele[24][26];
    ele[24][3] != ele[24][27];
    ele[24][3] != ele[24][28];
    ele[24][3] != ele[24][29];
    ele[24][3] != ele[24][30];
    ele[24][3] != ele[24][31];
    ele[24][3] != ele[24][32];
    ele[24][3] != ele[24][33];
    ele[24][3] != ele[24][34];
    ele[24][3] != ele[24][35];
    ele[24][3] != ele[24][4];
    ele[24][3] != ele[24][5];
    ele[24][3] != ele[24][6];
    ele[24][3] != ele[24][7];
    ele[24][3] != ele[24][8];
    ele[24][3] != ele[24][9];
    ele[24][3] != ele[25][0];
    ele[24][3] != ele[25][1];
    ele[24][3] != ele[25][2];
    ele[24][3] != ele[25][3];
    ele[24][3] != ele[25][4];
    ele[24][3] != ele[25][5];
    ele[24][3] != ele[26][0];
    ele[24][3] != ele[26][1];
    ele[24][3] != ele[26][2];
    ele[24][3] != ele[26][3];
    ele[24][3] != ele[26][4];
    ele[24][3] != ele[26][5];
    ele[24][3] != ele[27][0];
    ele[24][3] != ele[27][1];
    ele[24][3] != ele[27][2];
    ele[24][3] != ele[27][3];
    ele[24][3] != ele[27][4];
    ele[24][3] != ele[27][5];
    ele[24][3] != ele[28][0];
    ele[24][3] != ele[28][1];
    ele[24][3] != ele[28][2];
    ele[24][3] != ele[28][3];
    ele[24][3] != ele[28][4];
    ele[24][3] != ele[28][5];
    ele[24][3] != ele[29][0];
    ele[24][3] != ele[29][1];
    ele[24][3] != ele[29][2];
    ele[24][3] != ele[29][3];
    ele[24][3] != ele[29][4];
    ele[24][3] != ele[29][5];
    ele[24][3] != ele[30][3];
    ele[24][3] != ele[31][3];
    ele[24][3] != ele[32][3];
    ele[24][3] != ele[33][3];
    ele[24][3] != ele[34][3];
    ele[24][3] != ele[35][3];
    ele[24][30] != ele[24][31];
    ele[24][30] != ele[24][32];
    ele[24][30] != ele[24][33];
    ele[24][30] != ele[24][34];
    ele[24][30] != ele[24][35];
    ele[24][30] != ele[25][30];
    ele[24][30] != ele[25][31];
    ele[24][30] != ele[25][32];
    ele[24][30] != ele[25][33];
    ele[24][30] != ele[25][34];
    ele[24][30] != ele[25][35];
    ele[24][30] != ele[26][30];
    ele[24][30] != ele[26][31];
    ele[24][30] != ele[26][32];
    ele[24][30] != ele[26][33];
    ele[24][30] != ele[26][34];
    ele[24][30] != ele[26][35];
    ele[24][30] != ele[27][30];
    ele[24][30] != ele[27][31];
    ele[24][30] != ele[27][32];
    ele[24][30] != ele[27][33];
    ele[24][30] != ele[27][34];
    ele[24][30] != ele[27][35];
    ele[24][30] != ele[28][30];
    ele[24][30] != ele[28][31];
    ele[24][30] != ele[28][32];
    ele[24][30] != ele[28][33];
    ele[24][30] != ele[28][34];
    ele[24][30] != ele[28][35];
    ele[24][30] != ele[29][30];
    ele[24][30] != ele[29][31];
    ele[24][30] != ele[29][32];
    ele[24][30] != ele[29][33];
    ele[24][30] != ele[29][34];
    ele[24][30] != ele[29][35];
    ele[24][30] != ele[30][30];
    ele[24][30] != ele[31][30];
    ele[24][30] != ele[32][30];
    ele[24][30] != ele[33][30];
    ele[24][30] != ele[34][30];
    ele[24][30] != ele[35][30];
    ele[24][31] != ele[24][32];
    ele[24][31] != ele[24][33];
    ele[24][31] != ele[24][34];
    ele[24][31] != ele[24][35];
    ele[24][31] != ele[25][30];
    ele[24][31] != ele[25][31];
    ele[24][31] != ele[25][32];
    ele[24][31] != ele[25][33];
    ele[24][31] != ele[25][34];
    ele[24][31] != ele[25][35];
    ele[24][31] != ele[26][30];
    ele[24][31] != ele[26][31];
    ele[24][31] != ele[26][32];
    ele[24][31] != ele[26][33];
    ele[24][31] != ele[26][34];
    ele[24][31] != ele[26][35];
    ele[24][31] != ele[27][30];
    ele[24][31] != ele[27][31];
    ele[24][31] != ele[27][32];
    ele[24][31] != ele[27][33];
    ele[24][31] != ele[27][34];
    ele[24][31] != ele[27][35];
    ele[24][31] != ele[28][30];
    ele[24][31] != ele[28][31];
    ele[24][31] != ele[28][32];
    ele[24][31] != ele[28][33];
    ele[24][31] != ele[28][34];
    ele[24][31] != ele[28][35];
    ele[24][31] != ele[29][30];
    ele[24][31] != ele[29][31];
    ele[24][31] != ele[29][32];
    ele[24][31] != ele[29][33];
    ele[24][31] != ele[29][34];
    ele[24][31] != ele[29][35];
    ele[24][31] != ele[30][31];
    ele[24][31] != ele[31][31];
    ele[24][31] != ele[32][31];
    ele[24][31] != ele[33][31];
    ele[24][31] != ele[34][31];
    ele[24][31] != ele[35][31];
    ele[24][32] != ele[24][33];
    ele[24][32] != ele[24][34];
    ele[24][32] != ele[24][35];
    ele[24][32] != ele[25][30];
    ele[24][32] != ele[25][31];
    ele[24][32] != ele[25][32];
    ele[24][32] != ele[25][33];
    ele[24][32] != ele[25][34];
    ele[24][32] != ele[25][35];
    ele[24][32] != ele[26][30];
    ele[24][32] != ele[26][31];
    ele[24][32] != ele[26][32];
    ele[24][32] != ele[26][33];
    ele[24][32] != ele[26][34];
    ele[24][32] != ele[26][35];
    ele[24][32] != ele[27][30];
    ele[24][32] != ele[27][31];
    ele[24][32] != ele[27][32];
    ele[24][32] != ele[27][33];
    ele[24][32] != ele[27][34];
    ele[24][32] != ele[27][35];
    ele[24][32] != ele[28][30];
    ele[24][32] != ele[28][31];
    ele[24][32] != ele[28][32];
    ele[24][32] != ele[28][33];
    ele[24][32] != ele[28][34];
    ele[24][32] != ele[28][35];
    ele[24][32] != ele[29][30];
    ele[24][32] != ele[29][31];
    ele[24][32] != ele[29][32];
    ele[24][32] != ele[29][33];
    ele[24][32] != ele[29][34];
    ele[24][32] != ele[29][35];
    ele[24][32] != ele[30][32];
    ele[24][32] != ele[31][32];
    ele[24][32] != ele[32][32];
    ele[24][32] != ele[33][32];
    ele[24][32] != ele[34][32];
    ele[24][32] != ele[35][32];
    ele[24][33] != ele[24][34];
    ele[24][33] != ele[24][35];
    ele[24][33] != ele[25][30];
    ele[24][33] != ele[25][31];
    ele[24][33] != ele[25][32];
    ele[24][33] != ele[25][33];
    ele[24][33] != ele[25][34];
    ele[24][33] != ele[25][35];
    ele[24][33] != ele[26][30];
    ele[24][33] != ele[26][31];
    ele[24][33] != ele[26][32];
    ele[24][33] != ele[26][33];
    ele[24][33] != ele[26][34];
    ele[24][33] != ele[26][35];
    ele[24][33] != ele[27][30];
    ele[24][33] != ele[27][31];
    ele[24][33] != ele[27][32];
    ele[24][33] != ele[27][33];
    ele[24][33] != ele[27][34];
    ele[24][33] != ele[27][35];
    ele[24][33] != ele[28][30];
    ele[24][33] != ele[28][31];
    ele[24][33] != ele[28][32];
    ele[24][33] != ele[28][33];
    ele[24][33] != ele[28][34];
    ele[24][33] != ele[28][35];
    ele[24][33] != ele[29][30];
    ele[24][33] != ele[29][31];
    ele[24][33] != ele[29][32];
    ele[24][33] != ele[29][33];
    ele[24][33] != ele[29][34];
    ele[24][33] != ele[29][35];
    ele[24][33] != ele[30][33];
    ele[24][33] != ele[31][33];
    ele[24][33] != ele[32][33];
    ele[24][33] != ele[33][33];
    ele[24][33] != ele[34][33];
    ele[24][33] != ele[35][33];
    ele[24][34] != ele[24][35];
    ele[24][34] != ele[25][30];
    ele[24][34] != ele[25][31];
    ele[24][34] != ele[25][32];
    ele[24][34] != ele[25][33];
    ele[24][34] != ele[25][34];
    ele[24][34] != ele[25][35];
    ele[24][34] != ele[26][30];
    ele[24][34] != ele[26][31];
    ele[24][34] != ele[26][32];
    ele[24][34] != ele[26][33];
    ele[24][34] != ele[26][34];
    ele[24][34] != ele[26][35];
    ele[24][34] != ele[27][30];
    ele[24][34] != ele[27][31];
    ele[24][34] != ele[27][32];
    ele[24][34] != ele[27][33];
    ele[24][34] != ele[27][34];
    ele[24][34] != ele[27][35];
    ele[24][34] != ele[28][30];
    ele[24][34] != ele[28][31];
    ele[24][34] != ele[28][32];
    ele[24][34] != ele[28][33];
    ele[24][34] != ele[28][34];
    ele[24][34] != ele[28][35];
    ele[24][34] != ele[29][30];
    ele[24][34] != ele[29][31];
    ele[24][34] != ele[29][32];
    ele[24][34] != ele[29][33];
    ele[24][34] != ele[29][34];
    ele[24][34] != ele[29][35];
    ele[24][34] != ele[30][34];
    ele[24][34] != ele[31][34];
    ele[24][34] != ele[32][34];
    ele[24][34] != ele[33][34];
    ele[24][34] != ele[34][34];
    ele[24][34] != ele[35][34];
    ele[24][35] != ele[25][30];
    ele[24][35] != ele[25][31];
    ele[24][35] != ele[25][32];
    ele[24][35] != ele[25][33];
    ele[24][35] != ele[25][34];
    ele[24][35] != ele[25][35];
    ele[24][35] != ele[26][30];
    ele[24][35] != ele[26][31];
    ele[24][35] != ele[26][32];
    ele[24][35] != ele[26][33];
    ele[24][35] != ele[26][34];
    ele[24][35] != ele[26][35];
    ele[24][35] != ele[27][30];
    ele[24][35] != ele[27][31];
    ele[24][35] != ele[27][32];
    ele[24][35] != ele[27][33];
    ele[24][35] != ele[27][34];
    ele[24][35] != ele[27][35];
    ele[24][35] != ele[28][30];
    ele[24][35] != ele[28][31];
    ele[24][35] != ele[28][32];
    ele[24][35] != ele[28][33];
    ele[24][35] != ele[28][34];
    ele[24][35] != ele[28][35];
    ele[24][35] != ele[29][30];
    ele[24][35] != ele[29][31];
    ele[24][35] != ele[29][32];
    ele[24][35] != ele[29][33];
    ele[24][35] != ele[29][34];
    ele[24][35] != ele[29][35];
    ele[24][35] != ele[30][35];
    ele[24][35] != ele[31][35];
    ele[24][35] != ele[32][35];
    ele[24][35] != ele[33][35];
    ele[24][35] != ele[34][35];
    ele[24][35] != ele[35][35];
    ele[24][4] != ele[24][10];
    ele[24][4] != ele[24][11];
    ele[24][4] != ele[24][12];
    ele[24][4] != ele[24][13];
    ele[24][4] != ele[24][14];
    ele[24][4] != ele[24][15];
    ele[24][4] != ele[24][16];
    ele[24][4] != ele[24][17];
    ele[24][4] != ele[24][18];
    ele[24][4] != ele[24][19];
    ele[24][4] != ele[24][20];
    ele[24][4] != ele[24][21];
    ele[24][4] != ele[24][22];
    ele[24][4] != ele[24][23];
    ele[24][4] != ele[24][24];
    ele[24][4] != ele[24][25];
    ele[24][4] != ele[24][26];
    ele[24][4] != ele[24][27];
    ele[24][4] != ele[24][28];
    ele[24][4] != ele[24][29];
    ele[24][4] != ele[24][30];
    ele[24][4] != ele[24][31];
    ele[24][4] != ele[24][32];
    ele[24][4] != ele[24][33];
    ele[24][4] != ele[24][34];
    ele[24][4] != ele[24][35];
    ele[24][4] != ele[24][5];
    ele[24][4] != ele[24][6];
    ele[24][4] != ele[24][7];
    ele[24][4] != ele[24][8];
    ele[24][4] != ele[24][9];
    ele[24][4] != ele[25][0];
    ele[24][4] != ele[25][1];
    ele[24][4] != ele[25][2];
    ele[24][4] != ele[25][3];
    ele[24][4] != ele[25][4];
    ele[24][4] != ele[25][5];
    ele[24][4] != ele[26][0];
    ele[24][4] != ele[26][1];
    ele[24][4] != ele[26][2];
    ele[24][4] != ele[26][3];
    ele[24][4] != ele[26][4];
    ele[24][4] != ele[26][5];
    ele[24][4] != ele[27][0];
    ele[24][4] != ele[27][1];
    ele[24][4] != ele[27][2];
    ele[24][4] != ele[27][3];
    ele[24][4] != ele[27][4];
    ele[24][4] != ele[27][5];
    ele[24][4] != ele[28][0];
    ele[24][4] != ele[28][1];
    ele[24][4] != ele[28][2];
    ele[24][4] != ele[28][3];
    ele[24][4] != ele[28][4];
    ele[24][4] != ele[28][5];
    ele[24][4] != ele[29][0];
    ele[24][4] != ele[29][1];
    ele[24][4] != ele[29][2];
    ele[24][4] != ele[29][3];
    ele[24][4] != ele[29][4];
    ele[24][4] != ele[29][5];
    ele[24][4] != ele[30][4];
    ele[24][4] != ele[31][4];
    ele[24][4] != ele[32][4];
    ele[24][4] != ele[33][4];
    ele[24][4] != ele[34][4];
    ele[24][4] != ele[35][4];
    ele[24][5] != ele[24][10];
    ele[24][5] != ele[24][11];
    ele[24][5] != ele[24][12];
    ele[24][5] != ele[24][13];
    ele[24][5] != ele[24][14];
    ele[24][5] != ele[24][15];
    ele[24][5] != ele[24][16];
    ele[24][5] != ele[24][17];
    ele[24][5] != ele[24][18];
    ele[24][5] != ele[24][19];
    ele[24][5] != ele[24][20];
    ele[24][5] != ele[24][21];
    ele[24][5] != ele[24][22];
    ele[24][5] != ele[24][23];
    ele[24][5] != ele[24][24];
    ele[24][5] != ele[24][25];
    ele[24][5] != ele[24][26];
    ele[24][5] != ele[24][27];
    ele[24][5] != ele[24][28];
    ele[24][5] != ele[24][29];
    ele[24][5] != ele[24][30];
    ele[24][5] != ele[24][31];
    ele[24][5] != ele[24][32];
    ele[24][5] != ele[24][33];
    ele[24][5] != ele[24][34];
    ele[24][5] != ele[24][35];
    ele[24][5] != ele[24][6];
    ele[24][5] != ele[24][7];
    ele[24][5] != ele[24][8];
    ele[24][5] != ele[24][9];
    ele[24][5] != ele[25][0];
    ele[24][5] != ele[25][1];
    ele[24][5] != ele[25][2];
    ele[24][5] != ele[25][3];
    ele[24][5] != ele[25][4];
    ele[24][5] != ele[25][5];
    ele[24][5] != ele[26][0];
    ele[24][5] != ele[26][1];
    ele[24][5] != ele[26][2];
    ele[24][5] != ele[26][3];
    ele[24][5] != ele[26][4];
    ele[24][5] != ele[26][5];
    ele[24][5] != ele[27][0];
    ele[24][5] != ele[27][1];
    ele[24][5] != ele[27][2];
    ele[24][5] != ele[27][3];
    ele[24][5] != ele[27][4];
    ele[24][5] != ele[27][5];
    ele[24][5] != ele[28][0];
    ele[24][5] != ele[28][1];
    ele[24][5] != ele[28][2];
    ele[24][5] != ele[28][3];
    ele[24][5] != ele[28][4];
    ele[24][5] != ele[28][5];
    ele[24][5] != ele[29][0];
    ele[24][5] != ele[29][1];
    ele[24][5] != ele[29][2];
    ele[24][5] != ele[29][3];
    ele[24][5] != ele[29][4];
    ele[24][5] != ele[29][5];
    ele[24][5] != ele[30][5];
    ele[24][5] != ele[31][5];
    ele[24][5] != ele[32][5];
    ele[24][5] != ele[33][5];
    ele[24][5] != ele[34][5];
    ele[24][5] != ele[35][5];
    ele[24][6] != ele[24][10];
    ele[24][6] != ele[24][11];
    ele[24][6] != ele[24][12];
    ele[24][6] != ele[24][13];
    ele[24][6] != ele[24][14];
    ele[24][6] != ele[24][15];
    ele[24][6] != ele[24][16];
    ele[24][6] != ele[24][17];
    ele[24][6] != ele[24][18];
    ele[24][6] != ele[24][19];
    ele[24][6] != ele[24][20];
    ele[24][6] != ele[24][21];
    ele[24][6] != ele[24][22];
    ele[24][6] != ele[24][23];
    ele[24][6] != ele[24][24];
    ele[24][6] != ele[24][25];
    ele[24][6] != ele[24][26];
    ele[24][6] != ele[24][27];
    ele[24][6] != ele[24][28];
    ele[24][6] != ele[24][29];
    ele[24][6] != ele[24][30];
    ele[24][6] != ele[24][31];
    ele[24][6] != ele[24][32];
    ele[24][6] != ele[24][33];
    ele[24][6] != ele[24][34];
    ele[24][6] != ele[24][35];
    ele[24][6] != ele[24][7];
    ele[24][6] != ele[24][8];
    ele[24][6] != ele[24][9];
    ele[24][6] != ele[25][10];
    ele[24][6] != ele[25][11];
    ele[24][6] != ele[25][6];
    ele[24][6] != ele[25][7];
    ele[24][6] != ele[25][8];
    ele[24][6] != ele[25][9];
    ele[24][6] != ele[26][10];
    ele[24][6] != ele[26][11];
    ele[24][6] != ele[26][6];
    ele[24][6] != ele[26][7];
    ele[24][6] != ele[26][8];
    ele[24][6] != ele[26][9];
    ele[24][6] != ele[27][10];
    ele[24][6] != ele[27][11];
    ele[24][6] != ele[27][6];
    ele[24][6] != ele[27][7];
    ele[24][6] != ele[27][8];
    ele[24][6] != ele[27][9];
    ele[24][6] != ele[28][10];
    ele[24][6] != ele[28][11];
    ele[24][6] != ele[28][6];
    ele[24][6] != ele[28][7];
    ele[24][6] != ele[28][8];
    ele[24][6] != ele[28][9];
    ele[24][6] != ele[29][10];
    ele[24][6] != ele[29][11];
    ele[24][6] != ele[29][6];
    ele[24][6] != ele[29][7];
    ele[24][6] != ele[29][8];
    ele[24][6] != ele[29][9];
    ele[24][6] != ele[30][6];
    ele[24][6] != ele[31][6];
    ele[24][6] != ele[32][6];
    ele[24][6] != ele[33][6];
    ele[24][6] != ele[34][6];
    ele[24][6] != ele[35][6];
    ele[24][7] != ele[24][10];
    ele[24][7] != ele[24][11];
    ele[24][7] != ele[24][12];
    ele[24][7] != ele[24][13];
    ele[24][7] != ele[24][14];
    ele[24][7] != ele[24][15];
    ele[24][7] != ele[24][16];
    ele[24][7] != ele[24][17];
    ele[24][7] != ele[24][18];
    ele[24][7] != ele[24][19];
    ele[24][7] != ele[24][20];
    ele[24][7] != ele[24][21];
    ele[24][7] != ele[24][22];
    ele[24][7] != ele[24][23];
    ele[24][7] != ele[24][24];
    ele[24][7] != ele[24][25];
    ele[24][7] != ele[24][26];
    ele[24][7] != ele[24][27];
    ele[24][7] != ele[24][28];
    ele[24][7] != ele[24][29];
    ele[24][7] != ele[24][30];
    ele[24][7] != ele[24][31];
    ele[24][7] != ele[24][32];
    ele[24][7] != ele[24][33];
    ele[24][7] != ele[24][34];
    ele[24][7] != ele[24][35];
    ele[24][7] != ele[24][8];
    ele[24][7] != ele[24][9];
    ele[24][7] != ele[25][10];
    ele[24][7] != ele[25][11];
    ele[24][7] != ele[25][6];
    ele[24][7] != ele[25][7];
    ele[24][7] != ele[25][8];
    ele[24][7] != ele[25][9];
    ele[24][7] != ele[26][10];
    ele[24][7] != ele[26][11];
    ele[24][7] != ele[26][6];
    ele[24][7] != ele[26][7];
    ele[24][7] != ele[26][8];
    ele[24][7] != ele[26][9];
    ele[24][7] != ele[27][10];
    ele[24][7] != ele[27][11];
    ele[24][7] != ele[27][6];
    ele[24][7] != ele[27][7];
    ele[24][7] != ele[27][8];
    ele[24][7] != ele[27][9];
    ele[24][7] != ele[28][10];
    ele[24][7] != ele[28][11];
    ele[24][7] != ele[28][6];
    ele[24][7] != ele[28][7];
    ele[24][7] != ele[28][8];
    ele[24][7] != ele[28][9];
    ele[24][7] != ele[29][10];
    ele[24][7] != ele[29][11];
    ele[24][7] != ele[29][6];
    ele[24][7] != ele[29][7];
    ele[24][7] != ele[29][8];
    ele[24][7] != ele[29][9];
    ele[24][7] != ele[30][7];
    ele[24][7] != ele[31][7];
    ele[24][7] != ele[32][7];
    ele[24][7] != ele[33][7];
    ele[24][7] != ele[34][7];
    ele[24][7] != ele[35][7];
    ele[24][8] != ele[24][10];
    ele[24][8] != ele[24][11];
    ele[24][8] != ele[24][12];
    ele[24][8] != ele[24][13];
    ele[24][8] != ele[24][14];
    ele[24][8] != ele[24][15];
    ele[24][8] != ele[24][16];
    ele[24][8] != ele[24][17];
    ele[24][8] != ele[24][18];
    ele[24][8] != ele[24][19];
    ele[24][8] != ele[24][20];
    ele[24][8] != ele[24][21];
    ele[24][8] != ele[24][22];
    ele[24][8] != ele[24][23];
    ele[24][8] != ele[24][24];
    ele[24][8] != ele[24][25];
    ele[24][8] != ele[24][26];
    ele[24][8] != ele[24][27];
    ele[24][8] != ele[24][28];
    ele[24][8] != ele[24][29];
    ele[24][8] != ele[24][30];
    ele[24][8] != ele[24][31];
    ele[24][8] != ele[24][32];
    ele[24][8] != ele[24][33];
    ele[24][8] != ele[24][34];
    ele[24][8] != ele[24][35];
    ele[24][8] != ele[24][9];
    ele[24][8] != ele[25][10];
    ele[24][8] != ele[25][11];
    ele[24][8] != ele[25][6];
    ele[24][8] != ele[25][7];
    ele[24][8] != ele[25][8];
    ele[24][8] != ele[25][9];
    ele[24][8] != ele[26][10];
    ele[24][8] != ele[26][11];
    ele[24][8] != ele[26][6];
    ele[24][8] != ele[26][7];
    ele[24][8] != ele[26][8];
    ele[24][8] != ele[26][9];
    ele[24][8] != ele[27][10];
    ele[24][8] != ele[27][11];
    ele[24][8] != ele[27][6];
    ele[24][8] != ele[27][7];
    ele[24][8] != ele[27][8];
    ele[24][8] != ele[27][9];
    ele[24][8] != ele[28][10];
    ele[24][8] != ele[28][11];
    ele[24][8] != ele[28][6];
    ele[24][8] != ele[28][7];
    ele[24][8] != ele[28][8];
    ele[24][8] != ele[28][9];
    ele[24][8] != ele[29][10];
    ele[24][8] != ele[29][11];
    ele[24][8] != ele[29][6];
    ele[24][8] != ele[29][7];
    ele[24][8] != ele[29][8];
    ele[24][8] != ele[29][9];
    ele[24][8] != ele[30][8];
    ele[24][8] != ele[31][8];
    ele[24][8] != ele[32][8];
    ele[24][8] != ele[33][8];
    ele[24][8] != ele[34][8];
    ele[24][8] != ele[35][8];
    ele[24][9] != ele[24][10];
    ele[24][9] != ele[24][11];
    ele[24][9] != ele[24][12];
    ele[24][9] != ele[24][13];
    ele[24][9] != ele[24][14];
    ele[24][9] != ele[24][15];
    ele[24][9] != ele[24][16];
    ele[24][9] != ele[24][17];
    ele[24][9] != ele[24][18];
    ele[24][9] != ele[24][19];
    ele[24][9] != ele[24][20];
    ele[24][9] != ele[24][21];
    ele[24][9] != ele[24][22];
    ele[24][9] != ele[24][23];
    ele[24][9] != ele[24][24];
    ele[24][9] != ele[24][25];
    ele[24][9] != ele[24][26];
    ele[24][9] != ele[24][27];
    ele[24][9] != ele[24][28];
    ele[24][9] != ele[24][29];
    ele[24][9] != ele[24][30];
    ele[24][9] != ele[24][31];
    ele[24][9] != ele[24][32];
    ele[24][9] != ele[24][33];
    ele[24][9] != ele[24][34];
    ele[24][9] != ele[24][35];
    ele[24][9] != ele[25][10];
    ele[24][9] != ele[25][11];
    ele[24][9] != ele[25][6];
    ele[24][9] != ele[25][7];
    ele[24][9] != ele[25][8];
    ele[24][9] != ele[25][9];
    ele[24][9] != ele[26][10];
    ele[24][9] != ele[26][11];
    ele[24][9] != ele[26][6];
    ele[24][9] != ele[26][7];
    ele[24][9] != ele[26][8];
    ele[24][9] != ele[26][9];
    ele[24][9] != ele[27][10];
    ele[24][9] != ele[27][11];
    ele[24][9] != ele[27][6];
    ele[24][9] != ele[27][7];
    ele[24][9] != ele[27][8];
    ele[24][9] != ele[27][9];
    ele[24][9] != ele[28][10];
    ele[24][9] != ele[28][11];
    ele[24][9] != ele[28][6];
    ele[24][9] != ele[28][7];
    ele[24][9] != ele[28][8];
    ele[24][9] != ele[28][9];
    ele[24][9] != ele[29][10];
    ele[24][9] != ele[29][11];
    ele[24][9] != ele[29][6];
    ele[24][9] != ele[29][7];
    ele[24][9] != ele[29][8];
    ele[24][9] != ele[29][9];
    ele[24][9] != ele[30][9];
    ele[24][9] != ele[31][9];
    ele[24][9] != ele[32][9];
    ele[24][9] != ele[33][9];
    ele[24][9] != ele[34][9];
    ele[24][9] != ele[35][9];
    ele[25][0] != ele[25][1];
    ele[25][0] != ele[25][10];
    ele[25][0] != ele[25][11];
    ele[25][0] != ele[25][12];
    ele[25][0] != ele[25][13];
    ele[25][0] != ele[25][14];
    ele[25][0] != ele[25][15];
    ele[25][0] != ele[25][16];
    ele[25][0] != ele[25][17];
    ele[25][0] != ele[25][18];
    ele[25][0] != ele[25][19];
    ele[25][0] != ele[25][2];
    ele[25][0] != ele[25][20];
    ele[25][0] != ele[25][21];
    ele[25][0] != ele[25][22];
    ele[25][0] != ele[25][23];
    ele[25][0] != ele[25][24];
    ele[25][0] != ele[25][25];
    ele[25][0] != ele[25][26];
    ele[25][0] != ele[25][27];
    ele[25][0] != ele[25][28];
    ele[25][0] != ele[25][29];
    ele[25][0] != ele[25][3];
    ele[25][0] != ele[25][30];
    ele[25][0] != ele[25][31];
    ele[25][0] != ele[25][32];
    ele[25][0] != ele[25][33];
    ele[25][0] != ele[25][34];
    ele[25][0] != ele[25][35];
    ele[25][0] != ele[25][4];
    ele[25][0] != ele[25][5];
    ele[25][0] != ele[25][6];
    ele[25][0] != ele[25][7];
    ele[25][0] != ele[25][8];
    ele[25][0] != ele[25][9];
    ele[25][0] != ele[26][0];
    ele[25][0] != ele[26][1];
    ele[25][0] != ele[26][2];
    ele[25][0] != ele[26][3];
    ele[25][0] != ele[26][4];
    ele[25][0] != ele[26][5];
    ele[25][0] != ele[27][0];
    ele[25][0] != ele[27][1];
    ele[25][0] != ele[27][2];
    ele[25][0] != ele[27][3];
    ele[25][0] != ele[27][4];
    ele[25][0] != ele[27][5];
    ele[25][0] != ele[28][0];
    ele[25][0] != ele[28][1];
    ele[25][0] != ele[28][2];
    ele[25][0] != ele[28][3];
    ele[25][0] != ele[28][4];
    ele[25][0] != ele[28][5];
    ele[25][0] != ele[29][0];
    ele[25][0] != ele[29][1];
    ele[25][0] != ele[29][2];
    ele[25][0] != ele[29][3];
    ele[25][0] != ele[29][4];
    ele[25][0] != ele[29][5];
    ele[25][0] != ele[30][0];
    ele[25][0] != ele[31][0];
    ele[25][0] != ele[32][0];
    ele[25][0] != ele[33][0];
    ele[25][0] != ele[34][0];
    ele[25][0] != ele[35][0];
    ele[25][1] != ele[25][10];
    ele[25][1] != ele[25][11];
    ele[25][1] != ele[25][12];
    ele[25][1] != ele[25][13];
    ele[25][1] != ele[25][14];
    ele[25][1] != ele[25][15];
    ele[25][1] != ele[25][16];
    ele[25][1] != ele[25][17];
    ele[25][1] != ele[25][18];
    ele[25][1] != ele[25][19];
    ele[25][1] != ele[25][2];
    ele[25][1] != ele[25][20];
    ele[25][1] != ele[25][21];
    ele[25][1] != ele[25][22];
    ele[25][1] != ele[25][23];
    ele[25][1] != ele[25][24];
    ele[25][1] != ele[25][25];
    ele[25][1] != ele[25][26];
    ele[25][1] != ele[25][27];
    ele[25][1] != ele[25][28];
    ele[25][1] != ele[25][29];
    ele[25][1] != ele[25][3];
    ele[25][1] != ele[25][30];
    ele[25][1] != ele[25][31];
    ele[25][1] != ele[25][32];
    ele[25][1] != ele[25][33];
    ele[25][1] != ele[25][34];
    ele[25][1] != ele[25][35];
    ele[25][1] != ele[25][4];
    ele[25][1] != ele[25][5];
    ele[25][1] != ele[25][6];
    ele[25][1] != ele[25][7];
    ele[25][1] != ele[25][8];
    ele[25][1] != ele[25][9];
    ele[25][1] != ele[26][0];
    ele[25][1] != ele[26][1];
    ele[25][1] != ele[26][2];
    ele[25][1] != ele[26][3];
    ele[25][1] != ele[26][4];
    ele[25][1] != ele[26][5];
    ele[25][1] != ele[27][0];
    ele[25][1] != ele[27][1];
    ele[25][1] != ele[27][2];
    ele[25][1] != ele[27][3];
    ele[25][1] != ele[27][4];
    ele[25][1] != ele[27][5];
    ele[25][1] != ele[28][0];
    ele[25][1] != ele[28][1];
    ele[25][1] != ele[28][2];
    ele[25][1] != ele[28][3];
    ele[25][1] != ele[28][4];
    ele[25][1] != ele[28][5];
    ele[25][1] != ele[29][0];
    ele[25][1] != ele[29][1];
    ele[25][1] != ele[29][2];
    ele[25][1] != ele[29][3];
    ele[25][1] != ele[29][4];
    ele[25][1] != ele[29][5];
    ele[25][1] != ele[30][1];
    ele[25][1] != ele[31][1];
    ele[25][1] != ele[32][1];
    ele[25][1] != ele[33][1];
    ele[25][1] != ele[34][1];
    ele[25][1] != ele[35][1];
    ele[25][10] != ele[25][11];
    ele[25][10] != ele[25][12];
    ele[25][10] != ele[25][13];
    ele[25][10] != ele[25][14];
    ele[25][10] != ele[25][15];
    ele[25][10] != ele[25][16];
    ele[25][10] != ele[25][17];
    ele[25][10] != ele[25][18];
    ele[25][10] != ele[25][19];
    ele[25][10] != ele[25][20];
    ele[25][10] != ele[25][21];
    ele[25][10] != ele[25][22];
    ele[25][10] != ele[25][23];
    ele[25][10] != ele[25][24];
    ele[25][10] != ele[25][25];
    ele[25][10] != ele[25][26];
    ele[25][10] != ele[25][27];
    ele[25][10] != ele[25][28];
    ele[25][10] != ele[25][29];
    ele[25][10] != ele[25][30];
    ele[25][10] != ele[25][31];
    ele[25][10] != ele[25][32];
    ele[25][10] != ele[25][33];
    ele[25][10] != ele[25][34];
    ele[25][10] != ele[25][35];
    ele[25][10] != ele[26][10];
    ele[25][10] != ele[26][11];
    ele[25][10] != ele[26][6];
    ele[25][10] != ele[26][7];
    ele[25][10] != ele[26][8];
    ele[25][10] != ele[26][9];
    ele[25][10] != ele[27][10];
    ele[25][10] != ele[27][11];
    ele[25][10] != ele[27][6];
    ele[25][10] != ele[27][7];
    ele[25][10] != ele[27][8];
    ele[25][10] != ele[27][9];
    ele[25][10] != ele[28][10];
    ele[25][10] != ele[28][11];
    ele[25][10] != ele[28][6];
    ele[25][10] != ele[28][7];
    ele[25][10] != ele[28][8];
    ele[25][10] != ele[28][9];
    ele[25][10] != ele[29][10];
    ele[25][10] != ele[29][11];
    ele[25][10] != ele[29][6];
    ele[25][10] != ele[29][7];
    ele[25][10] != ele[29][8];
    ele[25][10] != ele[29][9];
    ele[25][10] != ele[30][10];
    ele[25][10] != ele[31][10];
    ele[25][10] != ele[32][10];
    ele[25][10] != ele[33][10];
    ele[25][10] != ele[34][10];
    ele[25][10] != ele[35][10];
    ele[25][11] != ele[25][12];
    ele[25][11] != ele[25][13];
    ele[25][11] != ele[25][14];
    ele[25][11] != ele[25][15];
    ele[25][11] != ele[25][16];
    ele[25][11] != ele[25][17];
    ele[25][11] != ele[25][18];
    ele[25][11] != ele[25][19];
    ele[25][11] != ele[25][20];
    ele[25][11] != ele[25][21];
    ele[25][11] != ele[25][22];
    ele[25][11] != ele[25][23];
    ele[25][11] != ele[25][24];
    ele[25][11] != ele[25][25];
    ele[25][11] != ele[25][26];
    ele[25][11] != ele[25][27];
    ele[25][11] != ele[25][28];
    ele[25][11] != ele[25][29];
    ele[25][11] != ele[25][30];
    ele[25][11] != ele[25][31];
    ele[25][11] != ele[25][32];
    ele[25][11] != ele[25][33];
    ele[25][11] != ele[25][34];
    ele[25][11] != ele[25][35];
    ele[25][11] != ele[26][10];
    ele[25][11] != ele[26][11];
    ele[25][11] != ele[26][6];
    ele[25][11] != ele[26][7];
    ele[25][11] != ele[26][8];
    ele[25][11] != ele[26][9];
    ele[25][11] != ele[27][10];
    ele[25][11] != ele[27][11];
    ele[25][11] != ele[27][6];
    ele[25][11] != ele[27][7];
    ele[25][11] != ele[27][8];
    ele[25][11] != ele[27][9];
    ele[25][11] != ele[28][10];
    ele[25][11] != ele[28][11];
    ele[25][11] != ele[28][6];
    ele[25][11] != ele[28][7];
    ele[25][11] != ele[28][8];
    ele[25][11] != ele[28][9];
    ele[25][11] != ele[29][10];
    ele[25][11] != ele[29][11];
    ele[25][11] != ele[29][6];
    ele[25][11] != ele[29][7];
    ele[25][11] != ele[29][8];
    ele[25][11] != ele[29][9];
    ele[25][11] != ele[30][11];
    ele[25][11] != ele[31][11];
    ele[25][11] != ele[32][11];
    ele[25][11] != ele[33][11];
    ele[25][11] != ele[34][11];
    ele[25][11] != ele[35][11];
    ele[25][12] != ele[25][13];
    ele[25][12] != ele[25][14];
    ele[25][12] != ele[25][15];
    ele[25][12] != ele[25][16];
    ele[25][12] != ele[25][17];
    ele[25][12] != ele[25][18];
    ele[25][12] != ele[25][19];
    ele[25][12] != ele[25][20];
    ele[25][12] != ele[25][21];
    ele[25][12] != ele[25][22];
    ele[25][12] != ele[25][23];
    ele[25][12] != ele[25][24];
    ele[25][12] != ele[25][25];
    ele[25][12] != ele[25][26];
    ele[25][12] != ele[25][27];
    ele[25][12] != ele[25][28];
    ele[25][12] != ele[25][29];
    ele[25][12] != ele[25][30];
    ele[25][12] != ele[25][31];
    ele[25][12] != ele[25][32];
    ele[25][12] != ele[25][33];
    ele[25][12] != ele[25][34];
    ele[25][12] != ele[25][35];
    ele[25][12] != ele[26][12];
    ele[25][12] != ele[26][13];
    ele[25][12] != ele[26][14];
    ele[25][12] != ele[26][15];
    ele[25][12] != ele[26][16];
    ele[25][12] != ele[26][17];
    ele[25][12] != ele[27][12];
    ele[25][12] != ele[27][13];
    ele[25][12] != ele[27][14];
    ele[25][12] != ele[27][15];
    ele[25][12] != ele[27][16];
    ele[25][12] != ele[27][17];
    ele[25][12] != ele[28][12];
    ele[25][12] != ele[28][13];
    ele[25][12] != ele[28][14];
    ele[25][12] != ele[28][15];
    ele[25][12] != ele[28][16];
    ele[25][12] != ele[28][17];
    ele[25][12] != ele[29][12];
    ele[25][12] != ele[29][13];
    ele[25][12] != ele[29][14];
    ele[25][12] != ele[29][15];
    ele[25][12] != ele[29][16];
    ele[25][12] != ele[29][17];
    ele[25][12] != ele[30][12];
    ele[25][12] != ele[31][12];
    ele[25][12] != ele[32][12];
    ele[25][12] != ele[33][12];
    ele[25][12] != ele[34][12];
    ele[25][12] != ele[35][12];
    ele[25][13] != ele[25][14];
    ele[25][13] != ele[25][15];
    ele[25][13] != ele[25][16];
    ele[25][13] != ele[25][17];
    ele[25][13] != ele[25][18];
    ele[25][13] != ele[25][19];
    ele[25][13] != ele[25][20];
    ele[25][13] != ele[25][21];
    ele[25][13] != ele[25][22];
    ele[25][13] != ele[25][23];
    ele[25][13] != ele[25][24];
    ele[25][13] != ele[25][25];
    ele[25][13] != ele[25][26];
    ele[25][13] != ele[25][27];
    ele[25][13] != ele[25][28];
    ele[25][13] != ele[25][29];
    ele[25][13] != ele[25][30];
    ele[25][13] != ele[25][31];
    ele[25][13] != ele[25][32];
    ele[25][13] != ele[25][33];
    ele[25][13] != ele[25][34];
    ele[25][13] != ele[25][35];
    ele[25][13] != ele[26][12];
    ele[25][13] != ele[26][13];
    ele[25][13] != ele[26][14];
    ele[25][13] != ele[26][15];
    ele[25][13] != ele[26][16];
    ele[25][13] != ele[26][17];
    ele[25][13] != ele[27][12];
    ele[25][13] != ele[27][13];
    ele[25][13] != ele[27][14];
    ele[25][13] != ele[27][15];
    ele[25][13] != ele[27][16];
    ele[25][13] != ele[27][17];
    ele[25][13] != ele[28][12];
    ele[25][13] != ele[28][13];
    ele[25][13] != ele[28][14];
    ele[25][13] != ele[28][15];
    ele[25][13] != ele[28][16];
    ele[25][13] != ele[28][17];
    ele[25][13] != ele[29][12];
    ele[25][13] != ele[29][13];
    ele[25][13] != ele[29][14];
    ele[25][13] != ele[29][15];
    ele[25][13] != ele[29][16];
    ele[25][13] != ele[29][17];
    ele[25][13] != ele[30][13];
    ele[25][13] != ele[31][13];
    ele[25][13] != ele[32][13];
    ele[25][13] != ele[33][13];
    ele[25][13] != ele[34][13];
    ele[25][13] != ele[35][13];
    ele[25][14] != ele[25][15];
    ele[25][14] != ele[25][16];
    ele[25][14] != ele[25][17];
    ele[25][14] != ele[25][18];
    ele[25][14] != ele[25][19];
    ele[25][14] != ele[25][20];
    ele[25][14] != ele[25][21];
    ele[25][14] != ele[25][22];
    ele[25][14] != ele[25][23];
    ele[25][14] != ele[25][24];
    ele[25][14] != ele[25][25];
    ele[25][14] != ele[25][26];
    ele[25][14] != ele[25][27];
    ele[25][14] != ele[25][28];
    ele[25][14] != ele[25][29];
    ele[25][14] != ele[25][30];
    ele[25][14] != ele[25][31];
    ele[25][14] != ele[25][32];
    ele[25][14] != ele[25][33];
    ele[25][14] != ele[25][34];
    ele[25][14] != ele[25][35];
    ele[25][14] != ele[26][12];
    ele[25][14] != ele[26][13];
    ele[25][14] != ele[26][14];
    ele[25][14] != ele[26][15];
    ele[25][14] != ele[26][16];
    ele[25][14] != ele[26][17];
    ele[25][14] != ele[27][12];
    ele[25][14] != ele[27][13];
    ele[25][14] != ele[27][14];
    ele[25][14] != ele[27][15];
    ele[25][14] != ele[27][16];
    ele[25][14] != ele[27][17];
    ele[25][14] != ele[28][12];
    ele[25][14] != ele[28][13];
    ele[25][14] != ele[28][14];
    ele[25][14] != ele[28][15];
    ele[25][14] != ele[28][16];
    ele[25][14] != ele[28][17];
    ele[25][14] != ele[29][12];
    ele[25][14] != ele[29][13];
    ele[25][14] != ele[29][14];
    ele[25][14] != ele[29][15];
    ele[25][14] != ele[29][16];
    ele[25][14] != ele[29][17];
    ele[25][14] != ele[30][14];
    ele[25][14] != ele[31][14];
    ele[25][14] != ele[32][14];
    ele[25][14] != ele[33][14];
    ele[25][14] != ele[34][14];
    ele[25][14] != ele[35][14];
    ele[25][15] != ele[25][16];
    ele[25][15] != ele[25][17];
    ele[25][15] != ele[25][18];
    ele[25][15] != ele[25][19];
    ele[25][15] != ele[25][20];
    ele[25][15] != ele[25][21];
    ele[25][15] != ele[25][22];
    ele[25][15] != ele[25][23];
    ele[25][15] != ele[25][24];
    ele[25][15] != ele[25][25];
    ele[25][15] != ele[25][26];
    ele[25][15] != ele[25][27];
    ele[25][15] != ele[25][28];
    ele[25][15] != ele[25][29];
    ele[25][15] != ele[25][30];
    ele[25][15] != ele[25][31];
    ele[25][15] != ele[25][32];
    ele[25][15] != ele[25][33];
    ele[25][15] != ele[25][34];
    ele[25][15] != ele[25][35];
    ele[25][15] != ele[26][12];
    ele[25][15] != ele[26][13];
    ele[25][15] != ele[26][14];
    ele[25][15] != ele[26][15];
    ele[25][15] != ele[26][16];
    ele[25][15] != ele[26][17];
    ele[25][15] != ele[27][12];
    ele[25][15] != ele[27][13];
    ele[25][15] != ele[27][14];
    ele[25][15] != ele[27][15];
    ele[25][15] != ele[27][16];
    ele[25][15] != ele[27][17];
    ele[25][15] != ele[28][12];
    ele[25][15] != ele[28][13];
    ele[25][15] != ele[28][14];
    ele[25][15] != ele[28][15];
    ele[25][15] != ele[28][16];
    ele[25][15] != ele[28][17];
    ele[25][15] != ele[29][12];
    ele[25][15] != ele[29][13];
    ele[25][15] != ele[29][14];
    ele[25][15] != ele[29][15];
    ele[25][15] != ele[29][16];
    ele[25][15] != ele[29][17];
    ele[25][15] != ele[30][15];
    ele[25][15] != ele[31][15];
    ele[25][15] != ele[32][15];
    ele[25][15] != ele[33][15];
    ele[25][15] != ele[34][15];
    ele[25][15] != ele[35][15];
    ele[25][16] != ele[25][17];
    ele[25][16] != ele[25][18];
    ele[25][16] != ele[25][19];
    ele[25][16] != ele[25][20];
    ele[25][16] != ele[25][21];
    ele[25][16] != ele[25][22];
    ele[25][16] != ele[25][23];
    ele[25][16] != ele[25][24];
    ele[25][16] != ele[25][25];
    ele[25][16] != ele[25][26];
    ele[25][16] != ele[25][27];
    ele[25][16] != ele[25][28];
    ele[25][16] != ele[25][29];
    ele[25][16] != ele[25][30];
    ele[25][16] != ele[25][31];
    ele[25][16] != ele[25][32];
    ele[25][16] != ele[25][33];
    ele[25][16] != ele[25][34];
    ele[25][16] != ele[25][35];
    ele[25][16] != ele[26][12];
    ele[25][16] != ele[26][13];
    ele[25][16] != ele[26][14];
    ele[25][16] != ele[26][15];
    ele[25][16] != ele[26][16];
    ele[25][16] != ele[26][17];
    ele[25][16] != ele[27][12];
    ele[25][16] != ele[27][13];
    ele[25][16] != ele[27][14];
    ele[25][16] != ele[27][15];
    ele[25][16] != ele[27][16];
    ele[25][16] != ele[27][17];
    ele[25][16] != ele[28][12];
    ele[25][16] != ele[28][13];
    ele[25][16] != ele[28][14];
    ele[25][16] != ele[28][15];
    ele[25][16] != ele[28][16];
    ele[25][16] != ele[28][17];
    ele[25][16] != ele[29][12];
    ele[25][16] != ele[29][13];
    ele[25][16] != ele[29][14];
    ele[25][16] != ele[29][15];
    ele[25][16] != ele[29][16];
    ele[25][16] != ele[29][17];
    ele[25][16] != ele[30][16];
    ele[25][16] != ele[31][16];
    ele[25][16] != ele[32][16];
    ele[25][16] != ele[33][16];
    ele[25][16] != ele[34][16];
    ele[25][16] != ele[35][16];
    ele[25][17] != ele[25][18];
    ele[25][17] != ele[25][19];
    ele[25][17] != ele[25][20];
    ele[25][17] != ele[25][21];
    ele[25][17] != ele[25][22];
    ele[25][17] != ele[25][23];
    ele[25][17] != ele[25][24];
    ele[25][17] != ele[25][25];
    ele[25][17] != ele[25][26];
    ele[25][17] != ele[25][27];
    ele[25][17] != ele[25][28];
    ele[25][17] != ele[25][29];
    ele[25][17] != ele[25][30];
    ele[25][17] != ele[25][31];
    ele[25][17] != ele[25][32];
    ele[25][17] != ele[25][33];
    ele[25][17] != ele[25][34];
    ele[25][17] != ele[25][35];
    ele[25][17] != ele[26][12];
    ele[25][17] != ele[26][13];
    ele[25][17] != ele[26][14];
    ele[25][17] != ele[26][15];
    ele[25][17] != ele[26][16];
    ele[25][17] != ele[26][17];
    ele[25][17] != ele[27][12];
    ele[25][17] != ele[27][13];
    ele[25][17] != ele[27][14];
    ele[25][17] != ele[27][15];
    ele[25][17] != ele[27][16];
    ele[25][17] != ele[27][17];
    ele[25][17] != ele[28][12];
    ele[25][17] != ele[28][13];
    ele[25][17] != ele[28][14];
    ele[25][17] != ele[28][15];
    ele[25][17] != ele[28][16];
    ele[25][17] != ele[28][17];
    ele[25][17] != ele[29][12];
    ele[25][17] != ele[29][13];
    ele[25][17] != ele[29][14];
    ele[25][17] != ele[29][15];
    ele[25][17] != ele[29][16];
    ele[25][17] != ele[29][17];
    ele[25][17] != ele[30][17];
    ele[25][17] != ele[31][17];
    ele[25][17] != ele[32][17];
    ele[25][17] != ele[33][17];
    ele[25][17] != ele[34][17];
    ele[25][17] != ele[35][17];
    ele[25][18] != ele[25][19];
    ele[25][18] != ele[25][20];
    ele[25][18] != ele[25][21];
    ele[25][18] != ele[25][22];
    ele[25][18] != ele[25][23];
    ele[25][18] != ele[25][24];
    ele[25][18] != ele[25][25];
    ele[25][18] != ele[25][26];
    ele[25][18] != ele[25][27];
    ele[25][18] != ele[25][28];
    ele[25][18] != ele[25][29];
    ele[25][18] != ele[25][30];
    ele[25][18] != ele[25][31];
    ele[25][18] != ele[25][32];
    ele[25][18] != ele[25][33];
    ele[25][18] != ele[25][34];
    ele[25][18] != ele[25][35];
    ele[25][18] != ele[26][18];
    ele[25][18] != ele[26][19];
    ele[25][18] != ele[26][20];
    ele[25][18] != ele[26][21];
    ele[25][18] != ele[26][22];
    ele[25][18] != ele[26][23];
    ele[25][18] != ele[27][18];
    ele[25][18] != ele[27][19];
    ele[25][18] != ele[27][20];
    ele[25][18] != ele[27][21];
    ele[25][18] != ele[27][22];
    ele[25][18] != ele[27][23];
    ele[25][18] != ele[28][18];
    ele[25][18] != ele[28][19];
    ele[25][18] != ele[28][20];
    ele[25][18] != ele[28][21];
    ele[25][18] != ele[28][22];
    ele[25][18] != ele[28][23];
    ele[25][18] != ele[29][18];
    ele[25][18] != ele[29][19];
    ele[25][18] != ele[29][20];
    ele[25][18] != ele[29][21];
    ele[25][18] != ele[29][22];
    ele[25][18] != ele[29][23];
    ele[25][18] != ele[30][18];
    ele[25][18] != ele[31][18];
    ele[25][18] != ele[32][18];
    ele[25][18] != ele[33][18];
    ele[25][18] != ele[34][18];
    ele[25][18] != ele[35][18];
    ele[25][19] != ele[25][20];
    ele[25][19] != ele[25][21];
    ele[25][19] != ele[25][22];
    ele[25][19] != ele[25][23];
    ele[25][19] != ele[25][24];
    ele[25][19] != ele[25][25];
    ele[25][19] != ele[25][26];
    ele[25][19] != ele[25][27];
    ele[25][19] != ele[25][28];
    ele[25][19] != ele[25][29];
    ele[25][19] != ele[25][30];
    ele[25][19] != ele[25][31];
    ele[25][19] != ele[25][32];
    ele[25][19] != ele[25][33];
    ele[25][19] != ele[25][34];
    ele[25][19] != ele[25][35];
    ele[25][19] != ele[26][18];
    ele[25][19] != ele[26][19];
    ele[25][19] != ele[26][20];
    ele[25][19] != ele[26][21];
    ele[25][19] != ele[26][22];
    ele[25][19] != ele[26][23];
    ele[25][19] != ele[27][18];
    ele[25][19] != ele[27][19];
    ele[25][19] != ele[27][20];
    ele[25][19] != ele[27][21];
    ele[25][19] != ele[27][22];
    ele[25][19] != ele[27][23];
    ele[25][19] != ele[28][18];
    ele[25][19] != ele[28][19];
    ele[25][19] != ele[28][20];
    ele[25][19] != ele[28][21];
    ele[25][19] != ele[28][22];
    ele[25][19] != ele[28][23];
    ele[25][19] != ele[29][18];
    ele[25][19] != ele[29][19];
    ele[25][19] != ele[29][20];
    ele[25][19] != ele[29][21];
    ele[25][19] != ele[29][22];
    ele[25][19] != ele[29][23];
    ele[25][19] != ele[30][19];
    ele[25][19] != ele[31][19];
    ele[25][19] != ele[32][19];
    ele[25][19] != ele[33][19];
    ele[25][19] != ele[34][19];
    ele[25][19] != ele[35][19];
    ele[25][2] != ele[25][10];
    ele[25][2] != ele[25][11];
    ele[25][2] != ele[25][12];
    ele[25][2] != ele[25][13];
    ele[25][2] != ele[25][14];
    ele[25][2] != ele[25][15];
    ele[25][2] != ele[25][16];
    ele[25][2] != ele[25][17];
    ele[25][2] != ele[25][18];
    ele[25][2] != ele[25][19];
    ele[25][2] != ele[25][20];
    ele[25][2] != ele[25][21];
    ele[25][2] != ele[25][22];
    ele[25][2] != ele[25][23];
    ele[25][2] != ele[25][24];
    ele[25][2] != ele[25][25];
    ele[25][2] != ele[25][26];
    ele[25][2] != ele[25][27];
    ele[25][2] != ele[25][28];
    ele[25][2] != ele[25][29];
    ele[25][2] != ele[25][3];
    ele[25][2] != ele[25][30];
    ele[25][2] != ele[25][31];
    ele[25][2] != ele[25][32];
    ele[25][2] != ele[25][33];
    ele[25][2] != ele[25][34];
    ele[25][2] != ele[25][35];
    ele[25][2] != ele[25][4];
    ele[25][2] != ele[25][5];
    ele[25][2] != ele[25][6];
    ele[25][2] != ele[25][7];
    ele[25][2] != ele[25][8];
    ele[25][2] != ele[25][9];
    ele[25][2] != ele[26][0];
    ele[25][2] != ele[26][1];
    ele[25][2] != ele[26][2];
    ele[25][2] != ele[26][3];
    ele[25][2] != ele[26][4];
    ele[25][2] != ele[26][5];
    ele[25][2] != ele[27][0];
    ele[25][2] != ele[27][1];
    ele[25][2] != ele[27][2];
    ele[25][2] != ele[27][3];
    ele[25][2] != ele[27][4];
    ele[25][2] != ele[27][5];
    ele[25][2] != ele[28][0];
    ele[25][2] != ele[28][1];
    ele[25][2] != ele[28][2];
    ele[25][2] != ele[28][3];
    ele[25][2] != ele[28][4];
    ele[25][2] != ele[28][5];
    ele[25][2] != ele[29][0];
    ele[25][2] != ele[29][1];
    ele[25][2] != ele[29][2];
    ele[25][2] != ele[29][3];
    ele[25][2] != ele[29][4];
    ele[25][2] != ele[29][5];
    ele[25][2] != ele[30][2];
    ele[25][2] != ele[31][2];
    ele[25][2] != ele[32][2];
    ele[25][2] != ele[33][2];
    ele[25][2] != ele[34][2];
    ele[25][2] != ele[35][2];
    ele[25][20] != ele[25][21];
    ele[25][20] != ele[25][22];
    ele[25][20] != ele[25][23];
    ele[25][20] != ele[25][24];
    ele[25][20] != ele[25][25];
    ele[25][20] != ele[25][26];
    ele[25][20] != ele[25][27];
    ele[25][20] != ele[25][28];
    ele[25][20] != ele[25][29];
    ele[25][20] != ele[25][30];
    ele[25][20] != ele[25][31];
    ele[25][20] != ele[25][32];
    ele[25][20] != ele[25][33];
    ele[25][20] != ele[25][34];
    ele[25][20] != ele[25][35];
    ele[25][20] != ele[26][18];
    ele[25][20] != ele[26][19];
    ele[25][20] != ele[26][20];
    ele[25][20] != ele[26][21];
    ele[25][20] != ele[26][22];
    ele[25][20] != ele[26][23];
    ele[25][20] != ele[27][18];
    ele[25][20] != ele[27][19];
    ele[25][20] != ele[27][20];
    ele[25][20] != ele[27][21];
    ele[25][20] != ele[27][22];
    ele[25][20] != ele[27][23];
    ele[25][20] != ele[28][18];
    ele[25][20] != ele[28][19];
    ele[25][20] != ele[28][20];
    ele[25][20] != ele[28][21];
    ele[25][20] != ele[28][22];
    ele[25][20] != ele[28][23];
    ele[25][20] != ele[29][18];
    ele[25][20] != ele[29][19];
    ele[25][20] != ele[29][20];
    ele[25][20] != ele[29][21];
    ele[25][20] != ele[29][22];
    ele[25][20] != ele[29][23];
    ele[25][20] != ele[30][20];
    ele[25][20] != ele[31][20];
    ele[25][20] != ele[32][20];
    ele[25][20] != ele[33][20];
    ele[25][20] != ele[34][20];
    ele[25][20] != ele[35][20];
    ele[25][21] != ele[25][22];
    ele[25][21] != ele[25][23];
    ele[25][21] != ele[25][24];
    ele[25][21] != ele[25][25];
    ele[25][21] != ele[25][26];
    ele[25][21] != ele[25][27];
    ele[25][21] != ele[25][28];
    ele[25][21] != ele[25][29];
    ele[25][21] != ele[25][30];
    ele[25][21] != ele[25][31];
    ele[25][21] != ele[25][32];
    ele[25][21] != ele[25][33];
    ele[25][21] != ele[25][34];
    ele[25][21] != ele[25][35];
    ele[25][21] != ele[26][18];
    ele[25][21] != ele[26][19];
    ele[25][21] != ele[26][20];
    ele[25][21] != ele[26][21];
    ele[25][21] != ele[26][22];
    ele[25][21] != ele[26][23];
    ele[25][21] != ele[27][18];
    ele[25][21] != ele[27][19];
    ele[25][21] != ele[27][20];
    ele[25][21] != ele[27][21];
    ele[25][21] != ele[27][22];
    ele[25][21] != ele[27][23];
    ele[25][21] != ele[28][18];
    ele[25][21] != ele[28][19];
    ele[25][21] != ele[28][20];
    ele[25][21] != ele[28][21];
    ele[25][21] != ele[28][22];
    ele[25][21] != ele[28][23];
    ele[25][21] != ele[29][18];
    ele[25][21] != ele[29][19];
    ele[25][21] != ele[29][20];
    ele[25][21] != ele[29][21];
    ele[25][21] != ele[29][22];
    ele[25][21] != ele[29][23];
    ele[25][21] != ele[30][21];
    ele[25][21] != ele[31][21];
    ele[25][21] != ele[32][21];
    ele[25][21] != ele[33][21];
    ele[25][21] != ele[34][21];
    ele[25][21] != ele[35][21];
    ele[25][22] != ele[25][23];
    ele[25][22] != ele[25][24];
    ele[25][22] != ele[25][25];
    ele[25][22] != ele[25][26];
    ele[25][22] != ele[25][27];
    ele[25][22] != ele[25][28];
    ele[25][22] != ele[25][29];
    ele[25][22] != ele[25][30];
    ele[25][22] != ele[25][31];
    ele[25][22] != ele[25][32];
    ele[25][22] != ele[25][33];
    ele[25][22] != ele[25][34];
    ele[25][22] != ele[25][35];
    ele[25][22] != ele[26][18];
    ele[25][22] != ele[26][19];
    ele[25][22] != ele[26][20];
    ele[25][22] != ele[26][21];
    ele[25][22] != ele[26][22];
    ele[25][22] != ele[26][23];
    ele[25][22] != ele[27][18];
    ele[25][22] != ele[27][19];
    ele[25][22] != ele[27][20];
    ele[25][22] != ele[27][21];
    ele[25][22] != ele[27][22];
    ele[25][22] != ele[27][23];
    ele[25][22] != ele[28][18];
    ele[25][22] != ele[28][19];
    ele[25][22] != ele[28][20];
    ele[25][22] != ele[28][21];
    ele[25][22] != ele[28][22];
    ele[25][22] != ele[28][23];
    ele[25][22] != ele[29][18];
    ele[25][22] != ele[29][19];
    ele[25][22] != ele[29][20];
    ele[25][22] != ele[29][21];
    ele[25][22] != ele[29][22];
    ele[25][22] != ele[29][23];
    ele[25][22] != ele[30][22];
    ele[25][22] != ele[31][22];
    ele[25][22] != ele[32][22];
    ele[25][22] != ele[33][22];
    ele[25][22] != ele[34][22];
    ele[25][22] != ele[35][22];
    ele[25][23] != ele[25][24];
    ele[25][23] != ele[25][25];
    ele[25][23] != ele[25][26];
    ele[25][23] != ele[25][27];
    ele[25][23] != ele[25][28];
    ele[25][23] != ele[25][29];
    ele[25][23] != ele[25][30];
    ele[25][23] != ele[25][31];
    ele[25][23] != ele[25][32];
    ele[25][23] != ele[25][33];
    ele[25][23] != ele[25][34];
    ele[25][23] != ele[25][35];
    ele[25][23] != ele[26][18];
    ele[25][23] != ele[26][19];
    ele[25][23] != ele[26][20];
    ele[25][23] != ele[26][21];
    ele[25][23] != ele[26][22];
    ele[25][23] != ele[26][23];
    ele[25][23] != ele[27][18];
    ele[25][23] != ele[27][19];
    ele[25][23] != ele[27][20];
    ele[25][23] != ele[27][21];
    ele[25][23] != ele[27][22];
    ele[25][23] != ele[27][23];
    ele[25][23] != ele[28][18];
    ele[25][23] != ele[28][19];
    ele[25][23] != ele[28][20];
    ele[25][23] != ele[28][21];
    ele[25][23] != ele[28][22];
    ele[25][23] != ele[28][23];
    ele[25][23] != ele[29][18];
    ele[25][23] != ele[29][19];
    ele[25][23] != ele[29][20];
    ele[25][23] != ele[29][21];
    ele[25][23] != ele[29][22];
    ele[25][23] != ele[29][23];
    ele[25][23] != ele[30][23];
    ele[25][23] != ele[31][23];
    ele[25][23] != ele[32][23];
    ele[25][23] != ele[33][23];
    ele[25][23] != ele[34][23];
    ele[25][23] != ele[35][23];
    ele[25][24] != ele[25][25];
    ele[25][24] != ele[25][26];
    ele[25][24] != ele[25][27];
    ele[25][24] != ele[25][28];
    ele[25][24] != ele[25][29];
    ele[25][24] != ele[25][30];
    ele[25][24] != ele[25][31];
    ele[25][24] != ele[25][32];
    ele[25][24] != ele[25][33];
    ele[25][24] != ele[25][34];
    ele[25][24] != ele[25][35];
    ele[25][24] != ele[26][24];
    ele[25][24] != ele[26][25];
    ele[25][24] != ele[26][26];
    ele[25][24] != ele[26][27];
    ele[25][24] != ele[26][28];
    ele[25][24] != ele[26][29];
    ele[25][24] != ele[27][24];
    ele[25][24] != ele[27][25];
    ele[25][24] != ele[27][26];
    ele[25][24] != ele[27][27];
    ele[25][24] != ele[27][28];
    ele[25][24] != ele[27][29];
    ele[25][24] != ele[28][24];
    ele[25][24] != ele[28][25];
    ele[25][24] != ele[28][26];
    ele[25][24] != ele[28][27];
    ele[25][24] != ele[28][28];
    ele[25][24] != ele[28][29];
    ele[25][24] != ele[29][24];
    ele[25][24] != ele[29][25];
    ele[25][24] != ele[29][26];
    ele[25][24] != ele[29][27];
    ele[25][24] != ele[29][28];
    ele[25][24] != ele[29][29];
    ele[25][24] != ele[30][24];
    ele[25][24] != ele[31][24];
    ele[25][24] != ele[32][24];
    ele[25][24] != ele[33][24];
    ele[25][24] != ele[34][24];
    ele[25][24] != ele[35][24];
    ele[25][25] != ele[25][26];
    ele[25][25] != ele[25][27];
    ele[25][25] != ele[25][28];
    ele[25][25] != ele[25][29];
    ele[25][25] != ele[25][30];
    ele[25][25] != ele[25][31];
    ele[25][25] != ele[25][32];
    ele[25][25] != ele[25][33];
    ele[25][25] != ele[25][34];
    ele[25][25] != ele[25][35];
    ele[25][25] != ele[26][24];
    ele[25][25] != ele[26][25];
    ele[25][25] != ele[26][26];
    ele[25][25] != ele[26][27];
    ele[25][25] != ele[26][28];
    ele[25][25] != ele[26][29];
    ele[25][25] != ele[27][24];
    ele[25][25] != ele[27][25];
    ele[25][25] != ele[27][26];
    ele[25][25] != ele[27][27];
    ele[25][25] != ele[27][28];
    ele[25][25] != ele[27][29];
    ele[25][25] != ele[28][24];
    ele[25][25] != ele[28][25];
    ele[25][25] != ele[28][26];
    ele[25][25] != ele[28][27];
    ele[25][25] != ele[28][28];
    ele[25][25] != ele[28][29];
    ele[25][25] != ele[29][24];
    ele[25][25] != ele[29][25];
    ele[25][25] != ele[29][26];
    ele[25][25] != ele[29][27];
    ele[25][25] != ele[29][28];
    ele[25][25] != ele[29][29];
    ele[25][25] != ele[30][25];
    ele[25][25] != ele[31][25];
    ele[25][25] != ele[32][25];
    ele[25][25] != ele[33][25];
    ele[25][25] != ele[34][25];
    ele[25][25] != ele[35][25];
    ele[25][26] != ele[25][27];
    ele[25][26] != ele[25][28];
    ele[25][26] != ele[25][29];
    ele[25][26] != ele[25][30];
    ele[25][26] != ele[25][31];
    ele[25][26] != ele[25][32];
    ele[25][26] != ele[25][33];
    ele[25][26] != ele[25][34];
    ele[25][26] != ele[25][35];
    ele[25][26] != ele[26][24];
    ele[25][26] != ele[26][25];
    ele[25][26] != ele[26][26];
    ele[25][26] != ele[26][27];
    ele[25][26] != ele[26][28];
    ele[25][26] != ele[26][29];
    ele[25][26] != ele[27][24];
    ele[25][26] != ele[27][25];
    ele[25][26] != ele[27][26];
    ele[25][26] != ele[27][27];
    ele[25][26] != ele[27][28];
    ele[25][26] != ele[27][29];
    ele[25][26] != ele[28][24];
    ele[25][26] != ele[28][25];
    ele[25][26] != ele[28][26];
    ele[25][26] != ele[28][27];
    ele[25][26] != ele[28][28];
    ele[25][26] != ele[28][29];
    ele[25][26] != ele[29][24];
    ele[25][26] != ele[29][25];
    ele[25][26] != ele[29][26];
    ele[25][26] != ele[29][27];
    ele[25][26] != ele[29][28];
    ele[25][26] != ele[29][29];
    ele[25][26] != ele[30][26];
    ele[25][26] != ele[31][26];
    ele[25][26] != ele[32][26];
    ele[25][26] != ele[33][26];
    ele[25][26] != ele[34][26];
    ele[25][26] != ele[35][26];
    ele[25][27] != ele[25][28];
    ele[25][27] != ele[25][29];
    ele[25][27] != ele[25][30];
    ele[25][27] != ele[25][31];
    ele[25][27] != ele[25][32];
    ele[25][27] != ele[25][33];
    ele[25][27] != ele[25][34];
    ele[25][27] != ele[25][35];
    ele[25][27] != ele[26][24];
    ele[25][27] != ele[26][25];
    ele[25][27] != ele[26][26];
    ele[25][27] != ele[26][27];
    ele[25][27] != ele[26][28];
    ele[25][27] != ele[26][29];
    ele[25][27] != ele[27][24];
    ele[25][27] != ele[27][25];
    ele[25][27] != ele[27][26];
    ele[25][27] != ele[27][27];
    ele[25][27] != ele[27][28];
    ele[25][27] != ele[27][29];
    ele[25][27] != ele[28][24];
    ele[25][27] != ele[28][25];
    ele[25][27] != ele[28][26];
    ele[25][27] != ele[28][27];
    ele[25][27] != ele[28][28];
    ele[25][27] != ele[28][29];
    ele[25][27] != ele[29][24];
    ele[25][27] != ele[29][25];
    ele[25][27] != ele[29][26];
    ele[25][27] != ele[29][27];
    ele[25][27] != ele[29][28];
    ele[25][27] != ele[29][29];
    ele[25][27] != ele[30][27];
    ele[25][27] != ele[31][27];
    ele[25][27] != ele[32][27];
    ele[25][27] != ele[33][27];
    ele[25][27] != ele[34][27];
    ele[25][27] != ele[35][27];
    ele[25][28] != ele[25][29];
    ele[25][28] != ele[25][30];
    ele[25][28] != ele[25][31];
    ele[25][28] != ele[25][32];
    ele[25][28] != ele[25][33];
    ele[25][28] != ele[25][34];
    ele[25][28] != ele[25][35];
    ele[25][28] != ele[26][24];
    ele[25][28] != ele[26][25];
    ele[25][28] != ele[26][26];
    ele[25][28] != ele[26][27];
    ele[25][28] != ele[26][28];
    ele[25][28] != ele[26][29];
    ele[25][28] != ele[27][24];
    ele[25][28] != ele[27][25];
    ele[25][28] != ele[27][26];
    ele[25][28] != ele[27][27];
    ele[25][28] != ele[27][28];
    ele[25][28] != ele[27][29];
    ele[25][28] != ele[28][24];
    ele[25][28] != ele[28][25];
    ele[25][28] != ele[28][26];
    ele[25][28] != ele[28][27];
    ele[25][28] != ele[28][28];
    ele[25][28] != ele[28][29];
    ele[25][28] != ele[29][24];
    ele[25][28] != ele[29][25];
    ele[25][28] != ele[29][26];
    ele[25][28] != ele[29][27];
    ele[25][28] != ele[29][28];
    ele[25][28] != ele[29][29];
    ele[25][28] != ele[30][28];
    ele[25][28] != ele[31][28];
    ele[25][28] != ele[32][28];
    ele[25][28] != ele[33][28];
    ele[25][28] != ele[34][28];
    ele[25][28] != ele[35][28];
    ele[25][29] != ele[25][30];
    ele[25][29] != ele[25][31];
    ele[25][29] != ele[25][32];
    ele[25][29] != ele[25][33];
    ele[25][29] != ele[25][34];
    ele[25][29] != ele[25][35];
    ele[25][29] != ele[26][24];
    ele[25][29] != ele[26][25];
    ele[25][29] != ele[26][26];
    ele[25][29] != ele[26][27];
    ele[25][29] != ele[26][28];
    ele[25][29] != ele[26][29];
    ele[25][29] != ele[27][24];
    ele[25][29] != ele[27][25];
    ele[25][29] != ele[27][26];
    ele[25][29] != ele[27][27];
    ele[25][29] != ele[27][28];
    ele[25][29] != ele[27][29];
    ele[25][29] != ele[28][24];
    ele[25][29] != ele[28][25];
    ele[25][29] != ele[28][26];
    ele[25][29] != ele[28][27];
    ele[25][29] != ele[28][28];
    ele[25][29] != ele[28][29];
    ele[25][29] != ele[29][24];
    ele[25][29] != ele[29][25];
    ele[25][29] != ele[29][26];
    ele[25][29] != ele[29][27];
    ele[25][29] != ele[29][28];
    ele[25][29] != ele[29][29];
    ele[25][29] != ele[30][29];
    ele[25][29] != ele[31][29];
    ele[25][29] != ele[32][29];
    ele[25][29] != ele[33][29];
    ele[25][29] != ele[34][29];
    ele[25][29] != ele[35][29];
    ele[25][3] != ele[25][10];
    ele[25][3] != ele[25][11];
    ele[25][3] != ele[25][12];
    ele[25][3] != ele[25][13];
    ele[25][3] != ele[25][14];
    ele[25][3] != ele[25][15];
    ele[25][3] != ele[25][16];
    ele[25][3] != ele[25][17];
    ele[25][3] != ele[25][18];
    ele[25][3] != ele[25][19];
    ele[25][3] != ele[25][20];
    ele[25][3] != ele[25][21];
    ele[25][3] != ele[25][22];
    ele[25][3] != ele[25][23];
    ele[25][3] != ele[25][24];
    ele[25][3] != ele[25][25];
    ele[25][3] != ele[25][26];
    ele[25][3] != ele[25][27];
    ele[25][3] != ele[25][28];
    ele[25][3] != ele[25][29];
    ele[25][3] != ele[25][30];
    ele[25][3] != ele[25][31];
    ele[25][3] != ele[25][32];
    ele[25][3] != ele[25][33];
    ele[25][3] != ele[25][34];
    ele[25][3] != ele[25][35];
    ele[25][3] != ele[25][4];
    ele[25][3] != ele[25][5];
    ele[25][3] != ele[25][6];
    ele[25][3] != ele[25][7];
    ele[25][3] != ele[25][8];
    ele[25][3] != ele[25][9];
    ele[25][3] != ele[26][0];
    ele[25][3] != ele[26][1];
    ele[25][3] != ele[26][2];
    ele[25][3] != ele[26][3];
    ele[25][3] != ele[26][4];
    ele[25][3] != ele[26][5];
    ele[25][3] != ele[27][0];
    ele[25][3] != ele[27][1];
    ele[25][3] != ele[27][2];
    ele[25][3] != ele[27][3];
    ele[25][3] != ele[27][4];
    ele[25][3] != ele[27][5];
    ele[25][3] != ele[28][0];
    ele[25][3] != ele[28][1];
    ele[25][3] != ele[28][2];
    ele[25][3] != ele[28][3];
    ele[25][3] != ele[28][4];
    ele[25][3] != ele[28][5];
    ele[25][3] != ele[29][0];
    ele[25][3] != ele[29][1];
    ele[25][3] != ele[29][2];
    ele[25][3] != ele[29][3];
    ele[25][3] != ele[29][4];
    ele[25][3] != ele[29][5];
    ele[25][3] != ele[30][3];
    ele[25][3] != ele[31][3];
    ele[25][3] != ele[32][3];
    ele[25][3] != ele[33][3];
    ele[25][3] != ele[34][3];
    ele[25][3] != ele[35][3];
    ele[25][30] != ele[25][31];
    ele[25][30] != ele[25][32];
    ele[25][30] != ele[25][33];
    ele[25][30] != ele[25][34];
    ele[25][30] != ele[25][35];
    ele[25][30] != ele[26][30];
    ele[25][30] != ele[26][31];
    ele[25][30] != ele[26][32];
    ele[25][30] != ele[26][33];
    ele[25][30] != ele[26][34];
    ele[25][30] != ele[26][35];
    ele[25][30] != ele[27][30];
    ele[25][30] != ele[27][31];
    ele[25][30] != ele[27][32];
    ele[25][30] != ele[27][33];
    ele[25][30] != ele[27][34];
    ele[25][30] != ele[27][35];
    ele[25][30] != ele[28][30];
    ele[25][30] != ele[28][31];
    ele[25][30] != ele[28][32];
    ele[25][30] != ele[28][33];
    ele[25][30] != ele[28][34];
    ele[25][30] != ele[28][35];
    ele[25][30] != ele[29][30];
    ele[25][30] != ele[29][31];
    ele[25][30] != ele[29][32];
    ele[25][30] != ele[29][33];
    ele[25][30] != ele[29][34];
    ele[25][30] != ele[29][35];
    ele[25][30] != ele[30][30];
    ele[25][30] != ele[31][30];
    ele[25][30] != ele[32][30];
    ele[25][30] != ele[33][30];
    ele[25][30] != ele[34][30];
    ele[25][30] != ele[35][30];
    ele[25][31] != ele[25][32];
    ele[25][31] != ele[25][33];
    ele[25][31] != ele[25][34];
    ele[25][31] != ele[25][35];
    ele[25][31] != ele[26][30];
    ele[25][31] != ele[26][31];
    ele[25][31] != ele[26][32];
    ele[25][31] != ele[26][33];
    ele[25][31] != ele[26][34];
    ele[25][31] != ele[26][35];
    ele[25][31] != ele[27][30];
    ele[25][31] != ele[27][31];
    ele[25][31] != ele[27][32];
    ele[25][31] != ele[27][33];
    ele[25][31] != ele[27][34];
    ele[25][31] != ele[27][35];
    ele[25][31] != ele[28][30];
    ele[25][31] != ele[28][31];
    ele[25][31] != ele[28][32];
    ele[25][31] != ele[28][33];
    ele[25][31] != ele[28][34];
    ele[25][31] != ele[28][35];
    ele[25][31] != ele[29][30];
    ele[25][31] != ele[29][31];
    ele[25][31] != ele[29][32];
    ele[25][31] != ele[29][33];
    ele[25][31] != ele[29][34];
    ele[25][31] != ele[29][35];
    ele[25][31] != ele[30][31];
    ele[25][31] != ele[31][31];
    ele[25][31] != ele[32][31];
    ele[25][31] != ele[33][31];
    ele[25][31] != ele[34][31];
    ele[25][31] != ele[35][31];
    ele[25][32] != ele[25][33];
    ele[25][32] != ele[25][34];
    ele[25][32] != ele[25][35];
    ele[25][32] != ele[26][30];
    ele[25][32] != ele[26][31];
    ele[25][32] != ele[26][32];
    ele[25][32] != ele[26][33];
    ele[25][32] != ele[26][34];
    ele[25][32] != ele[26][35];
    ele[25][32] != ele[27][30];
    ele[25][32] != ele[27][31];
    ele[25][32] != ele[27][32];
    ele[25][32] != ele[27][33];
    ele[25][32] != ele[27][34];
    ele[25][32] != ele[27][35];
    ele[25][32] != ele[28][30];
    ele[25][32] != ele[28][31];
    ele[25][32] != ele[28][32];
    ele[25][32] != ele[28][33];
    ele[25][32] != ele[28][34];
    ele[25][32] != ele[28][35];
    ele[25][32] != ele[29][30];
    ele[25][32] != ele[29][31];
    ele[25][32] != ele[29][32];
    ele[25][32] != ele[29][33];
    ele[25][32] != ele[29][34];
    ele[25][32] != ele[29][35];
    ele[25][32] != ele[30][32];
    ele[25][32] != ele[31][32];
    ele[25][32] != ele[32][32];
    ele[25][32] != ele[33][32];
    ele[25][32] != ele[34][32];
    ele[25][32] != ele[35][32];
    ele[25][33] != ele[25][34];
    ele[25][33] != ele[25][35];
    ele[25][33] != ele[26][30];
    ele[25][33] != ele[26][31];
    ele[25][33] != ele[26][32];
    ele[25][33] != ele[26][33];
    ele[25][33] != ele[26][34];
    ele[25][33] != ele[26][35];
    ele[25][33] != ele[27][30];
    ele[25][33] != ele[27][31];
    ele[25][33] != ele[27][32];
    ele[25][33] != ele[27][33];
    ele[25][33] != ele[27][34];
    ele[25][33] != ele[27][35];
    ele[25][33] != ele[28][30];
    ele[25][33] != ele[28][31];
    ele[25][33] != ele[28][32];
    ele[25][33] != ele[28][33];
    ele[25][33] != ele[28][34];
    ele[25][33] != ele[28][35];
    ele[25][33] != ele[29][30];
    ele[25][33] != ele[29][31];
    ele[25][33] != ele[29][32];
    ele[25][33] != ele[29][33];
    ele[25][33] != ele[29][34];
    ele[25][33] != ele[29][35];
    ele[25][33] != ele[30][33];
    ele[25][33] != ele[31][33];
    ele[25][33] != ele[32][33];
    ele[25][33] != ele[33][33];
    ele[25][33] != ele[34][33];
    ele[25][33] != ele[35][33];
    ele[25][34] != ele[25][35];
    ele[25][34] != ele[26][30];
    ele[25][34] != ele[26][31];
    ele[25][34] != ele[26][32];
    ele[25][34] != ele[26][33];
    ele[25][34] != ele[26][34];
    ele[25][34] != ele[26][35];
    ele[25][34] != ele[27][30];
    ele[25][34] != ele[27][31];
    ele[25][34] != ele[27][32];
    ele[25][34] != ele[27][33];
    ele[25][34] != ele[27][34];
    ele[25][34] != ele[27][35];
    ele[25][34] != ele[28][30];
    ele[25][34] != ele[28][31];
    ele[25][34] != ele[28][32];
    ele[25][34] != ele[28][33];
    ele[25][34] != ele[28][34];
    ele[25][34] != ele[28][35];
    ele[25][34] != ele[29][30];
    ele[25][34] != ele[29][31];
    ele[25][34] != ele[29][32];
    ele[25][34] != ele[29][33];
    ele[25][34] != ele[29][34];
    ele[25][34] != ele[29][35];
    ele[25][34] != ele[30][34];
    ele[25][34] != ele[31][34];
    ele[25][34] != ele[32][34];
    ele[25][34] != ele[33][34];
    ele[25][34] != ele[34][34];
    ele[25][34] != ele[35][34];
    ele[25][35] != ele[26][30];
    ele[25][35] != ele[26][31];
    ele[25][35] != ele[26][32];
    ele[25][35] != ele[26][33];
    ele[25][35] != ele[26][34];
    ele[25][35] != ele[26][35];
    ele[25][35] != ele[27][30];
    ele[25][35] != ele[27][31];
    ele[25][35] != ele[27][32];
    ele[25][35] != ele[27][33];
    ele[25][35] != ele[27][34];
    ele[25][35] != ele[27][35];
    ele[25][35] != ele[28][30];
    ele[25][35] != ele[28][31];
    ele[25][35] != ele[28][32];
    ele[25][35] != ele[28][33];
    ele[25][35] != ele[28][34];
    ele[25][35] != ele[28][35];
    ele[25][35] != ele[29][30];
    ele[25][35] != ele[29][31];
    ele[25][35] != ele[29][32];
    ele[25][35] != ele[29][33];
    ele[25][35] != ele[29][34];
    ele[25][35] != ele[29][35];
    ele[25][35] != ele[30][35];
    ele[25][35] != ele[31][35];
    ele[25][35] != ele[32][35];
    ele[25][35] != ele[33][35];
    ele[25][35] != ele[34][35];
    ele[25][35] != ele[35][35];
    ele[25][4] != ele[25][10];
    ele[25][4] != ele[25][11];
    ele[25][4] != ele[25][12];
    ele[25][4] != ele[25][13];
    ele[25][4] != ele[25][14];
    ele[25][4] != ele[25][15];
    ele[25][4] != ele[25][16];
    ele[25][4] != ele[25][17];
    ele[25][4] != ele[25][18];
    ele[25][4] != ele[25][19];
    ele[25][4] != ele[25][20];
    ele[25][4] != ele[25][21];
    ele[25][4] != ele[25][22];
    ele[25][4] != ele[25][23];
    ele[25][4] != ele[25][24];
    ele[25][4] != ele[25][25];
    ele[25][4] != ele[25][26];
    ele[25][4] != ele[25][27];
    ele[25][4] != ele[25][28];
    ele[25][4] != ele[25][29];
    ele[25][4] != ele[25][30];
    ele[25][4] != ele[25][31];
    ele[25][4] != ele[25][32];
    ele[25][4] != ele[25][33];
    ele[25][4] != ele[25][34];
    ele[25][4] != ele[25][35];
    ele[25][4] != ele[25][5];
    ele[25][4] != ele[25][6];
    ele[25][4] != ele[25][7];
    ele[25][4] != ele[25][8];
    ele[25][4] != ele[25][9];
    ele[25][4] != ele[26][0];
    ele[25][4] != ele[26][1];
    ele[25][4] != ele[26][2];
    ele[25][4] != ele[26][3];
    ele[25][4] != ele[26][4];
    ele[25][4] != ele[26][5];
    ele[25][4] != ele[27][0];
    ele[25][4] != ele[27][1];
    ele[25][4] != ele[27][2];
    ele[25][4] != ele[27][3];
    ele[25][4] != ele[27][4];
    ele[25][4] != ele[27][5];
    ele[25][4] != ele[28][0];
    ele[25][4] != ele[28][1];
    ele[25][4] != ele[28][2];
    ele[25][4] != ele[28][3];
    ele[25][4] != ele[28][4];
    ele[25][4] != ele[28][5];
    ele[25][4] != ele[29][0];
    ele[25][4] != ele[29][1];
    ele[25][4] != ele[29][2];
    ele[25][4] != ele[29][3];
    ele[25][4] != ele[29][4];
    ele[25][4] != ele[29][5];
    ele[25][4] != ele[30][4];
    ele[25][4] != ele[31][4];
    ele[25][4] != ele[32][4];
    ele[25][4] != ele[33][4];
    ele[25][4] != ele[34][4];
    ele[25][4] != ele[35][4];
    ele[25][5] != ele[25][10];
    ele[25][5] != ele[25][11];
    ele[25][5] != ele[25][12];
    ele[25][5] != ele[25][13];
    ele[25][5] != ele[25][14];
    ele[25][5] != ele[25][15];
    ele[25][5] != ele[25][16];
    ele[25][5] != ele[25][17];
    ele[25][5] != ele[25][18];
    ele[25][5] != ele[25][19];
    ele[25][5] != ele[25][20];
    ele[25][5] != ele[25][21];
    ele[25][5] != ele[25][22];
    ele[25][5] != ele[25][23];
    ele[25][5] != ele[25][24];
    ele[25][5] != ele[25][25];
    ele[25][5] != ele[25][26];
    ele[25][5] != ele[25][27];
    ele[25][5] != ele[25][28];
    ele[25][5] != ele[25][29];
    ele[25][5] != ele[25][30];
    ele[25][5] != ele[25][31];
    ele[25][5] != ele[25][32];
    ele[25][5] != ele[25][33];
    ele[25][5] != ele[25][34];
    ele[25][5] != ele[25][35];
    ele[25][5] != ele[25][6];
    ele[25][5] != ele[25][7];
    ele[25][5] != ele[25][8];
    ele[25][5] != ele[25][9];
    ele[25][5] != ele[26][0];
    ele[25][5] != ele[26][1];
    ele[25][5] != ele[26][2];
    ele[25][5] != ele[26][3];
    ele[25][5] != ele[26][4];
    ele[25][5] != ele[26][5];
    ele[25][5] != ele[27][0];
    ele[25][5] != ele[27][1];
    ele[25][5] != ele[27][2];
    ele[25][5] != ele[27][3];
    ele[25][5] != ele[27][4];
    ele[25][5] != ele[27][5];
    ele[25][5] != ele[28][0];
    ele[25][5] != ele[28][1];
    ele[25][5] != ele[28][2];
    ele[25][5] != ele[28][3];
    ele[25][5] != ele[28][4];
    ele[25][5] != ele[28][5];
    ele[25][5] != ele[29][0];
    ele[25][5] != ele[29][1];
    ele[25][5] != ele[29][2];
    ele[25][5] != ele[29][3];
    ele[25][5] != ele[29][4];
    ele[25][5] != ele[29][5];
    ele[25][5] != ele[30][5];
    ele[25][5] != ele[31][5];
    ele[25][5] != ele[32][5];
    ele[25][5] != ele[33][5];
    ele[25][5] != ele[34][5];
    ele[25][5] != ele[35][5];
    ele[25][6] != ele[25][10];
    ele[25][6] != ele[25][11];
    ele[25][6] != ele[25][12];
    ele[25][6] != ele[25][13];
    ele[25][6] != ele[25][14];
    ele[25][6] != ele[25][15];
    ele[25][6] != ele[25][16];
    ele[25][6] != ele[25][17];
    ele[25][6] != ele[25][18];
    ele[25][6] != ele[25][19];
    ele[25][6] != ele[25][20];
    ele[25][6] != ele[25][21];
    ele[25][6] != ele[25][22];
    ele[25][6] != ele[25][23];
    ele[25][6] != ele[25][24];
    ele[25][6] != ele[25][25];
    ele[25][6] != ele[25][26];
    ele[25][6] != ele[25][27];
    ele[25][6] != ele[25][28];
    ele[25][6] != ele[25][29];
    ele[25][6] != ele[25][30];
    ele[25][6] != ele[25][31];
    ele[25][6] != ele[25][32];
    ele[25][6] != ele[25][33];
    ele[25][6] != ele[25][34];
    ele[25][6] != ele[25][35];
    ele[25][6] != ele[25][7];
    ele[25][6] != ele[25][8];
    ele[25][6] != ele[25][9];
    ele[25][6] != ele[26][10];
    ele[25][6] != ele[26][11];
    ele[25][6] != ele[26][6];
    ele[25][6] != ele[26][7];
    ele[25][6] != ele[26][8];
    ele[25][6] != ele[26][9];
    ele[25][6] != ele[27][10];
    ele[25][6] != ele[27][11];
    ele[25][6] != ele[27][6];
    ele[25][6] != ele[27][7];
    ele[25][6] != ele[27][8];
    ele[25][6] != ele[27][9];
    ele[25][6] != ele[28][10];
    ele[25][6] != ele[28][11];
    ele[25][6] != ele[28][6];
    ele[25][6] != ele[28][7];
    ele[25][6] != ele[28][8];
    ele[25][6] != ele[28][9];
    ele[25][6] != ele[29][10];
    ele[25][6] != ele[29][11];
    ele[25][6] != ele[29][6];
    ele[25][6] != ele[29][7];
    ele[25][6] != ele[29][8];
    ele[25][6] != ele[29][9];
    ele[25][6] != ele[30][6];
    ele[25][6] != ele[31][6];
    ele[25][6] != ele[32][6];
    ele[25][6] != ele[33][6];
    ele[25][6] != ele[34][6];
    ele[25][6] != ele[35][6];
    ele[25][7] != ele[25][10];
    ele[25][7] != ele[25][11];
    ele[25][7] != ele[25][12];
    ele[25][7] != ele[25][13];
    ele[25][7] != ele[25][14];
    ele[25][7] != ele[25][15];
    ele[25][7] != ele[25][16];
    ele[25][7] != ele[25][17];
    ele[25][7] != ele[25][18];
    ele[25][7] != ele[25][19];
    ele[25][7] != ele[25][20];
    ele[25][7] != ele[25][21];
    ele[25][7] != ele[25][22];
    ele[25][7] != ele[25][23];
    ele[25][7] != ele[25][24];
    ele[25][7] != ele[25][25];
    ele[25][7] != ele[25][26];
    ele[25][7] != ele[25][27];
    ele[25][7] != ele[25][28];
    ele[25][7] != ele[25][29];
    ele[25][7] != ele[25][30];
    ele[25][7] != ele[25][31];
    ele[25][7] != ele[25][32];
    ele[25][7] != ele[25][33];
    ele[25][7] != ele[25][34];
    ele[25][7] != ele[25][35];
    ele[25][7] != ele[25][8];
    ele[25][7] != ele[25][9];
    ele[25][7] != ele[26][10];
    ele[25][7] != ele[26][11];
    ele[25][7] != ele[26][6];
    ele[25][7] != ele[26][7];
    ele[25][7] != ele[26][8];
    ele[25][7] != ele[26][9];
    ele[25][7] != ele[27][10];
    ele[25][7] != ele[27][11];
    ele[25][7] != ele[27][6];
    ele[25][7] != ele[27][7];
    ele[25][7] != ele[27][8];
    ele[25][7] != ele[27][9];
    ele[25][7] != ele[28][10];
    ele[25][7] != ele[28][11];
    ele[25][7] != ele[28][6];
    ele[25][7] != ele[28][7];
    ele[25][7] != ele[28][8];
    ele[25][7] != ele[28][9];
    ele[25][7] != ele[29][10];
    ele[25][7] != ele[29][11];
    ele[25][7] != ele[29][6];
    ele[25][7] != ele[29][7];
    ele[25][7] != ele[29][8];
    ele[25][7] != ele[29][9];
    ele[25][7] != ele[30][7];
    ele[25][7] != ele[31][7];
    ele[25][7] != ele[32][7];
    ele[25][7] != ele[33][7];
    ele[25][7] != ele[34][7];
    ele[25][7] != ele[35][7];
    ele[25][8] != ele[25][10];
    ele[25][8] != ele[25][11];
    ele[25][8] != ele[25][12];
    ele[25][8] != ele[25][13];
    ele[25][8] != ele[25][14];
    ele[25][8] != ele[25][15];
    ele[25][8] != ele[25][16];
    ele[25][8] != ele[25][17];
    ele[25][8] != ele[25][18];
    ele[25][8] != ele[25][19];
    ele[25][8] != ele[25][20];
    ele[25][8] != ele[25][21];
    ele[25][8] != ele[25][22];
    ele[25][8] != ele[25][23];
    ele[25][8] != ele[25][24];
    ele[25][8] != ele[25][25];
    ele[25][8] != ele[25][26];
    ele[25][8] != ele[25][27];
    ele[25][8] != ele[25][28];
    ele[25][8] != ele[25][29];
    ele[25][8] != ele[25][30];
    ele[25][8] != ele[25][31];
    ele[25][8] != ele[25][32];
    ele[25][8] != ele[25][33];
    ele[25][8] != ele[25][34];
    ele[25][8] != ele[25][35];
    ele[25][8] != ele[25][9];
    ele[25][8] != ele[26][10];
    ele[25][8] != ele[26][11];
    ele[25][8] != ele[26][6];
    ele[25][8] != ele[26][7];
    ele[25][8] != ele[26][8];
    ele[25][8] != ele[26][9];
    ele[25][8] != ele[27][10];
    ele[25][8] != ele[27][11];
    ele[25][8] != ele[27][6];
    ele[25][8] != ele[27][7];
    ele[25][8] != ele[27][8];
    ele[25][8] != ele[27][9];
    ele[25][8] != ele[28][10];
    ele[25][8] != ele[28][11];
    ele[25][8] != ele[28][6];
    ele[25][8] != ele[28][7];
    ele[25][8] != ele[28][8];
    ele[25][8] != ele[28][9];
    ele[25][8] != ele[29][10];
    ele[25][8] != ele[29][11];
    ele[25][8] != ele[29][6];
    ele[25][8] != ele[29][7];
    ele[25][8] != ele[29][8];
    ele[25][8] != ele[29][9];
    ele[25][8] != ele[30][8];
    ele[25][8] != ele[31][8];
    ele[25][8] != ele[32][8];
    ele[25][8] != ele[33][8];
    ele[25][8] != ele[34][8];
    ele[25][8] != ele[35][8];
    ele[25][9] != ele[25][10];
    ele[25][9] != ele[25][11];
    ele[25][9] != ele[25][12];
    ele[25][9] != ele[25][13];
    ele[25][9] != ele[25][14];
    ele[25][9] != ele[25][15];
    ele[25][9] != ele[25][16];
    ele[25][9] != ele[25][17];
    ele[25][9] != ele[25][18];
    ele[25][9] != ele[25][19];
    ele[25][9] != ele[25][20];
    ele[25][9] != ele[25][21];
    ele[25][9] != ele[25][22];
    ele[25][9] != ele[25][23];
    ele[25][9] != ele[25][24];
    ele[25][9] != ele[25][25];
    ele[25][9] != ele[25][26];
    ele[25][9] != ele[25][27];
    ele[25][9] != ele[25][28];
    ele[25][9] != ele[25][29];
    ele[25][9] != ele[25][30];
    ele[25][9] != ele[25][31];
    ele[25][9] != ele[25][32];
    ele[25][9] != ele[25][33];
    ele[25][9] != ele[25][34];
    ele[25][9] != ele[25][35];
    ele[25][9] != ele[26][10];
    ele[25][9] != ele[26][11];
    ele[25][9] != ele[26][6];
    ele[25][9] != ele[26][7];
    ele[25][9] != ele[26][8];
    ele[25][9] != ele[26][9];
    ele[25][9] != ele[27][10];
    ele[25][9] != ele[27][11];
    ele[25][9] != ele[27][6];
    ele[25][9] != ele[27][7];
    ele[25][9] != ele[27][8];
    ele[25][9] != ele[27][9];
    ele[25][9] != ele[28][10];
    ele[25][9] != ele[28][11];
    ele[25][9] != ele[28][6];
    ele[25][9] != ele[28][7];
    ele[25][9] != ele[28][8];
    ele[25][9] != ele[28][9];
    ele[25][9] != ele[29][10];
    ele[25][9] != ele[29][11];
    ele[25][9] != ele[29][6];
    ele[25][9] != ele[29][7];
    ele[25][9] != ele[29][8];
    ele[25][9] != ele[29][9];
    ele[25][9] != ele[30][9];
    ele[25][9] != ele[31][9];
    ele[25][9] != ele[32][9];
    ele[25][9] != ele[33][9];
    ele[25][9] != ele[34][9];
    ele[25][9] != ele[35][9];
    ele[26][0] != ele[26][1];
    ele[26][0] != ele[26][10];
    ele[26][0] != ele[26][11];
    ele[26][0] != ele[26][12];
    ele[26][0] != ele[26][13];
    ele[26][0] != ele[26][14];
    ele[26][0] != ele[26][15];
    ele[26][0] != ele[26][16];
    ele[26][0] != ele[26][17];
    ele[26][0] != ele[26][18];
    ele[26][0] != ele[26][19];
    ele[26][0] != ele[26][2];
    ele[26][0] != ele[26][20];
    ele[26][0] != ele[26][21];
    ele[26][0] != ele[26][22];
    ele[26][0] != ele[26][23];
    ele[26][0] != ele[26][24];
    ele[26][0] != ele[26][25];
    ele[26][0] != ele[26][26];
    ele[26][0] != ele[26][27];
    ele[26][0] != ele[26][28];
    ele[26][0] != ele[26][29];
    ele[26][0] != ele[26][3];
    ele[26][0] != ele[26][30];
    ele[26][0] != ele[26][31];
    ele[26][0] != ele[26][32];
    ele[26][0] != ele[26][33];
    ele[26][0] != ele[26][34];
    ele[26][0] != ele[26][35];
    ele[26][0] != ele[26][4];
    ele[26][0] != ele[26][5];
    ele[26][0] != ele[26][6];
    ele[26][0] != ele[26][7];
    ele[26][0] != ele[26][8];
    ele[26][0] != ele[26][9];
    ele[26][0] != ele[27][0];
    ele[26][0] != ele[27][1];
    ele[26][0] != ele[27][2];
    ele[26][0] != ele[27][3];
    ele[26][0] != ele[27][4];
    ele[26][0] != ele[27][5];
    ele[26][0] != ele[28][0];
    ele[26][0] != ele[28][1];
    ele[26][0] != ele[28][2];
    ele[26][0] != ele[28][3];
    ele[26][0] != ele[28][4];
    ele[26][0] != ele[28][5];
    ele[26][0] != ele[29][0];
    ele[26][0] != ele[29][1];
    ele[26][0] != ele[29][2];
    ele[26][0] != ele[29][3];
    ele[26][0] != ele[29][4];
    ele[26][0] != ele[29][5];
    ele[26][0] != ele[30][0];
    ele[26][0] != ele[31][0];
    ele[26][0] != ele[32][0];
    ele[26][0] != ele[33][0];
    ele[26][0] != ele[34][0];
    ele[26][0] != ele[35][0];
    ele[26][1] != ele[26][10];
    ele[26][1] != ele[26][11];
    ele[26][1] != ele[26][12];
    ele[26][1] != ele[26][13];
    ele[26][1] != ele[26][14];
    ele[26][1] != ele[26][15];
    ele[26][1] != ele[26][16];
    ele[26][1] != ele[26][17];
    ele[26][1] != ele[26][18];
    ele[26][1] != ele[26][19];
    ele[26][1] != ele[26][2];
    ele[26][1] != ele[26][20];
    ele[26][1] != ele[26][21];
    ele[26][1] != ele[26][22];
    ele[26][1] != ele[26][23];
    ele[26][1] != ele[26][24];
    ele[26][1] != ele[26][25];
    ele[26][1] != ele[26][26];
    ele[26][1] != ele[26][27];
    ele[26][1] != ele[26][28];
    ele[26][1] != ele[26][29];
    ele[26][1] != ele[26][3];
    ele[26][1] != ele[26][30];
    ele[26][1] != ele[26][31];
    ele[26][1] != ele[26][32];
    ele[26][1] != ele[26][33];
    ele[26][1] != ele[26][34];
    ele[26][1] != ele[26][35];
    ele[26][1] != ele[26][4];
    ele[26][1] != ele[26][5];
    ele[26][1] != ele[26][6];
    ele[26][1] != ele[26][7];
    ele[26][1] != ele[26][8];
    ele[26][1] != ele[26][9];
    ele[26][1] != ele[27][0];
    ele[26][1] != ele[27][1];
    ele[26][1] != ele[27][2];
    ele[26][1] != ele[27][3];
    ele[26][1] != ele[27][4];
    ele[26][1] != ele[27][5];
    ele[26][1] != ele[28][0];
    ele[26][1] != ele[28][1];
    ele[26][1] != ele[28][2];
    ele[26][1] != ele[28][3];
    ele[26][1] != ele[28][4];
    ele[26][1] != ele[28][5];
    ele[26][1] != ele[29][0];
    ele[26][1] != ele[29][1];
    ele[26][1] != ele[29][2];
    ele[26][1] != ele[29][3];
    ele[26][1] != ele[29][4];
    ele[26][1] != ele[29][5];
    ele[26][1] != ele[30][1];
    ele[26][1] != ele[31][1];
    ele[26][1] != ele[32][1];
    ele[26][1] != ele[33][1];
    ele[26][1] != ele[34][1];
    ele[26][1] != ele[35][1];
    ele[26][10] != ele[26][11];
    ele[26][10] != ele[26][12];
    ele[26][10] != ele[26][13];
    ele[26][10] != ele[26][14];
    ele[26][10] != ele[26][15];
    ele[26][10] != ele[26][16];
    ele[26][10] != ele[26][17];
    ele[26][10] != ele[26][18];
    ele[26][10] != ele[26][19];
    ele[26][10] != ele[26][20];
    ele[26][10] != ele[26][21];
    ele[26][10] != ele[26][22];
    ele[26][10] != ele[26][23];
    ele[26][10] != ele[26][24];
    ele[26][10] != ele[26][25];
    ele[26][10] != ele[26][26];
    ele[26][10] != ele[26][27];
    ele[26][10] != ele[26][28];
    ele[26][10] != ele[26][29];
    ele[26][10] != ele[26][30];
    ele[26][10] != ele[26][31];
    ele[26][10] != ele[26][32];
    ele[26][10] != ele[26][33];
    ele[26][10] != ele[26][34];
    ele[26][10] != ele[26][35];
    ele[26][10] != ele[27][10];
    ele[26][10] != ele[27][11];
    ele[26][10] != ele[27][6];
    ele[26][10] != ele[27][7];
    ele[26][10] != ele[27][8];
    ele[26][10] != ele[27][9];
    ele[26][10] != ele[28][10];
    ele[26][10] != ele[28][11];
    ele[26][10] != ele[28][6];
    ele[26][10] != ele[28][7];
    ele[26][10] != ele[28][8];
    ele[26][10] != ele[28][9];
    ele[26][10] != ele[29][10];
    ele[26][10] != ele[29][11];
    ele[26][10] != ele[29][6];
    ele[26][10] != ele[29][7];
    ele[26][10] != ele[29][8];
    ele[26][10] != ele[29][9];
    ele[26][10] != ele[30][10];
    ele[26][10] != ele[31][10];
    ele[26][10] != ele[32][10];
    ele[26][10] != ele[33][10];
    ele[26][10] != ele[34][10];
    ele[26][10] != ele[35][10];
    ele[26][11] != ele[26][12];
    ele[26][11] != ele[26][13];
    ele[26][11] != ele[26][14];
    ele[26][11] != ele[26][15];
    ele[26][11] != ele[26][16];
    ele[26][11] != ele[26][17];
    ele[26][11] != ele[26][18];
    ele[26][11] != ele[26][19];
    ele[26][11] != ele[26][20];
    ele[26][11] != ele[26][21];
    ele[26][11] != ele[26][22];
    ele[26][11] != ele[26][23];
    ele[26][11] != ele[26][24];
    ele[26][11] != ele[26][25];
    ele[26][11] != ele[26][26];
    ele[26][11] != ele[26][27];
    ele[26][11] != ele[26][28];
    ele[26][11] != ele[26][29];
    ele[26][11] != ele[26][30];
    ele[26][11] != ele[26][31];
    ele[26][11] != ele[26][32];
    ele[26][11] != ele[26][33];
    ele[26][11] != ele[26][34];
    ele[26][11] != ele[26][35];
    ele[26][11] != ele[27][10];
    ele[26][11] != ele[27][11];
    ele[26][11] != ele[27][6];
    ele[26][11] != ele[27][7];
    ele[26][11] != ele[27][8];
    ele[26][11] != ele[27][9];
    ele[26][11] != ele[28][10];
    ele[26][11] != ele[28][11];
    ele[26][11] != ele[28][6];
    ele[26][11] != ele[28][7];
    ele[26][11] != ele[28][8];
    ele[26][11] != ele[28][9];
    ele[26][11] != ele[29][10];
    ele[26][11] != ele[29][11];
    ele[26][11] != ele[29][6];
    ele[26][11] != ele[29][7];
    ele[26][11] != ele[29][8];
    ele[26][11] != ele[29][9];
    ele[26][11] != ele[30][11];
    ele[26][11] != ele[31][11];
    ele[26][11] != ele[32][11];
    ele[26][11] != ele[33][11];
    ele[26][11] != ele[34][11];
    ele[26][11] != ele[35][11];
    ele[26][12] != ele[26][13];
    ele[26][12] != ele[26][14];
    ele[26][12] != ele[26][15];
    ele[26][12] != ele[26][16];
    ele[26][12] != ele[26][17];
    ele[26][12] != ele[26][18];
    ele[26][12] != ele[26][19];
    ele[26][12] != ele[26][20];
    ele[26][12] != ele[26][21];
    ele[26][12] != ele[26][22];
    ele[26][12] != ele[26][23];
    ele[26][12] != ele[26][24];
    ele[26][12] != ele[26][25];
    ele[26][12] != ele[26][26];
    ele[26][12] != ele[26][27];
    ele[26][12] != ele[26][28];
    ele[26][12] != ele[26][29];
    ele[26][12] != ele[26][30];
    ele[26][12] != ele[26][31];
    ele[26][12] != ele[26][32];
    ele[26][12] != ele[26][33];
    ele[26][12] != ele[26][34];
    ele[26][12] != ele[26][35];
    ele[26][12] != ele[27][12];
    ele[26][12] != ele[27][13];
    ele[26][12] != ele[27][14];
    ele[26][12] != ele[27][15];
    ele[26][12] != ele[27][16];
    ele[26][12] != ele[27][17];
    ele[26][12] != ele[28][12];
    ele[26][12] != ele[28][13];
    ele[26][12] != ele[28][14];
    ele[26][12] != ele[28][15];
    ele[26][12] != ele[28][16];
    ele[26][12] != ele[28][17];
    ele[26][12] != ele[29][12];
    ele[26][12] != ele[29][13];
    ele[26][12] != ele[29][14];
    ele[26][12] != ele[29][15];
    ele[26][12] != ele[29][16];
    ele[26][12] != ele[29][17];
    ele[26][12] != ele[30][12];
    ele[26][12] != ele[31][12];
    ele[26][12] != ele[32][12];
    ele[26][12] != ele[33][12];
    ele[26][12] != ele[34][12];
    ele[26][12] != ele[35][12];
    ele[26][13] != ele[26][14];
    ele[26][13] != ele[26][15];
    ele[26][13] != ele[26][16];
    ele[26][13] != ele[26][17];
    ele[26][13] != ele[26][18];
    ele[26][13] != ele[26][19];
    ele[26][13] != ele[26][20];
    ele[26][13] != ele[26][21];
    ele[26][13] != ele[26][22];
    ele[26][13] != ele[26][23];
    ele[26][13] != ele[26][24];
    ele[26][13] != ele[26][25];
    ele[26][13] != ele[26][26];
    ele[26][13] != ele[26][27];
    ele[26][13] != ele[26][28];
    ele[26][13] != ele[26][29];
    ele[26][13] != ele[26][30];
    ele[26][13] != ele[26][31];
    ele[26][13] != ele[26][32];
    ele[26][13] != ele[26][33];
    ele[26][13] != ele[26][34];
    ele[26][13] != ele[26][35];
    ele[26][13] != ele[27][12];
    ele[26][13] != ele[27][13];
    ele[26][13] != ele[27][14];
    ele[26][13] != ele[27][15];
    ele[26][13] != ele[27][16];
    ele[26][13] != ele[27][17];
    ele[26][13] != ele[28][12];
    ele[26][13] != ele[28][13];
    ele[26][13] != ele[28][14];
    ele[26][13] != ele[28][15];
    ele[26][13] != ele[28][16];
    ele[26][13] != ele[28][17];
    ele[26][13] != ele[29][12];
    ele[26][13] != ele[29][13];
    ele[26][13] != ele[29][14];
    ele[26][13] != ele[29][15];
    ele[26][13] != ele[29][16];
    ele[26][13] != ele[29][17];
    ele[26][13] != ele[30][13];
    ele[26][13] != ele[31][13];
    ele[26][13] != ele[32][13];
    ele[26][13] != ele[33][13];
    ele[26][13] != ele[34][13];
    ele[26][13] != ele[35][13];
    ele[26][14] != ele[26][15];
    ele[26][14] != ele[26][16];
    ele[26][14] != ele[26][17];
    ele[26][14] != ele[26][18];
    ele[26][14] != ele[26][19];
    ele[26][14] != ele[26][20];
    ele[26][14] != ele[26][21];
    ele[26][14] != ele[26][22];
    ele[26][14] != ele[26][23];
    ele[26][14] != ele[26][24];
    ele[26][14] != ele[26][25];
    ele[26][14] != ele[26][26];
    ele[26][14] != ele[26][27];
    ele[26][14] != ele[26][28];
    ele[26][14] != ele[26][29];
    ele[26][14] != ele[26][30];
    ele[26][14] != ele[26][31];
    ele[26][14] != ele[26][32];
    ele[26][14] != ele[26][33];
    ele[26][14] != ele[26][34];
    ele[26][14] != ele[26][35];
    ele[26][14] != ele[27][12];
    ele[26][14] != ele[27][13];
    ele[26][14] != ele[27][14];
    ele[26][14] != ele[27][15];
    ele[26][14] != ele[27][16];
    ele[26][14] != ele[27][17];
    ele[26][14] != ele[28][12];
    ele[26][14] != ele[28][13];
    ele[26][14] != ele[28][14];
    ele[26][14] != ele[28][15];
    ele[26][14] != ele[28][16];
    ele[26][14] != ele[28][17];
    ele[26][14] != ele[29][12];
    ele[26][14] != ele[29][13];
    ele[26][14] != ele[29][14];
    ele[26][14] != ele[29][15];
    ele[26][14] != ele[29][16];
    ele[26][14] != ele[29][17];
    ele[26][14] != ele[30][14];
    ele[26][14] != ele[31][14];
    ele[26][14] != ele[32][14];
    ele[26][14] != ele[33][14];
    ele[26][14] != ele[34][14];
    ele[26][14] != ele[35][14];
    ele[26][15] != ele[26][16];
    ele[26][15] != ele[26][17];
    ele[26][15] != ele[26][18];
    ele[26][15] != ele[26][19];
    ele[26][15] != ele[26][20];
    ele[26][15] != ele[26][21];
    ele[26][15] != ele[26][22];
    ele[26][15] != ele[26][23];
    ele[26][15] != ele[26][24];
    ele[26][15] != ele[26][25];
    ele[26][15] != ele[26][26];
    ele[26][15] != ele[26][27];
    ele[26][15] != ele[26][28];
    ele[26][15] != ele[26][29];
    ele[26][15] != ele[26][30];
    ele[26][15] != ele[26][31];
    ele[26][15] != ele[26][32];
    ele[26][15] != ele[26][33];
    ele[26][15] != ele[26][34];
    ele[26][15] != ele[26][35];
    ele[26][15] != ele[27][12];
    ele[26][15] != ele[27][13];
    ele[26][15] != ele[27][14];
    ele[26][15] != ele[27][15];
    ele[26][15] != ele[27][16];
    ele[26][15] != ele[27][17];
    ele[26][15] != ele[28][12];
    ele[26][15] != ele[28][13];
    ele[26][15] != ele[28][14];
    ele[26][15] != ele[28][15];
    ele[26][15] != ele[28][16];
    ele[26][15] != ele[28][17];
    ele[26][15] != ele[29][12];
    ele[26][15] != ele[29][13];
    ele[26][15] != ele[29][14];
    ele[26][15] != ele[29][15];
    ele[26][15] != ele[29][16];
    ele[26][15] != ele[29][17];
    ele[26][15] != ele[30][15];
    ele[26][15] != ele[31][15];
    ele[26][15] != ele[32][15];
    ele[26][15] != ele[33][15];
    ele[26][15] != ele[34][15];
    ele[26][15] != ele[35][15];
    ele[26][16] != ele[26][17];
    ele[26][16] != ele[26][18];
    ele[26][16] != ele[26][19];
    ele[26][16] != ele[26][20];
    ele[26][16] != ele[26][21];
    ele[26][16] != ele[26][22];
    ele[26][16] != ele[26][23];
    ele[26][16] != ele[26][24];
    ele[26][16] != ele[26][25];
    ele[26][16] != ele[26][26];
    ele[26][16] != ele[26][27];
    ele[26][16] != ele[26][28];
    ele[26][16] != ele[26][29];
    ele[26][16] != ele[26][30];
    ele[26][16] != ele[26][31];
    ele[26][16] != ele[26][32];
    ele[26][16] != ele[26][33];
    ele[26][16] != ele[26][34];
    ele[26][16] != ele[26][35];
    ele[26][16] != ele[27][12];
    ele[26][16] != ele[27][13];
    ele[26][16] != ele[27][14];
    ele[26][16] != ele[27][15];
    ele[26][16] != ele[27][16];
    ele[26][16] != ele[27][17];
    ele[26][16] != ele[28][12];
    ele[26][16] != ele[28][13];
    ele[26][16] != ele[28][14];
    ele[26][16] != ele[28][15];
    ele[26][16] != ele[28][16];
    ele[26][16] != ele[28][17];
    ele[26][16] != ele[29][12];
    ele[26][16] != ele[29][13];
    ele[26][16] != ele[29][14];
    ele[26][16] != ele[29][15];
    ele[26][16] != ele[29][16];
    ele[26][16] != ele[29][17];
    ele[26][16] != ele[30][16];
    ele[26][16] != ele[31][16];
    ele[26][16] != ele[32][16];
    ele[26][16] != ele[33][16];
    ele[26][16] != ele[34][16];
    ele[26][16] != ele[35][16];
    ele[26][17] != ele[26][18];
    ele[26][17] != ele[26][19];
    ele[26][17] != ele[26][20];
    ele[26][17] != ele[26][21];
    ele[26][17] != ele[26][22];
    ele[26][17] != ele[26][23];
    ele[26][17] != ele[26][24];
    ele[26][17] != ele[26][25];
    ele[26][17] != ele[26][26];
    ele[26][17] != ele[26][27];
    ele[26][17] != ele[26][28];
    ele[26][17] != ele[26][29];
    ele[26][17] != ele[26][30];
    ele[26][17] != ele[26][31];
    ele[26][17] != ele[26][32];
    ele[26][17] != ele[26][33];
    ele[26][17] != ele[26][34];
    ele[26][17] != ele[26][35];
    ele[26][17] != ele[27][12];
    ele[26][17] != ele[27][13];
    ele[26][17] != ele[27][14];
    ele[26][17] != ele[27][15];
    ele[26][17] != ele[27][16];
    ele[26][17] != ele[27][17];
    ele[26][17] != ele[28][12];
    ele[26][17] != ele[28][13];
    ele[26][17] != ele[28][14];
    ele[26][17] != ele[28][15];
    ele[26][17] != ele[28][16];
    ele[26][17] != ele[28][17];
    ele[26][17] != ele[29][12];
    ele[26][17] != ele[29][13];
    ele[26][17] != ele[29][14];
    ele[26][17] != ele[29][15];
    ele[26][17] != ele[29][16];
    ele[26][17] != ele[29][17];
    ele[26][17] != ele[30][17];
    ele[26][17] != ele[31][17];
    ele[26][17] != ele[32][17];
    ele[26][17] != ele[33][17];
    ele[26][17] != ele[34][17];
    ele[26][17] != ele[35][17];
    ele[26][18] != ele[26][19];
    ele[26][18] != ele[26][20];
    ele[26][18] != ele[26][21];
    ele[26][18] != ele[26][22];
    ele[26][18] != ele[26][23];
    ele[26][18] != ele[26][24];
    ele[26][18] != ele[26][25];
    ele[26][18] != ele[26][26];
    ele[26][18] != ele[26][27];
    ele[26][18] != ele[26][28];
    ele[26][18] != ele[26][29];
    ele[26][18] != ele[26][30];
    ele[26][18] != ele[26][31];
    ele[26][18] != ele[26][32];
    ele[26][18] != ele[26][33];
    ele[26][18] != ele[26][34];
    ele[26][18] != ele[26][35];
    ele[26][18] != ele[27][18];
    ele[26][18] != ele[27][19];
    ele[26][18] != ele[27][20];
    ele[26][18] != ele[27][21];
    ele[26][18] != ele[27][22];
    ele[26][18] != ele[27][23];
    ele[26][18] != ele[28][18];
    ele[26][18] != ele[28][19];
    ele[26][18] != ele[28][20];
    ele[26][18] != ele[28][21];
    ele[26][18] != ele[28][22];
    ele[26][18] != ele[28][23];
    ele[26][18] != ele[29][18];
    ele[26][18] != ele[29][19];
    ele[26][18] != ele[29][20];
    ele[26][18] != ele[29][21];
    ele[26][18] != ele[29][22];
    ele[26][18] != ele[29][23];
    ele[26][18] != ele[30][18];
    ele[26][18] != ele[31][18];
    ele[26][18] != ele[32][18];
    ele[26][18] != ele[33][18];
    ele[26][18] != ele[34][18];
    ele[26][18] != ele[35][18];
    ele[26][19] != ele[26][20];
    ele[26][19] != ele[26][21];
    ele[26][19] != ele[26][22];
    ele[26][19] != ele[26][23];
    ele[26][19] != ele[26][24];
    ele[26][19] != ele[26][25];
    ele[26][19] != ele[26][26];
    ele[26][19] != ele[26][27];
    ele[26][19] != ele[26][28];
    ele[26][19] != ele[26][29];
    ele[26][19] != ele[26][30];
    ele[26][19] != ele[26][31];
    ele[26][19] != ele[26][32];
    ele[26][19] != ele[26][33];
    ele[26][19] != ele[26][34];
    ele[26][19] != ele[26][35];
    ele[26][19] != ele[27][18];
    ele[26][19] != ele[27][19];
    ele[26][19] != ele[27][20];
    ele[26][19] != ele[27][21];
    ele[26][19] != ele[27][22];
    ele[26][19] != ele[27][23];
    ele[26][19] != ele[28][18];
    ele[26][19] != ele[28][19];
    ele[26][19] != ele[28][20];
    ele[26][19] != ele[28][21];
    ele[26][19] != ele[28][22];
    ele[26][19] != ele[28][23];
    ele[26][19] != ele[29][18];
    ele[26][19] != ele[29][19];
    ele[26][19] != ele[29][20];
    ele[26][19] != ele[29][21];
    ele[26][19] != ele[29][22];
    ele[26][19] != ele[29][23];
    ele[26][19] != ele[30][19];
    ele[26][19] != ele[31][19];
    ele[26][19] != ele[32][19];
    ele[26][19] != ele[33][19];
    ele[26][19] != ele[34][19];
    ele[26][19] != ele[35][19];
    ele[26][2] != ele[26][10];
    ele[26][2] != ele[26][11];
    ele[26][2] != ele[26][12];
    ele[26][2] != ele[26][13];
    ele[26][2] != ele[26][14];
    ele[26][2] != ele[26][15];
    ele[26][2] != ele[26][16];
    ele[26][2] != ele[26][17];
    ele[26][2] != ele[26][18];
    ele[26][2] != ele[26][19];
    ele[26][2] != ele[26][20];
    ele[26][2] != ele[26][21];
    ele[26][2] != ele[26][22];
    ele[26][2] != ele[26][23];
    ele[26][2] != ele[26][24];
    ele[26][2] != ele[26][25];
    ele[26][2] != ele[26][26];
    ele[26][2] != ele[26][27];
    ele[26][2] != ele[26][28];
    ele[26][2] != ele[26][29];
    ele[26][2] != ele[26][3];
    ele[26][2] != ele[26][30];
    ele[26][2] != ele[26][31];
    ele[26][2] != ele[26][32];
    ele[26][2] != ele[26][33];
    ele[26][2] != ele[26][34];
    ele[26][2] != ele[26][35];
    ele[26][2] != ele[26][4];
    ele[26][2] != ele[26][5];
    ele[26][2] != ele[26][6];
    ele[26][2] != ele[26][7];
    ele[26][2] != ele[26][8];
    ele[26][2] != ele[26][9];
    ele[26][2] != ele[27][0];
    ele[26][2] != ele[27][1];
    ele[26][2] != ele[27][2];
    ele[26][2] != ele[27][3];
    ele[26][2] != ele[27][4];
    ele[26][2] != ele[27][5];
    ele[26][2] != ele[28][0];
    ele[26][2] != ele[28][1];
    ele[26][2] != ele[28][2];
    ele[26][2] != ele[28][3];
    ele[26][2] != ele[28][4];
    ele[26][2] != ele[28][5];
    ele[26][2] != ele[29][0];
    ele[26][2] != ele[29][1];
    ele[26][2] != ele[29][2];
    ele[26][2] != ele[29][3];
    ele[26][2] != ele[29][4];
    ele[26][2] != ele[29][5];
    ele[26][2] != ele[30][2];
    ele[26][2] != ele[31][2];
    ele[26][2] != ele[32][2];
    ele[26][2] != ele[33][2];
    ele[26][2] != ele[34][2];
    ele[26][2] != ele[35][2];
    ele[26][20] != ele[26][21];
    ele[26][20] != ele[26][22];
    ele[26][20] != ele[26][23];
    ele[26][20] != ele[26][24];
    ele[26][20] != ele[26][25];
    ele[26][20] != ele[26][26];
    ele[26][20] != ele[26][27];
    ele[26][20] != ele[26][28];
    ele[26][20] != ele[26][29];
    ele[26][20] != ele[26][30];
    ele[26][20] != ele[26][31];
    ele[26][20] != ele[26][32];
    ele[26][20] != ele[26][33];
    ele[26][20] != ele[26][34];
    ele[26][20] != ele[26][35];
    ele[26][20] != ele[27][18];
    ele[26][20] != ele[27][19];
    ele[26][20] != ele[27][20];
    ele[26][20] != ele[27][21];
    ele[26][20] != ele[27][22];
    ele[26][20] != ele[27][23];
    ele[26][20] != ele[28][18];
    ele[26][20] != ele[28][19];
    ele[26][20] != ele[28][20];
    ele[26][20] != ele[28][21];
    ele[26][20] != ele[28][22];
    ele[26][20] != ele[28][23];
    ele[26][20] != ele[29][18];
    ele[26][20] != ele[29][19];
    ele[26][20] != ele[29][20];
    ele[26][20] != ele[29][21];
    ele[26][20] != ele[29][22];
    ele[26][20] != ele[29][23];
    ele[26][20] != ele[30][20];
    ele[26][20] != ele[31][20];
    ele[26][20] != ele[32][20];
    ele[26][20] != ele[33][20];
    ele[26][20] != ele[34][20];
    ele[26][20] != ele[35][20];
    ele[26][21] != ele[26][22];
    ele[26][21] != ele[26][23];
    ele[26][21] != ele[26][24];
    ele[26][21] != ele[26][25];
    ele[26][21] != ele[26][26];
    ele[26][21] != ele[26][27];
    ele[26][21] != ele[26][28];
    ele[26][21] != ele[26][29];
    ele[26][21] != ele[26][30];
    ele[26][21] != ele[26][31];
    ele[26][21] != ele[26][32];
    ele[26][21] != ele[26][33];
    ele[26][21] != ele[26][34];
    ele[26][21] != ele[26][35];
    ele[26][21] != ele[27][18];
    ele[26][21] != ele[27][19];
    ele[26][21] != ele[27][20];
    ele[26][21] != ele[27][21];
    ele[26][21] != ele[27][22];
    ele[26][21] != ele[27][23];
    ele[26][21] != ele[28][18];
    ele[26][21] != ele[28][19];
    ele[26][21] != ele[28][20];
    ele[26][21] != ele[28][21];
    ele[26][21] != ele[28][22];
    ele[26][21] != ele[28][23];
    ele[26][21] != ele[29][18];
    ele[26][21] != ele[29][19];
    ele[26][21] != ele[29][20];
    ele[26][21] != ele[29][21];
    ele[26][21] != ele[29][22];
    ele[26][21] != ele[29][23];
    ele[26][21] != ele[30][21];
    ele[26][21] != ele[31][21];
    ele[26][21] != ele[32][21];
    ele[26][21] != ele[33][21];
    ele[26][21] != ele[34][21];
    ele[26][21] != ele[35][21];
    ele[26][22] != ele[26][23];
    ele[26][22] != ele[26][24];
    ele[26][22] != ele[26][25];
    ele[26][22] != ele[26][26];
    ele[26][22] != ele[26][27];
    ele[26][22] != ele[26][28];
    ele[26][22] != ele[26][29];
    ele[26][22] != ele[26][30];
    ele[26][22] != ele[26][31];
    ele[26][22] != ele[26][32];
    ele[26][22] != ele[26][33];
    ele[26][22] != ele[26][34];
    ele[26][22] != ele[26][35];
    ele[26][22] != ele[27][18];
    ele[26][22] != ele[27][19];
    ele[26][22] != ele[27][20];
    ele[26][22] != ele[27][21];
    ele[26][22] != ele[27][22];
    ele[26][22] != ele[27][23];
    ele[26][22] != ele[28][18];
    ele[26][22] != ele[28][19];
    ele[26][22] != ele[28][20];
    ele[26][22] != ele[28][21];
    ele[26][22] != ele[28][22];
    ele[26][22] != ele[28][23];
    ele[26][22] != ele[29][18];
    ele[26][22] != ele[29][19];
    ele[26][22] != ele[29][20];
    ele[26][22] != ele[29][21];
    ele[26][22] != ele[29][22];
    ele[26][22] != ele[29][23];
    ele[26][22] != ele[30][22];
    ele[26][22] != ele[31][22];
    ele[26][22] != ele[32][22];
    ele[26][22] != ele[33][22];
    ele[26][22] != ele[34][22];
    ele[26][22] != ele[35][22];
    ele[26][23] != ele[26][24];
    ele[26][23] != ele[26][25];
    ele[26][23] != ele[26][26];
    ele[26][23] != ele[26][27];
    ele[26][23] != ele[26][28];
    ele[26][23] != ele[26][29];
    ele[26][23] != ele[26][30];
    ele[26][23] != ele[26][31];
    ele[26][23] != ele[26][32];
    ele[26][23] != ele[26][33];
    ele[26][23] != ele[26][34];
    ele[26][23] != ele[26][35];
    ele[26][23] != ele[27][18];
    ele[26][23] != ele[27][19];
    ele[26][23] != ele[27][20];
    ele[26][23] != ele[27][21];
    ele[26][23] != ele[27][22];
    ele[26][23] != ele[27][23];
    ele[26][23] != ele[28][18];
    ele[26][23] != ele[28][19];
    ele[26][23] != ele[28][20];
    ele[26][23] != ele[28][21];
    ele[26][23] != ele[28][22];
    ele[26][23] != ele[28][23];
    ele[26][23] != ele[29][18];
    ele[26][23] != ele[29][19];
    ele[26][23] != ele[29][20];
    ele[26][23] != ele[29][21];
    ele[26][23] != ele[29][22];
    ele[26][23] != ele[29][23];
    ele[26][23] != ele[30][23];
    ele[26][23] != ele[31][23];
    ele[26][23] != ele[32][23];
    ele[26][23] != ele[33][23];
    ele[26][23] != ele[34][23];
    ele[26][23] != ele[35][23];
    ele[26][24] != ele[26][25];
    ele[26][24] != ele[26][26];
    ele[26][24] != ele[26][27];
    ele[26][24] != ele[26][28];
    ele[26][24] != ele[26][29];
    ele[26][24] != ele[26][30];
    ele[26][24] != ele[26][31];
    ele[26][24] != ele[26][32];
    ele[26][24] != ele[26][33];
    ele[26][24] != ele[26][34];
    ele[26][24] != ele[26][35];
    ele[26][24] != ele[27][24];
    ele[26][24] != ele[27][25];
    ele[26][24] != ele[27][26];
    ele[26][24] != ele[27][27];
    ele[26][24] != ele[27][28];
    ele[26][24] != ele[27][29];
    ele[26][24] != ele[28][24];
    ele[26][24] != ele[28][25];
    ele[26][24] != ele[28][26];
    ele[26][24] != ele[28][27];
    ele[26][24] != ele[28][28];
    ele[26][24] != ele[28][29];
    ele[26][24] != ele[29][24];
    ele[26][24] != ele[29][25];
    ele[26][24] != ele[29][26];
    ele[26][24] != ele[29][27];
    ele[26][24] != ele[29][28];
    ele[26][24] != ele[29][29];
    ele[26][24] != ele[30][24];
    ele[26][24] != ele[31][24];
    ele[26][24] != ele[32][24];
    ele[26][24] != ele[33][24];
    ele[26][24] != ele[34][24];
    ele[26][24] != ele[35][24];
    ele[26][25] != ele[26][26];
    ele[26][25] != ele[26][27];
    ele[26][25] != ele[26][28];
    ele[26][25] != ele[26][29];
    ele[26][25] != ele[26][30];
    ele[26][25] != ele[26][31];
    ele[26][25] != ele[26][32];
    ele[26][25] != ele[26][33];
    ele[26][25] != ele[26][34];
    ele[26][25] != ele[26][35];
    ele[26][25] != ele[27][24];
    ele[26][25] != ele[27][25];
    ele[26][25] != ele[27][26];
    ele[26][25] != ele[27][27];
    ele[26][25] != ele[27][28];
    ele[26][25] != ele[27][29];
    ele[26][25] != ele[28][24];
    ele[26][25] != ele[28][25];
    ele[26][25] != ele[28][26];
    ele[26][25] != ele[28][27];
    ele[26][25] != ele[28][28];
    ele[26][25] != ele[28][29];
    ele[26][25] != ele[29][24];
    ele[26][25] != ele[29][25];
    ele[26][25] != ele[29][26];
    ele[26][25] != ele[29][27];
    ele[26][25] != ele[29][28];
    ele[26][25] != ele[29][29];
    ele[26][25] != ele[30][25];
    ele[26][25] != ele[31][25];
    ele[26][25] != ele[32][25];
    ele[26][25] != ele[33][25];
    ele[26][25] != ele[34][25];
    ele[26][25] != ele[35][25];
    ele[26][26] != ele[26][27];
    ele[26][26] != ele[26][28];
    ele[26][26] != ele[26][29];
    ele[26][26] != ele[26][30];
    ele[26][26] != ele[26][31];
    ele[26][26] != ele[26][32];
    ele[26][26] != ele[26][33];
    ele[26][26] != ele[26][34];
    ele[26][26] != ele[26][35];
    ele[26][26] != ele[27][24];
    ele[26][26] != ele[27][25];
    ele[26][26] != ele[27][26];
    ele[26][26] != ele[27][27];
    ele[26][26] != ele[27][28];
    ele[26][26] != ele[27][29];
    ele[26][26] != ele[28][24];
    ele[26][26] != ele[28][25];
    ele[26][26] != ele[28][26];
    ele[26][26] != ele[28][27];
    ele[26][26] != ele[28][28];
    ele[26][26] != ele[28][29];
    ele[26][26] != ele[29][24];
    ele[26][26] != ele[29][25];
    ele[26][26] != ele[29][26];
    ele[26][26] != ele[29][27];
    ele[26][26] != ele[29][28];
    ele[26][26] != ele[29][29];
    ele[26][26] != ele[30][26];
    ele[26][26] != ele[31][26];
    ele[26][26] != ele[32][26];
    ele[26][26] != ele[33][26];
    ele[26][26] != ele[34][26];
    ele[26][26] != ele[35][26];
    ele[26][27] != ele[26][28];
    ele[26][27] != ele[26][29];
    ele[26][27] != ele[26][30];
    ele[26][27] != ele[26][31];
    ele[26][27] != ele[26][32];
    ele[26][27] != ele[26][33];
    ele[26][27] != ele[26][34];
    ele[26][27] != ele[26][35];
    ele[26][27] != ele[27][24];
    ele[26][27] != ele[27][25];
    ele[26][27] != ele[27][26];
    ele[26][27] != ele[27][27];
    ele[26][27] != ele[27][28];
    ele[26][27] != ele[27][29];
    ele[26][27] != ele[28][24];
    ele[26][27] != ele[28][25];
    ele[26][27] != ele[28][26];
    ele[26][27] != ele[28][27];
    ele[26][27] != ele[28][28];
    ele[26][27] != ele[28][29];
    ele[26][27] != ele[29][24];
    ele[26][27] != ele[29][25];
    ele[26][27] != ele[29][26];
    ele[26][27] != ele[29][27];
    ele[26][27] != ele[29][28];
    ele[26][27] != ele[29][29];
    ele[26][27] != ele[30][27];
    ele[26][27] != ele[31][27];
    ele[26][27] != ele[32][27];
    ele[26][27] != ele[33][27];
    ele[26][27] != ele[34][27];
    ele[26][27] != ele[35][27];
    ele[26][28] != ele[26][29];
    ele[26][28] != ele[26][30];
    ele[26][28] != ele[26][31];
    ele[26][28] != ele[26][32];
    ele[26][28] != ele[26][33];
    ele[26][28] != ele[26][34];
    ele[26][28] != ele[26][35];
    ele[26][28] != ele[27][24];
    ele[26][28] != ele[27][25];
    ele[26][28] != ele[27][26];
    ele[26][28] != ele[27][27];
    ele[26][28] != ele[27][28];
    ele[26][28] != ele[27][29];
    ele[26][28] != ele[28][24];
    ele[26][28] != ele[28][25];
    ele[26][28] != ele[28][26];
    ele[26][28] != ele[28][27];
    ele[26][28] != ele[28][28];
    ele[26][28] != ele[28][29];
    ele[26][28] != ele[29][24];
    ele[26][28] != ele[29][25];
    ele[26][28] != ele[29][26];
    ele[26][28] != ele[29][27];
    ele[26][28] != ele[29][28];
    ele[26][28] != ele[29][29];
    ele[26][28] != ele[30][28];
    ele[26][28] != ele[31][28];
    ele[26][28] != ele[32][28];
    ele[26][28] != ele[33][28];
    ele[26][28] != ele[34][28];
    ele[26][28] != ele[35][28];
    ele[26][29] != ele[26][30];
    ele[26][29] != ele[26][31];
    ele[26][29] != ele[26][32];
    ele[26][29] != ele[26][33];
    ele[26][29] != ele[26][34];
    ele[26][29] != ele[26][35];
    ele[26][29] != ele[27][24];
    ele[26][29] != ele[27][25];
    ele[26][29] != ele[27][26];
    ele[26][29] != ele[27][27];
    ele[26][29] != ele[27][28];
    ele[26][29] != ele[27][29];
    ele[26][29] != ele[28][24];
    ele[26][29] != ele[28][25];
    ele[26][29] != ele[28][26];
    ele[26][29] != ele[28][27];
    ele[26][29] != ele[28][28];
    ele[26][29] != ele[28][29];
    ele[26][29] != ele[29][24];
    ele[26][29] != ele[29][25];
    ele[26][29] != ele[29][26];
    ele[26][29] != ele[29][27];
    ele[26][29] != ele[29][28];
    ele[26][29] != ele[29][29];
    ele[26][29] != ele[30][29];
    ele[26][29] != ele[31][29];
    ele[26][29] != ele[32][29];
    ele[26][29] != ele[33][29];
    ele[26][29] != ele[34][29];
    ele[26][29] != ele[35][29];
    ele[26][3] != ele[26][10];
    ele[26][3] != ele[26][11];
    ele[26][3] != ele[26][12];
    ele[26][3] != ele[26][13];
    ele[26][3] != ele[26][14];
    ele[26][3] != ele[26][15];
    ele[26][3] != ele[26][16];
    ele[26][3] != ele[26][17];
    ele[26][3] != ele[26][18];
    ele[26][3] != ele[26][19];
    ele[26][3] != ele[26][20];
    ele[26][3] != ele[26][21];
    ele[26][3] != ele[26][22];
    ele[26][3] != ele[26][23];
    ele[26][3] != ele[26][24];
    ele[26][3] != ele[26][25];
    ele[26][3] != ele[26][26];
    ele[26][3] != ele[26][27];
    ele[26][3] != ele[26][28];
    ele[26][3] != ele[26][29];
    ele[26][3] != ele[26][30];
    ele[26][3] != ele[26][31];
    ele[26][3] != ele[26][32];
    ele[26][3] != ele[26][33];
    ele[26][3] != ele[26][34];
    ele[26][3] != ele[26][35];
    ele[26][3] != ele[26][4];
    ele[26][3] != ele[26][5];
    ele[26][3] != ele[26][6];
    ele[26][3] != ele[26][7];
    ele[26][3] != ele[26][8];
    ele[26][3] != ele[26][9];
    ele[26][3] != ele[27][0];
    ele[26][3] != ele[27][1];
    ele[26][3] != ele[27][2];
    ele[26][3] != ele[27][3];
    ele[26][3] != ele[27][4];
    ele[26][3] != ele[27][5];
    ele[26][3] != ele[28][0];
    ele[26][3] != ele[28][1];
    ele[26][3] != ele[28][2];
    ele[26][3] != ele[28][3];
    ele[26][3] != ele[28][4];
    ele[26][3] != ele[28][5];
    ele[26][3] != ele[29][0];
    ele[26][3] != ele[29][1];
    ele[26][3] != ele[29][2];
    ele[26][3] != ele[29][3];
    ele[26][3] != ele[29][4];
    ele[26][3] != ele[29][5];
    ele[26][3] != ele[30][3];
    ele[26][3] != ele[31][3];
    ele[26][3] != ele[32][3];
    ele[26][3] != ele[33][3];
    ele[26][3] != ele[34][3];
    ele[26][3] != ele[35][3];
    ele[26][30] != ele[26][31];
    ele[26][30] != ele[26][32];
    ele[26][30] != ele[26][33];
    ele[26][30] != ele[26][34];
    ele[26][30] != ele[26][35];
    ele[26][30] != ele[27][30];
    ele[26][30] != ele[27][31];
    ele[26][30] != ele[27][32];
    ele[26][30] != ele[27][33];
    ele[26][30] != ele[27][34];
    ele[26][30] != ele[27][35];
    ele[26][30] != ele[28][30];
    ele[26][30] != ele[28][31];
    ele[26][30] != ele[28][32];
    ele[26][30] != ele[28][33];
    ele[26][30] != ele[28][34];
    ele[26][30] != ele[28][35];
    ele[26][30] != ele[29][30];
    ele[26][30] != ele[29][31];
    ele[26][30] != ele[29][32];
    ele[26][30] != ele[29][33];
    ele[26][30] != ele[29][34];
    ele[26][30] != ele[29][35];
    ele[26][30] != ele[30][30];
    ele[26][30] != ele[31][30];
    ele[26][30] != ele[32][30];
    ele[26][30] != ele[33][30];
    ele[26][30] != ele[34][30];
    ele[26][30] != ele[35][30];
    ele[26][31] != ele[26][32];
    ele[26][31] != ele[26][33];
    ele[26][31] != ele[26][34];
    ele[26][31] != ele[26][35];
    ele[26][31] != ele[27][30];
    ele[26][31] != ele[27][31];
    ele[26][31] != ele[27][32];
    ele[26][31] != ele[27][33];
    ele[26][31] != ele[27][34];
    ele[26][31] != ele[27][35];
    ele[26][31] != ele[28][30];
    ele[26][31] != ele[28][31];
    ele[26][31] != ele[28][32];
    ele[26][31] != ele[28][33];
    ele[26][31] != ele[28][34];
    ele[26][31] != ele[28][35];
    ele[26][31] != ele[29][30];
    ele[26][31] != ele[29][31];
    ele[26][31] != ele[29][32];
    ele[26][31] != ele[29][33];
    ele[26][31] != ele[29][34];
    ele[26][31] != ele[29][35];
    ele[26][31] != ele[30][31];
    ele[26][31] != ele[31][31];
    ele[26][31] != ele[32][31];
    ele[26][31] != ele[33][31];
    ele[26][31] != ele[34][31];
    ele[26][31] != ele[35][31];
    ele[26][32] != ele[26][33];
    ele[26][32] != ele[26][34];
    ele[26][32] != ele[26][35];
    ele[26][32] != ele[27][30];
    ele[26][32] != ele[27][31];
    ele[26][32] != ele[27][32];
    ele[26][32] != ele[27][33];
    ele[26][32] != ele[27][34];
    ele[26][32] != ele[27][35];
    ele[26][32] != ele[28][30];
    ele[26][32] != ele[28][31];
    ele[26][32] != ele[28][32];
    ele[26][32] != ele[28][33];
    ele[26][32] != ele[28][34];
    ele[26][32] != ele[28][35];
    ele[26][32] != ele[29][30];
    ele[26][32] != ele[29][31];
    ele[26][32] != ele[29][32];
    ele[26][32] != ele[29][33];
    ele[26][32] != ele[29][34];
    ele[26][32] != ele[29][35];
    ele[26][32] != ele[30][32];
    ele[26][32] != ele[31][32];
    ele[26][32] != ele[32][32];
    ele[26][32] != ele[33][32];
    ele[26][32] != ele[34][32];
    ele[26][32] != ele[35][32];
    ele[26][33] != ele[26][34];
    ele[26][33] != ele[26][35];
    ele[26][33] != ele[27][30];
    ele[26][33] != ele[27][31];
    ele[26][33] != ele[27][32];
    ele[26][33] != ele[27][33];
    ele[26][33] != ele[27][34];
    ele[26][33] != ele[27][35];
    ele[26][33] != ele[28][30];
    ele[26][33] != ele[28][31];
    ele[26][33] != ele[28][32];
    ele[26][33] != ele[28][33];
    ele[26][33] != ele[28][34];
    ele[26][33] != ele[28][35];
    ele[26][33] != ele[29][30];
    ele[26][33] != ele[29][31];
    ele[26][33] != ele[29][32];
    ele[26][33] != ele[29][33];
    ele[26][33] != ele[29][34];
    ele[26][33] != ele[29][35];
    ele[26][33] != ele[30][33];
    ele[26][33] != ele[31][33];
    ele[26][33] != ele[32][33];
    ele[26][33] != ele[33][33];
    ele[26][33] != ele[34][33];
    ele[26][33] != ele[35][33];
    ele[26][34] != ele[26][35];
    ele[26][34] != ele[27][30];
    ele[26][34] != ele[27][31];
    ele[26][34] != ele[27][32];
    ele[26][34] != ele[27][33];
    ele[26][34] != ele[27][34];
    ele[26][34] != ele[27][35];
    ele[26][34] != ele[28][30];
    ele[26][34] != ele[28][31];
    ele[26][34] != ele[28][32];
    ele[26][34] != ele[28][33];
    ele[26][34] != ele[28][34];
    ele[26][34] != ele[28][35];
    ele[26][34] != ele[29][30];
    ele[26][34] != ele[29][31];
    ele[26][34] != ele[29][32];
    ele[26][34] != ele[29][33];
    ele[26][34] != ele[29][34];
    ele[26][34] != ele[29][35];
    ele[26][34] != ele[30][34];
    ele[26][34] != ele[31][34];
    ele[26][34] != ele[32][34];
    ele[26][34] != ele[33][34];
    ele[26][34] != ele[34][34];
    ele[26][34] != ele[35][34];
    ele[26][35] != ele[27][30];
    ele[26][35] != ele[27][31];
    ele[26][35] != ele[27][32];
    ele[26][35] != ele[27][33];
    ele[26][35] != ele[27][34];
    ele[26][35] != ele[27][35];
    ele[26][35] != ele[28][30];
    ele[26][35] != ele[28][31];
    ele[26][35] != ele[28][32];
    ele[26][35] != ele[28][33];
    ele[26][35] != ele[28][34];
    ele[26][35] != ele[28][35];
    ele[26][35] != ele[29][30];
    ele[26][35] != ele[29][31];
    ele[26][35] != ele[29][32];
    ele[26][35] != ele[29][33];
    ele[26][35] != ele[29][34];
    ele[26][35] != ele[29][35];
    ele[26][35] != ele[30][35];
    ele[26][35] != ele[31][35];
    ele[26][35] != ele[32][35];
    ele[26][35] != ele[33][35];
    ele[26][35] != ele[34][35];
    ele[26][35] != ele[35][35];
    ele[26][4] != ele[26][10];
    ele[26][4] != ele[26][11];
    ele[26][4] != ele[26][12];
    ele[26][4] != ele[26][13];
    ele[26][4] != ele[26][14];
    ele[26][4] != ele[26][15];
    ele[26][4] != ele[26][16];
    ele[26][4] != ele[26][17];
    ele[26][4] != ele[26][18];
    ele[26][4] != ele[26][19];
    ele[26][4] != ele[26][20];
    ele[26][4] != ele[26][21];
    ele[26][4] != ele[26][22];
    ele[26][4] != ele[26][23];
    ele[26][4] != ele[26][24];
    ele[26][4] != ele[26][25];
    ele[26][4] != ele[26][26];
    ele[26][4] != ele[26][27];
    ele[26][4] != ele[26][28];
    ele[26][4] != ele[26][29];
    ele[26][4] != ele[26][30];
    ele[26][4] != ele[26][31];
    ele[26][4] != ele[26][32];
    ele[26][4] != ele[26][33];
    ele[26][4] != ele[26][34];
    ele[26][4] != ele[26][35];
    ele[26][4] != ele[26][5];
    ele[26][4] != ele[26][6];
    ele[26][4] != ele[26][7];
    ele[26][4] != ele[26][8];
    ele[26][4] != ele[26][9];
    ele[26][4] != ele[27][0];
    ele[26][4] != ele[27][1];
    ele[26][4] != ele[27][2];
    ele[26][4] != ele[27][3];
    ele[26][4] != ele[27][4];
    ele[26][4] != ele[27][5];
    ele[26][4] != ele[28][0];
    ele[26][4] != ele[28][1];
    ele[26][4] != ele[28][2];
    ele[26][4] != ele[28][3];
    ele[26][4] != ele[28][4];
    ele[26][4] != ele[28][5];
    ele[26][4] != ele[29][0];
    ele[26][4] != ele[29][1];
    ele[26][4] != ele[29][2];
    ele[26][4] != ele[29][3];
    ele[26][4] != ele[29][4];
    ele[26][4] != ele[29][5];
    ele[26][4] != ele[30][4];
    ele[26][4] != ele[31][4];
    ele[26][4] != ele[32][4];
    ele[26][4] != ele[33][4];
    ele[26][4] != ele[34][4];
    ele[26][4] != ele[35][4];
    ele[26][5] != ele[26][10];
    ele[26][5] != ele[26][11];
    ele[26][5] != ele[26][12];
    ele[26][5] != ele[26][13];
    ele[26][5] != ele[26][14];
    ele[26][5] != ele[26][15];
    ele[26][5] != ele[26][16];
    ele[26][5] != ele[26][17];
    ele[26][5] != ele[26][18];
    ele[26][5] != ele[26][19];
    ele[26][5] != ele[26][20];
    ele[26][5] != ele[26][21];
    ele[26][5] != ele[26][22];
    ele[26][5] != ele[26][23];
    ele[26][5] != ele[26][24];
    ele[26][5] != ele[26][25];
    ele[26][5] != ele[26][26];
    ele[26][5] != ele[26][27];
    ele[26][5] != ele[26][28];
    ele[26][5] != ele[26][29];
    ele[26][5] != ele[26][30];
    ele[26][5] != ele[26][31];
    ele[26][5] != ele[26][32];
    ele[26][5] != ele[26][33];
    ele[26][5] != ele[26][34];
    ele[26][5] != ele[26][35];
    ele[26][5] != ele[26][6];
    ele[26][5] != ele[26][7];
    ele[26][5] != ele[26][8];
    ele[26][5] != ele[26][9];
    ele[26][5] != ele[27][0];
    ele[26][5] != ele[27][1];
    ele[26][5] != ele[27][2];
    ele[26][5] != ele[27][3];
    ele[26][5] != ele[27][4];
    ele[26][5] != ele[27][5];
    ele[26][5] != ele[28][0];
    ele[26][5] != ele[28][1];
    ele[26][5] != ele[28][2];
    ele[26][5] != ele[28][3];
    ele[26][5] != ele[28][4];
    ele[26][5] != ele[28][5];
    ele[26][5] != ele[29][0];
    ele[26][5] != ele[29][1];
    ele[26][5] != ele[29][2];
    ele[26][5] != ele[29][3];
    ele[26][5] != ele[29][4];
    ele[26][5] != ele[29][5];
    ele[26][5] != ele[30][5];
    ele[26][5] != ele[31][5];
    ele[26][5] != ele[32][5];
    ele[26][5] != ele[33][5];
    ele[26][5] != ele[34][5];
    ele[26][5] != ele[35][5];
    ele[26][6] != ele[26][10];
    ele[26][6] != ele[26][11];
    ele[26][6] != ele[26][12];
    ele[26][6] != ele[26][13];
    ele[26][6] != ele[26][14];
    ele[26][6] != ele[26][15];
    ele[26][6] != ele[26][16];
    ele[26][6] != ele[26][17];
    ele[26][6] != ele[26][18];
    ele[26][6] != ele[26][19];
    ele[26][6] != ele[26][20];
    ele[26][6] != ele[26][21];
    ele[26][6] != ele[26][22];
    ele[26][6] != ele[26][23];
    ele[26][6] != ele[26][24];
    ele[26][6] != ele[26][25];
    ele[26][6] != ele[26][26];
    ele[26][6] != ele[26][27];
    ele[26][6] != ele[26][28];
    ele[26][6] != ele[26][29];
    ele[26][6] != ele[26][30];
    ele[26][6] != ele[26][31];
    ele[26][6] != ele[26][32];
    ele[26][6] != ele[26][33];
    ele[26][6] != ele[26][34];
    ele[26][6] != ele[26][35];
    ele[26][6] != ele[26][7];
    ele[26][6] != ele[26][8];
    ele[26][6] != ele[26][9];
    ele[26][6] != ele[27][10];
    ele[26][6] != ele[27][11];
    ele[26][6] != ele[27][6];
    ele[26][6] != ele[27][7];
    ele[26][6] != ele[27][8];
    ele[26][6] != ele[27][9];
    ele[26][6] != ele[28][10];
    ele[26][6] != ele[28][11];
    ele[26][6] != ele[28][6];
    ele[26][6] != ele[28][7];
    ele[26][6] != ele[28][8];
    ele[26][6] != ele[28][9];
    ele[26][6] != ele[29][10];
    ele[26][6] != ele[29][11];
    ele[26][6] != ele[29][6];
    ele[26][6] != ele[29][7];
    ele[26][6] != ele[29][8];
    ele[26][6] != ele[29][9];
    ele[26][6] != ele[30][6];
    ele[26][6] != ele[31][6];
    ele[26][6] != ele[32][6];
    ele[26][6] != ele[33][6];
    ele[26][6] != ele[34][6];
    ele[26][6] != ele[35][6];
    ele[26][7] != ele[26][10];
    ele[26][7] != ele[26][11];
    ele[26][7] != ele[26][12];
    ele[26][7] != ele[26][13];
    ele[26][7] != ele[26][14];
    ele[26][7] != ele[26][15];
    ele[26][7] != ele[26][16];
    ele[26][7] != ele[26][17];
    ele[26][7] != ele[26][18];
    ele[26][7] != ele[26][19];
    ele[26][7] != ele[26][20];
    ele[26][7] != ele[26][21];
    ele[26][7] != ele[26][22];
    ele[26][7] != ele[26][23];
    ele[26][7] != ele[26][24];
    ele[26][7] != ele[26][25];
    ele[26][7] != ele[26][26];
    ele[26][7] != ele[26][27];
    ele[26][7] != ele[26][28];
    ele[26][7] != ele[26][29];
    ele[26][7] != ele[26][30];
    ele[26][7] != ele[26][31];
    ele[26][7] != ele[26][32];
    ele[26][7] != ele[26][33];
    ele[26][7] != ele[26][34];
    ele[26][7] != ele[26][35];
    ele[26][7] != ele[26][8];
    ele[26][7] != ele[26][9];
    ele[26][7] != ele[27][10];
    ele[26][7] != ele[27][11];
    ele[26][7] != ele[27][6];
    ele[26][7] != ele[27][7];
    ele[26][7] != ele[27][8];
    ele[26][7] != ele[27][9];
    ele[26][7] != ele[28][10];
    ele[26][7] != ele[28][11];
    ele[26][7] != ele[28][6];
    ele[26][7] != ele[28][7];
    ele[26][7] != ele[28][8];
    ele[26][7] != ele[28][9];
    ele[26][7] != ele[29][10];
    ele[26][7] != ele[29][11];
    ele[26][7] != ele[29][6];
    ele[26][7] != ele[29][7];
    ele[26][7] != ele[29][8];
    ele[26][7] != ele[29][9];
    ele[26][7] != ele[30][7];
    ele[26][7] != ele[31][7];
    ele[26][7] != ele[32][7];
    ele[26][7] != ele[33][7];
    ele[26][7] != ele[34][7];
    ele[26][7] != ele[35][7];
    ele[26][8] != ele[26][10];
    ele[26][8] != ele[26][11];
    ele[26][8] != ele[26][12];
    ele[26][8] != ele[26][13];
    ele[26][8] != ele[26][14];
    ele[26][8] != ele[26][15];
    ele[26][8] != ele[26][16];
    ele[26][8] != ele[26][17];
    ele[26][8] != ele[26][18];
    ele[26][8] != ele[26][19];
    ele[26][8] != ele[26][20];
    ele[26][8] != ele[26][21];
    ele[26][8] != ele[26][22];
    ele[26][8] != ele[26][23];
    ele[26][8] != ele[26][24];
    ele[26][8] != ele[26][25];
    ele[26][8] != ele[26][26];
    ele[26][8] != ele[26][27];
    ele[26][8] != ele[26][28];
    ele[26][8] != ele[26][29];
    ele[26][8] != ele[26][30];
    ele[26][8] != ele[26][31];
    ele[26][8] != ele[26][32];
    ele[26][8] != ele[26][33];
    ele[26][8] != ele[26][34];
    ele[26][8] != ele[26][35];
    ele[26][8] != ele[26][9];
    ele[26][8] != ele[27][10];
    ele[26][8] != ele[27][11];
    ele[26][8] != ele[27][6];
    ele[26][8] != ele[27][7];
    ele[26][8] != ele[27][8];
    ele[26][8] != ele[27][9];
    ele[26][8] != ele[28][10];
    ele[26][8] != ele[28][11];
    ele[26][8] != ele[28][6];
    ele[26][8] != ele[28][7];
    ele[26][8] != ele[28][8];
    ele[26][8] != ele[28][9];
    ele[26][8] != ele[29][10];
    ele[26][8] != ele[29][11];
    ele[26][8] != ele[29][6];
    ele[26][8] != ele[29][7];
    ele[26][8] != ele[29][8];
    ele[26][8] != ele[29][9];
    ele[26][8] != ele[30][8];
    ele[26][8] != ele[31][8];
    ele[26][8] != ele[32][8];
    ele[26][8] != ele[33][8];
    ele[26][8] != ele[34][8];
    ele[26][8] != ele[35][8];
    ele[26][9] != ele[26][10];
    ele[26][9] != ele[26][11];
    ele[26][9] != ele[26][12];
    ele[26][9] != ele[26][13];
    ele[26][9] != ele[26][14];
    ele[26][9] != ele[26][15];
    ele[26][9] != ele[26][16];
    ele[26][9] != ele[26][17];
    ele[26][9] != ele[26][18];
    ele[26][9] != ele[26][19];
    ele[26][9] != ele[26][20];
    ele[26][9] != ele[26][21];
    ele[26][9] != ele[26][22];
    ele[26][9] != ele[26][23];
    ele[26][9] != ele[26][24];
    ele[26][9] != ele[26][25];
    ele[26][9] != ele[26][26];
    ele[26][9] != ele[26][27];
    ele[26][9] != ele[26][28];
    ele[26][9] != ele[26][29];
    ele[26][9] != ele[26][30];
    ele[26][9] != ele[26][31];
    ele[26][9] != ele[26][32];
    ele[26][9] != ele[26][33];
    ele[26][9] != ele[26][34];
    ele[26][9] != ele[26][35];
    ele[26][9] != ele[27][10];
    ele[26][9] != ele[27][11];
    ele[26][9] != ele[27][6];
    ele[26][9] != ele[27][7];
    ele[26][9] != ele[27][8];
    ele[26][9] != ele[27][9];
    ele[26][9] != ele[28][10];
    ele[26][9] != ele[28][11];
    ele[26][9] != ele[28][6];
    ele[26][9] != ele[28][7];
    ele[26][9] != ele[28][8];
    ele[26][9] != ele[28][9];
    ele[26][9] != ele[29][10];
    ele[26][9] != ele[29][11];
    ele[26][9] != ele[29][6];
    ele[26][9] != ele[29][7];
    ele[26][9] != ele[29][8];
    ele[26][9] != ele[29][9];
    ele[26][9] != ele[30][9];
    ele[26][9] != ele[31][9];
    ele[26][9] != ele[32][9];
    ele[26][9] != ele[33][9];
    ele[26][9] != ele[34][9];
    ele[26][9] != ele[35][9];
    ele[27][0] != ele[27][1];
    ele[27][0] != ele[27][10];
    ele[27][0] != ele[27][11];
    ele[27][0] != ele[27][12];
    ele[27][0] != ele[27][13];
    ele[27][0] != ele[27][14];
    ele[27][0] != ele[27][15];
    ele[27][0] != ele[27][16];
    ele[27][0] != ele[27][17];
    ele[27][0] != ele[27][18];
    ele[27][0] != ele[27][19];
    ele[27][0] != ele[27][2];
    ele[27][0] != ele[27][20];
    ele[27][0] != ele[27][21];
    ele[27][0] != ele[27][22];
    ele[27][0] != ele[27][23];
    ele[27][0] != ele[27][24];
    ele[27][0] != ele[27][25];
    ele[27][0] != ele[27][26];
    ele[27][0] != ele[27][27];
    ele[27][0] != ele[27][28];
    ele[27][0] != ele[27][29];
    ele[27][0] != ele[27][3];
    ele[27][0] != ele[27][30];
    ele[27][0] != ele[27][31];
    ele[27][0] != ele[27][32];
    ele[27][0] != ele[27][33];
    ele[27][0] != ele[27][34];
    ele[27][0] != ele[27][35];
    ele[27][0] != ele[27][4];
    ele[27][0] != ele[27][5];
    ele[27][0] != ele[27][6];
    ele[27][0] != ele[27][7];
    ele[27][0] != ele[27][8];
    ele[27][0] != ele[27][9];
    ele[27][0] != ele[28][0];
    ele[27][0] != ele[28][1];
    ele[27][0] != ele[28][2];
    ele[27][0] != ele[28][3];
    ele[27][0] != ele[28][4];
    ele[27][0] != ele[28][5];
    ele[27][0] != ele[29][0];
    ele[27][0] != ele[29][1];
    ele[27][0] != ele[29][2];
    ele[27][0] != ele[29][3];
    ele[27][0] != ele[29][4];
    ele[27][0] != ele[29][5];
    ele[27][0] != ele[30][0];
    ele[27][0] != ele[31][0];
    ele[27][0] != ele[32][0];
    ele[27][0] != ele[33][0];
    ele[27][0] != ele[34][0];
    ele[27][0] != ele[35][0];
    ele[27][1] != ele[27][10];
    ele[27][1] != ele[27][11];
    ele[27][1] != ele[27][12];
    ele[27][1] != ele[27][13];
    ele[27][1] != ele[27][14];
    ele[27][1] != ele[27][15];
    ele[27][1] != ele[27][16];
    ele[27][1] != ele[27][17];
    ele[27][1] != ele[27][18];
    ele[27][1] != ele[27][19];
    ele[27][1] != ele[27][2];
    ele[27][1] != ele[27][20];
    ele[27][1] != ele[27][21];
    ele[27][1] != ele[27][22];
    ele[27][1] != ele[27][23];
    ele[27][1] != ele[27][24];
    ele[27][1] != ele[27][25];
    ele[27][1] != ele[27][26];
    ele[27][1] != ele[27][27];
    ele[27][1] != ele[27][28];
    ele[27][1] != ele[27][29];
    ele[27][1] != ele[27][3];
    ele[27][1] != ele[27][30];
    ele[27][1] != ele[27][31];
    ele[27][1] != ele[27][32];
    ele[27][1] != ele[27][33];
    ele[27][1] != ele[27][34];
    ele[27][1] != ele[27][35];
    ele[27][1] != ele[27][4];
    ele[27][1] != ele[27][5];
    ele[27][1] != ele[27][6];
    ele[27][1] != ele[27][7];
    ele[27][1] != ele[27][8];
    ele[27][1] != ele[27][9];
    ele[27][1] != ele[28][0];
    ele[27][1] != ele[28][1];
    ele[27][1] != ele[28][2];
    ele[27][1] != ele[28][3];
    ele[27][1] != ele[28][4];
    ele[27][1] != ele[28][5];
    ele[27][1] != ele[29][0];
    ele[27][1] != ele[29][1];
    ele[27][1] != ele[29][2];
    ele[27][1] != ele[29][3];
    ele[27][1] != ele[29][4];
    ele[27][1] != ele[29][5];
    ele[27][1] != ele[30][1];
    ele[27][1] != ele[31][1];
    ele[27][1] != ele[32][1];
    ele[27][1] != ele[33][1];
    ele[27][1] != ele[34][1];
    ele[27][1] != ele[35][1];
    ele[27][10] != ele[27][11];
    ele[27][10] != ele[27][12];
    ele[27][10] != ele[27][13];
    ele[27][10] != ele[27][14];
    ele[27][10] != ele[27][15];
    ele[27][10] != ele[27][16];
    ele[27][10] != ele[27][17];
    ele[27][10] != ele[27][18];
    ele[27][10] != ele[27][19];
    ele[27][10] != ele[27][20];
    ele[27][10] != ele[27][21];
    ele[27][10] != ele[27][22];
    ele[27][10] != ele[27][23];
    ele[27][10] != ele[27][24];
    ele[27][10] != ele[27][25];
    ele[27][10] != ele[27][26];
    ele[27][10] != ele[27][27];
    ele[27][10] != ele[27][28];
    ele[27][10] != ele[27][29];
    ele[27][10] != ele[27][30];
    ele[27][10] != ele[27][31];
    ele[27][10] != ele[27][32];
    ele[27][10] != ele[27][33];
    ele[27][10] != ele[27][34];
    ele[27][10] != ele[27][35];
    ele[27][10] != ele[28][10];
    ele[27][10] != ele[28][11];
    ele[27][10] != ele[28][6];
    ele[27][10] != ele[28][7];
    ele[27][10] != ele[28][8];
    ele[27][10] != ele[28][9];
    ele[27][10] != ele[29][10];
    ele[27][10] != ele[29][11];
    ele[27][10] != ele[29][6];
    ele[27][10] != ele[29][7];
    ele[27][10] != ele[29][8];
    ele[27][10] != ele[29][9];
    ele[27][10] != ele[30][10];
    ele[27][10] != ele[31][10];
    ele[27][10] != ele[32][10];
    ele[27][10] != ele[33][10];
    ele[27][10] != ele[34][10];
    ele[27][10] != ele[35][10];
    ele[27][11] != ele[27][12];
    ele[27][11] != ele[27][13];
    ele[27][11] != ele[27][14];
    ele[27][11] != ele[27][15];
    ele[27][11] != ele[27][16];
    ele[27][11] != ele[27][17];
    ele[27][11] != ele[27][18];
    ele[27][11] != ele[27][19];
    ele[27][11] != ele[27][20];
    ele[27][11] != ele[27][21];
    ele[27][11] != ele[27][22];
    ele[27][11] != ele[27][23];
    ele[27][11] != ele[27][24];
    ele[27][11] != ele[27][25];
    ele[27][11] != ele[27][26];
    ele[27][11] != ele[27][27];
    ele[27][11] != ele[27][28];
    ele[27][11] != ele[27][29];
    ele[27][11] != ele[27][30];
    ele[27][11] != ele[27][31];
    ele[27][11] != ele[27][32];
    ele[27][11] != ele[27][33];
    ele[27][11] != ele[27][34];
    ele[27][11] != ele[27][35];
    ele[27][11] != ele[28][10];
    ele[27][11] != ele[28][11];
    ele[27][11] != ele[28][6];
    ele[27][11] != ele[28][7];
    ele[27][11] != ele[28][8];
    ele[27][11] != ele[28][9];
    ele[27][11] != ele[29][10];
    ele[27][11] != ele[29][11];
    ele[27][11] != ele[29][6];
    ele[27][11] != ele[29][7];
    ele[27][11] != ele[29][8];
    ele[27][11] != ele[29][9];
    ele[27][11] != ele[30][11];
    ele[27][11] != ele[31][11];
    ele[27][11] != ele[32][11];
    ele[27][11] != ele[33][11];
    ele[27][11] != ele[34][11];
    ele[27][11] != ele[35][11];
    ele[27][12] != ele[27][13];
    ele[27][12] != ele[27][14];
    ele[27][12] != ele[27][15];
    ele[27][12] != ele[27][16];
    ele[27][12] != ele[27][17];
    ele[27][12] != ele[27][18];
    ele[27][12] != ele[27][19];
    ele[27][12] != ele[27][20];
    ele[27][12] != ele[27][21];
    ele[27][12] != ele[27][22];
    ele[27][12] != ele[27][23];
    ele[27][12] != ele[27][24];
    ele[27][12] != ele[27][25];
    ele[27][12] != ele[27][26];
    ele[27][12] != ele[27][27];
    ele[27][12] != ele[27][28];
    ele[27][12] != ele[27][29];
    ele[27][12] != ele[27][30];
    ele[27][12] != ele[27][31];
    ele[27][12] != ele[27][32];
    ele[27][12] != ele[27][33];
    ele[27][12] != ele[27][34];
    ele[27][12] != ele[27][35];
    ele[27][12] != ele[28][12];
    ele[27][12] != ele[28][13];
    ele[27][12] != ele[28][14];
    ele[27][12] != ele[28][15];
    ele[27][12] != ele[28][16];
    ele[27][12] != ele[28][17];
    ele[27][12] != ele[29][12];
    ele[27][12] != ele[29][13];
    ele[27][12] != ele[29][14];
    ele[27][12] != ele[29][15];
    ele[27][12] != ele[29][16];
    ele[27][12] != ele[29][17];
    ele[27][12] != ele[30][12];
    ele[27][12] != ele[31][12];
    ele[27][12] != ele[32][12];
    ele[27][12] != ele[33][12];
    ele[27][12] != ele[34][12];
    ele[27][12] != ele[35][12];
    ele[27][13] != ele[27][14];
    ele[27][13] != ele[27][15];
    ele[27][13] != ele[27][16];
    ele[27][13] != ele[27][17];
    ele[27][13] != ele[27][18];
    ele[27][13] != ele[27][19];
    ele[27][13] != ele[27][20];
    ele[27][13] != ele[27][21];
    ele[27][13] != ele[27][22];
    ele[27][13] != ele[27][23];
    ele[27][13] != ele[27][24];
    ele[27][13] != ele[27][25];
    ele[27][13] != ele[27][26];
    ele[27][13] != ele[27][27];
    ele[27][13] != ele[27][28];
    ele[27][13] != ele[27][29];
    ele[27][13] != ele[27][30];
    ele[27][13] != ele[27][31];
    ele[27][13] != ele[27][32];
    ele[27][13] != ele[27][33];
    ele[27][13] != ele[27][34];
    ele[27][13] != ele[27][35];
    ele[27][13] != ele[28][12];
    ele[27][13] != ele[28][13];
    ele[27][13] != ele[28][14];
    ele[27][13] != ele[28][15];
    ele[27][13] != ele[28][16];
    ele[27][13] != ele[28][17];
    ele[27][13] != ele[29][12];
    ele[27][13] != ele[29][13];
    ele[27][13] != ele[29][14];
    ele[27][13] != ele[29][15];
    ele[27][13] != ele[29][16];
    ele[27][13] != ele[29][17];
    ele[27][13] != ele[30][13];
    ele[27][13] != ele[31][13];
    ele[27][13] != ele[32][13];
    ele[27][13] != ele[33][13];
    ele[27][13] != ele[34][13];
    ele[27][13] != ele[35][13];
    ele[27][14] != ele[27][15];
    ele[27][14] != ele[27][16];
    ele[27][14] != ele[27][17];
    ele[27][14] != ele[27][18];
    ele[27][14] != ele[27][19];
    ele[27][14] != ele[27][20];
    ele[27][14] != ele[27][21];
    ele[27][14] != ele[27][22];
    ele[27][14] != ele[27][23];
    ele[27][14] != ele[27][24];
    ele[27][14] != ele[27][25];
    ele[27][14] != ele[27][26];
    ele[27][14] != ele[27][27];
    ele[27][14] != ele[27][28];
    ele[27][14] != ele[27][29];
    ele[27][14] != ele[27][30];
    ele[27][14] != ele[27][31];
    ele[27][14] != ele[27][32];
    ele[27][14] != ele[27][33];
    ele[27][14] != ele[27][34];
    ele[27][14] != ele[27][35];
    ele[27][14] != ele[28][12];
    ele[27][14] != ele[28][13];
    ele[27][14] != ele[28][14];
    ele[27][14] != ele[28][15];
    ele[27][14] != ele[28][16];
    ele[27][14] != ele[28][17];
    ele[27][14] != ele[29][12];
    ele[27][14] != ele[29][13];
    ele[27][14] != ele[29][14];
    ele[27][14] != ele[29][15];
    ele[27][14] != ele[29][16];
    ele[27][14] != ele[29][17];
    ele[27][14] != ele[30][14];
    ele[27][14] != ele[31][14];
    ele[27][14] != ele[32][14];
    ele[27][14] != ele[33][14];
    ele[27][14] != ele[34][14];
    ele[27][14] != ele[35][14];
    ele[27][15] != ele[27][16];
    ele[27][15] != ele[27][17];
    ele[27][15] != ele[27][18];
    ele[27][15] != ele[27][19];
    ele[27][15] != ele[27][20];
    ele[27][15] != ele[27][21];
    ele[27][15] != ele[27][22];
    ele[27][15] != ele[27][23];
    ele[27][15] != ele[27][24];
    ele[27][15] != ele[27][25];
    ele[27][15] != ele[27][26];
    ele[27][15] != ele[27][27];
    ele[27][15] != ele[27][28];
    ele[27][15] != ele[27][29];
    ele[27][15] != ele[27][30];
    ele[27][15] != ele[27][31];
    ele[27][15] != ele[27][32];
    ele[27][15] != ele[27][33];
    ele[27][15] != ele[27][34];
    ele[27][15] != ele[27][35];
    ele[27][15] != ele[28][12];
    ele[27][15] != ele[28][13];
    ele[27][15] != ele[28][14];
    ele[27][15] != ele[28][15];
    ele[27][15] != ele[28][16];
    ele[27][15] != ele[28][17];
    ele[27][15] != ele[29][12];
    ele[27][15] != ele[29][13];
    ele[27][15] != ele[29][14];
    ele[27][15] != ele[29][15];
    ele[27][15] != ele[29][16];
    ele[27][15] != ele[29][17];
    ele[27][15] != ele[30][15];
    ele[27][15] != ele[31][15];
    ele[27][15] != ele[32][15];
    ele[27][15] != ele[33][15];
    ele[27][15] != ele[34][15];
    ele[27][15] != ele[35][15];
    ele[27][16] != ele[27][17];
    ele[27][16] != ele[27][18];
    ele[27][16] != ele[27][19];
    ele[27][16] != ele[27][20];
    ele[27][16] != ele[27][21];
    ele[27][16] != ele[27][22];
    ele[27][16] != ele[27][23];
    ele[27][16] != ele[27][24];
    ele[27][16] != ele[27][25];
    ele[27][16] != ele[27][26];
    ele[27][16] != ele[27][27];
    ele[27][16] != ele[27][28];
    ele[27][16] != ele[27][29];
    ele[27][16] != ele[27][30];
    ele[27][16] != ele[27][31];
    ele[27][16] != ele[27][32];
    ele[27][16] != ele[27][33];
    ele[27][16] != ele[27][34];
    ele[27][16] != ele[27][35];
    ele[27][16] != ele[28][12];
    ele[27][16] != ele[28][13];
    ele[27][16] != ele[28][14];
    ele[27][16] != ele[28][15];
    ele[27][16] != ele[28][16];
    ele[27][16] != ele[28][17];
    ele[27][16] != ele[29][12];
    ele[27][16] != ele[29][13];
    ele[27][16] != ele[29][14];
    ele[27][16] != ele[29][15];
    ele[27][16] != ele[29][16];
    ele[27][16] != ele[29][17];
    ele[27][16] != ele[30][16];
    ele[27][16] != ele[31][16];
    ele[27][16] != ele[32][16];
    ele[27][16] != ele[33][16];
    ele[27][16] != ele[34][16];
    ele[27][16] != ele[35][16];
    ele[27][17] != ele[27][18];
    ele[27][17] != ele[27][19];
    ele[27][17] != ele[27][20];
    ele[27][17] != ele[27][21];
    ele[27][17] != ele[27][22];
    ele[27][17] != ele[27][23];
    ele[27][17] != ele[27][24];
    ele[27][17] != ele[27][25];
    ele[27][17] != ele[27][26];
    ele[27][17] != ele[27][27];
    ele[27][17] != ele[27][28];
    ele[27][17] != ele[27][29];
    ele[27][17] != ele[27][30];
    ele[27][17] != ele[27][31];
    ele[27][17] != ele[27][32];
    ele[27][17] != ele[27][33];
    ele[27][17] != ele[27][34];
    ele[27][17] != ele[27][35];
    ele[27][17] != ele[28][12];
    ele[27][17] != ele[28][13];
    ele[27][17] != ele[28][14];
    ele[27][17] != ele[28][15];
    ele[27][17] != ele[28][16];
    ele[27][17] != ele[28][17];
    ele[27][17] != ele[29][12];
    ele[27][17] != ele[29][13];
    ele[27][17] != ele[29][14];
    ele[27][17] != ele[29][15];
    ele[27][17] != ele[29][16];
    ele[27][17] != ele[29][17];
    ele[27][17] != ele[30][17];
    ele[27][17] != ele[31][17];
    ele[27][17] != ele[32][17];
    ele[27][17] != ele[33][17];
    ele[27][17] != ele[34][17];
    ele[27][17] != ele[35][17];
    ele[27][18] != ele[27][19];
    ele[27][18] != ele[27][20];
    ele[27][18] != ele[27][21];
    ele[27][18] != ele[27][22];
    ele[27][18] != ele[27][23];
    ele[27][18] != ele[27][24];
    ele[27][18] != ele[27][25];
    ele[27][18] != ele[27][26];
    ele[27][18] != ele[27][27];
    ele[27][18] != ele[27][28];
    ele[27][18] != ele[27][29];
    ele[27][18] != ele[27][30];
    ele[27][18] != ele[27][31];
    ele[27][18] != ele[27][32];
    ele[27][18] != ele[27][33];
    ele[27][18] != ele[27][34];
    ele[27][18] != ele[27][35];
    ele[27][18] != ele[28][18];
    ele[27][18] != ele[28][19];
    ele[27][18] != ele[28][20];
    ele[27][18] != ele[28][21];
    ele[27][18] != ele[28][22];
    ele[27][18] != ele[28][23];
    ele[27][18] != ele[29][18];
    ele[27][18] != ele[29][19];
    ele[27][18] != ele[29][20];
    ele[27][18] != ele[29][21];
    ele[27][18] != ele[29][22];
    ele[27][18] != ele[29][23];
    ele[27][18] != ele[30][18];
    ele[27][18] != ele[31][18];
    ele[27][18] != ele[32][18];
    ele[27][18] != ele[33][18];
    ele[27][18] != ele[34][18];
    ele[27][18] != ele[35][18];
    ele[27][19] != ele[27][20];
    ele[27][19] != ele[27][21];
    ele[27][19] != ele[27][22];
    ele[27][19] != ele[27][23];
    ele[27][19] != ele[27][24];
    ele[27][19] != ele[27][25];
    ele[27][19] != ele[27][26];
    ele[27][19] != ele[27][27];
    ele[27][19] != ele[27][28];
    ele[27][19] != ele[27][29];
    ele[27][19] != ele[27][30];
    ele[27][19] != ele[27][31];
    ele[27][19] != ele[27][32];
    ele[27][19] != ele[27][33];
    ele[27][19] != ele[27][34];
    ele[27][19] != ele[27][35];
    ele[27][19] != ele[28][18];
    ele[27][19] != ele[28][19];
    ele[27][19] != ele[28][20];
    ele[27][19] != ele[28][21];
    ele[27][19] != ele[28][22];
    ele[27][19] != ele[28][23];
    ele[27][19] != ele[29][18];
    ele[27][19] != ele[29][19];
    ele[27][19] != ele[29][20];
    ele[27][19] != ele[29][21];
    ele[27][19] != ele[29][22];
    ele[27][19] != ele[29][23];
    ele[27][19] != ele[30][19];
    ele[27][19] != ele[31][19];
    ele[27][19] != ele[32][19];
    ele[27][19] != ele[33][19];
    ele[27][19] != ele[34][19];
    ele[27][19] != ele[35][19];
    ele[27][2] != ele[27][10];
    ele[27][2] != ele[27][11];
    ele[27][2] != ele[27][12];
    ele[27][2] != ele[27][13];
    ele[27][2] != ele[27][14];
    ele[27][2] != ele[27][15];
    ele[27][2] != ele[27][16];
    ele[27][2] != ele[27][17];
    ele[27][2] != ele[27][18];
    ele[27][2] != ele[27][19];
    ele[27][2] != ele[27][20];
    ele[27][2] != ele[27][21];
    ele[27][2] != ele[27][22];
    ele[27][2] != ele[27][23];
    ele[27][2] != ele[27][24];
    ele[27][2] != ele[27][25];
    ele[27][2] != ele[27][26];
    ele[27][2] != ele[27][27];
    ele[27][2] != ele[27][28];
    ele[27][2] != ele[27][29];
    ele[27][2] != ele[27][3];
    ele[27][2] != ele[27][30];
    ele[27][2] != ele[27][31];
    ele[27][2] != ele[27][32];
    ele[27][2] != ele[27][33];
    ele[27][2] != ele[27][34];
    ele[27][2] != ele[27][35];
    ele[27][2] != ele[27][4];
    ele[27][2] != ele[27][5];
    ele[27][2] != ele[27][6];
    ele[27][2] != ele[27][7];
    ele[27][2] != ele[27][8];
    ele[27][2] != ele[27][9];
    ele[27][2] != ele[28][0];
    ele[27][2] != ele[28][1];
    ele[27][2] != ele[28][2];
    ele[27][2] != ele[28][3];
    ele[27][2] != ele[28][4];
    ele[27][2] != ele[28][5];
    ele[27][2] != ele[29][0];
    ele[27][2] != ele[29][1];
    ele[27][2] != ele[29][2];
    ele[27][2] != ele[29][3];
    ele[27][2] != ele[29][4];
    ele[27][2] != ele[29][5];
    ele[27][2] != ele[30][2];
    ele[27][2] != ele[31][2];
    ele[27][2] != ele[32][2];
    ele[27][2] != ele[33][2];
    ele[27][2] != ele[34][2];
    ele[27][2] != ele[35][2];
    ele[27][20] != ele[27][21];
    ele[27][20] != ele[27][22];
    ele[27][20] != ele[27][23];
    ele[27][20] != ele[27][24];
    ele[27][20] != ele[27][25];
    ele[27][20] != ele[27][26];
    ele[27][20] != ele[27][27];
    ele[27][20] != ele[27][28];
    ele[27][20] != ele[27][29];
    ele[27][20] != ele[27][30];
    ele[27][20] != ele[27][31];
    ele[27][20] != ele[27][32];
    ele[27][20] != ele[27][33];
    ele[27][20] != ele[27][34];
    ele[27][20] != ele[27][35];
    ele[27][20] != ele[28][18];
    ele[27][20] != ele[28][19];
    ele[27][20] != ele[28][20];
    ele[27][20] != ele[28][21];
    ele[27][20] != ele[28][22];
    ele[27][20] != ele[28][23];
    ele[27][20] != ele[29][18];
    ele[27][20] != ele[29][19];
    ele[27][20] != ele[29][20];
    ele[27][20] != ele[29][21];
    ele[27][20] != ele[29][22];
    ele[27][20] != ele[29][23];
    ele[27][20] != ele[30][20];
    ele[27][20] != ele[31][20];
    ele[27][20] != ele[32][20];
    ele[27][20] != ele[33][20];
    ele[27][20] != ele[34][20];
    ele[27][20] != ele[35][20];
    ele[27][21] != ele[27][22];
    ele[27][21] != ele[27][23];
    ele[27][21] != ele[27][24];
    ele[27][21] != ele[27][25];
    ele[27][21] != ele[27][26];
    ele[27][21] != ele[27][27];
    ele[27][21] != ele[27][28];
    ele[27][21] != ele[27][29];
    ele[27][21] != ele[27][30];
    ele[27][21] != ele[27][31];
    ele[27][21] != ele[27][32];
    ele[27][21] != ele[27][33];
    ele[27][21] != ele[27][34];
    ele[27][21] != ele[27][35];
    ele[27][21] != ele[28][18];
    ele[27][21] != ele[28][19];
    ele[27][21] != ele[28][20];
    ele[27][21] != ele[28][21];
    ele[27][21] != ele[28][22];
    ele[27][21] != ele[28][23];
    ele[27][21] != ele[29][18];
    ele[27][21] != ele[29][19];
    ele[27][21] != ele[29][20];
    ele[27][21] != ele[29][21];
    ele[27][21] != ele[29][22];
    ele[27][21] != ele[29][23];
    ele[27][21] != ele[30][21];
    ele[27][21] != ele[31][21];
    ele[27][21] != ele[32][21];
    ele[27][21] != ele[33][21];
    ele[27][21] != ele[34][21];
    ele[27][21] != ele[35][21];
    ele[27][22] != ele[27][23];
    ele[27][22] != ele[27][24];
    ele[27][22] != ele[27][25];
    ele[27][22] != ele[27][26];
    ele[27][22] != ele[27][27];
    ele[27][22] != ele[27][28];
    ele[27][22] != ele[27][29];
    ele[27][22] != ele[27][30];
    ele[27][22] != ele[27][31];
    ele[27][22] != ele[27][32];
    ele[27][22] != ele[27][33];
    ele[27][22] != ele[27][34];
    ele[27][22] != ele[27][35];
    ele[27][22] != ele[28][18];
    ele[27][22] != ele[28][19];
    ele[27][22] != ele[28][20];
    ele[27][22] != ele[28][21];
    ele[27][22] != ele[28][22];
    ele[27][22] != ele[28][23];
    ele[27][22] != ele[29][18];
    ele[27][22] != ele[29][19];
    ele[27][22] != ele[29][20];
    ele[27][22] != ele[29][21];
    ele[27][22] != ele[29][22];
    ele[27][22] != ele[29][23];
    ele[27][22] != ele[30][22];
    ele[27][22] != ele[31][22];
    ele[27][22] != ele[32][22];
    ele[27][22] != ele[33][22];
    ele[27][22] != ele[34][22];
    ele[27][22] != ele[35][22];
    ele[27][23] != ele[27][24];
    ele[27][23] != ele[27][25];
    ele[27][23] != ele[27][26];
    ele[27][23] != ele[27][27];
    ele[27][23] != ele[27][28];
    ele[27][23] != ele[27][29];
    ele[27][23] != ele[27][30];
    ele[27][23] != ele[27][31];
    ele[27][23] != ele[27][32];
    ele[27][23] != ele[27][33];
    ele[27][23] != ele[27][34];
    ele[27][23] != ele[27][35];
    ele[27][23] != ele[28][18];
    ele[27][23] != ele[28][19];
    ele[27][23] != ele[28][20];
    ele[27][23] != ele[28][21];
    ele[27][23] != ele[28][22];
    ele[27][23] != ele[28][23];
    ele[27][23] != ele[29][18];
    ele[27][23] != ele[29][19];
    ele[27][23] != ele[29][20];
    ele[27][23] != ele[29][21];
    ele[27][23] != ele[29][22];
    ele[27][23] != ele[29][23];
    ele[27][23] != ele[30][23];
    ele[27][23] != ele[31][23];
    ele[27][23] != ele[32][23];
    ele[27][23] != ele[33][23];
    ele[27][23] != ele[34][23];
    ele[27][23] != ele[35][23];
    ele[27][24] != ele[27][25];
    ele[27][24] != ele[27][26];
    ele[27][24] != ele[27][27];
    ele[27][24] != ele[27][28];
    ele[27][24] != ele[27][29];
    ele[27][24] != ele[27][30];
    ele[27][24] != ele[27][31];
    ele[27][24] != ele[27][32];
    ele[27][24] != ele[27][33];
    ele[27][24] != ele[27][34];
    ele[27][24] != ele[27][35];
    ele[27][24] != ele[28][24];
    ele[27][24] != ele[28][25];
    ele[27][24] != ele[28][26];
    ele[27][24] != ele[28][27];
    ele[27][24] != ele[28][28];
    ele[27][24] != ele[28][29];
    ele[27][24] != ele[29][24];
    ele[27][24] != ele[29][25];
    ele[27][24] != ele[29][26];
    ele[27][24] != ele[29][27];
    ele[27][24] != ele[29][28];
    ele[27][24] != ele[29][29];
    ele[27][24] != ele[30][24];
    ele[27][24] != ele[31][24];
    ele[27][24] != ele[32][24];
    ele[27][24] != ele[33][24];
    ele[27][24] != ele[34][24];
    ele[27][24] != ele[35][24];
    ele[27][25] != ele[27][26];
    ele[27][25] != ele[27][27];
    ele[27][25] != ele[27][28];
    ele[27][25] != ele[27][29];
    ele[27][25] != ele[27][30];
    ele[27][25] != ele[27][31];
    ele[27][25] != ele[27][32];
    ele[27][25] != ele[27][33];
    ele[27][25] != ele[27][34];
    ele[27][25] != ele[27][35];
    ele[27][25] != ele[28][24];
    ele[27][25] != ele[28][25];
    ele[27][25] != ele[28][26];
    ele[27][25] != ele[28][27];
    ele[27][25] != ele[28][28];
    ele[27][25] != ele[28][29];
    ele[27][25] != ele[29][24];
    ele[27][25] != ele[29][25];
    ele[27][25] != ele[29][26];
    ele[27][25] != ele[29][27];
    ele[27][25] != ele[29][28];
    ele[27][25] != ele[29][29];
    ele[27][25] != ele[30][25];
    ele[27][25] != ele[31][25];
    ele[27][25] != ele[32][25];
    ele[27][25] != ele[33][25];
    ele[27][25] != ele[34][25];
    ele[27][25] != ele[35][25];
    ele[27][26] != ele[27][27];
    ele[27][26] != ele[27][28];
    ele[27][26] != ele[27][29];
    ele[27][26] != ele[27][30];
    ele[27][26] != ele[27][31];
    ele[27][26] != ele[27][32];
    ele[27][26] != ele[27][33];
    ele[27][26] != ele[27][34];
    ele[27][26] != ele[27][35];
    ele[27][26] != ele[28][24];
    ele[27][26] != ele[28][25];
    ele[27][26] != ele[28][26];
    ele[27][26] != ele[28][27];
    ele[27][26] != ele[28][28];
    ele[27][26] != ele[28][29];
    ele[27][26] != ele[29][24];
    ele[27][26] != ele[29][25];
    ele[27][26] != ele[29][26];
    ele[27][26] != ele[29][27];
    ele[27][26] != ele[29][28];
    ele[27][26] != ele[29][29];
    ele[27][26] != ele[30][26];
    ele[27][26] != ele[31][26];
    ele[27][26] != ele[32][26];
    ele[27][26] != ele[33][26];
    ele[27][26] != ele[34][26];
    ele[27][26] != ele[35][26];
    ele[27][27] != ele[27][28];
    ele[27][27] != ele[27][29];
    ele[27][27] != ele[27][30];
    ele[27][27] != ele[27][31];
    ele[27][27] != ele[27][32];
    ele[27][27] != ele[27][33];
    ele[27][27] != ele[27][34];
    ele[27][27] != ele[27][35];
    ele[27][27] != ele[28][24];
    ele[27][27] != ele[28][25];
    ele[27][27] != ele[28][26];
    ele[27][27] != ele[28][27];
    ele[27][27] != ele[28][28];
    ele[27][27] != ele[28][29];
    ele[27][27] != ele[29][24];
    ele[27][27] != ele[29][25];
    ele[27][27] != ele[29][26];
    ele[27][27] != ele[29][27];
    ele[27][27] != ele[29][28];
    ele[27][27] != ele[29][29];
    ele[27][27] != ele[30][27];
    ele[27][27] != ele[31][27];
    ele[27][27] != ele[32][27];
    ele[27][27] != ele[33][27];
    ele[27][27] != ele[34][27];
    ele[27][27] != ele[35][27];
    ele[27][28] != ele[27][29];
    ele[27][28] != ele[27][30];
    ele[27][28] != ele[27][31];
    ele[27][28] != ele[27][32];
    ele[27][28] != ele[27][33];
    ele[27][28] != ele[27][34];
    ele[27][28] != ele[27][35];
    ele[27][28] != ele[28][24];
    ele[27][28] != ele[28][25];
    ele[27][28] != ele[28][26];
    ele[27][28] != ele[28][27];
    ele[27][28] != ele[28][28];
    ele[27][28] != ele[28][29];
    ele[27][28] != ele[29][24];
    ele[27][28] != ele[29][25];
    ele[27][28] != ele[29][26];
    ele[27][28] != ele[29][27];
    ele[27][28] != ele[29][28];
    ele[27][28] != ele[29][29];
    ele[27][28] != ele[30][28];
    ele[27][28] != ele[31][28];
    ele[27][28] != ele[32][28];
    ele[27][28] != ele[33][28];
    ele[27][28] != ele[34][28];
    ele[27][28] != ele[35][28];
    ele[27][29] != ele[27][30];
    ele[27][29] != ele[27][31];
    ele[27][29] != ele[27][32];
    ele[27][29] != ele[27][33];
    ele[27][29] != ele[27][34];
    ele[27][29] != ele[27][35];
    ele[27][29] != ele[28][24];
    ele[27][29] != ele[28][25];
    ele[27][29] != ele[28][26];
    ele[27][29] != ele[28][27];
    ele[27][29] != ele[28][28];
    ele[27][29] != ele[28][29];
    ele[27][29] != ele[29][24];
    ele[27][29] != ele[29][25];
    ele[27][29] != ele[29][26];
    ele[27][29] != ele[29][27];
    ele[27][29] != ele[29][28];
    ele[27][29] != ele[29][29];
    ele[27][29] != ele[30][29];
    ele[27][29] != ele[31][29];
    ele[27][29] != ele[32][29];
    ele[27][29] != ele[33][29];
    ele[27][29] != ele[34][29];
    ele[27][29] != ele[35][29];
    ele[27][3] != ele[27][10];
    ele[27][3] != ele[27][11];
    ele[27][3] != ele[27][12];
    ele[27][3] != ele[27][13];
    ele[27][3] != ele[27][14];
    ele[27][3] != ele[27][15];
    ele[27][3] != ele[27][16];
    ele[27][3] != ele[27][17];
    ele[27][3] != ele[27][18];
    ele[27][3] != ele[27][19];
    ele[27][3] != ele[27][20];
    ele[27][3] != ele[27][21];
    ele[27][3] != ele[27][22];
    ele[27][3] != ele[27][23];
    ele[27][3] != ele[27][24];
    ele[27][3] != ele[27][25];
    ele[27][3] != ele[27][26];
    ele[27][3] != ele[27][27];
    ele[27][3] != ele[27][28];
    ele[27][3] != ele[27][29];
    ele[27][3] != ele[27][30];
    ele[27][3] != ele[27][31];
    ele[27][3] != ele[27][32];
    ele[27][3] != ele[27][33];
    ele[27][3] != ele[27][34];
    ele[27][3] != ele[27][35];
    ele[27][3] != ele[27][4];
    ele[27][3] != ele[27][5];
    ele[27][3] != ele[27][6];
    ele[27][3] != ele[27][7];
    ele[27][3] != ele[27][8];
    ele[27][3] != ele[27][9];
    ele[27][3] != ele[28][0];
    ele[27][3] != ele[28][1];
    ele[27][3] != ele[28][2];
    ele[27][3] != ele[28][3];
    ele[27][3] != ele[28][4];
    ele[27][3] != ele[28][5];
    ele[27][3] != ele[29][0];
    ele[27][3] != ele[29][1];
    ele[27][3] != ele[29][2];
    ele[27][3] != ele[29][3];
    ele[27][3] != ele[29][4];
    ele[27][3] != ele[29][5];
    ele[27][3] != ele[30][3];
    ele[27][3] != ele[31][3];
    ele[27][3] != ele[32][3];
    ele[27][3] != ele[33][3];
    ele[27][3] != ele[34][3];
    ele[27][3] != ele[35][3];
    ele[27][30] != ele[27][31];
    ele[27][30] != ele[27][32];
    ele[27][30] != ele[27][33];
    ele[27][30] != ele[27][34];
    ele[27][30] != ele[27][35];
    ele[27][30] != ele[28][30];
    ele[27][30] != ele[28][31];
    ele[27][30] != ele[28][32];
    ele[27][30] != ele[28][33];
    ele[27][30] != ele[28][34];
    ele[27][30] != ele[28][35];
    ele[27][30] != ele[29][30];
    ele[27][30] != ele[29][31];
    ele[27][30] != ele[29][32];
    ele[27][30] != ele[29][33];
    ele[27][30] != ele[29][34];
    ele[27][30] != ele[29][35];
    ele[27][30] != ele[30][30];
    ele[27][30] != ele[31][30];
    ele[27][30] != ele[32][30];
    ele[27][30] != ele[33][30];
    ele[27][30] != ele[34][30];
    ele[27][30] != ele[35][30];
    ele[27][31] != ele[27][32];
    ele[27][31] != ele[27][33];
    ele[27][31] != ele[27][34];
    ele[27][31] != ele[27][35];
    ele[27][31] != ele[28][30];
    ele[27][31] != ele[28][31];
    ele[27][31] != ele[28][32];
    ele[27][31] != ele[28][33];
    ele[27][31] != ele[28][34];
    ele[27][31] != ele[28][35];
    ele[27][31] != ele[29][30];
    ele[27][31] != ele[29][31];
    ele[27][31] != ele[29][32];
    ele[27][31] != ele[29][33];
    ele[27][31] != ele[29][34];
    ele[27][31] != ele[29][35];
    ele[27][31] != ele[30][31];
    ele[27][31] != ele[31][31];
    ele[27][31] != ele[32][31];
    ele[27][31] != ele[33][31];
    ele[27][31] != ele[34][31];
    ele[27][31] != ele[35][31];
    ele[27][32] != ele[27][33];
    ele[27][32] != ele[27][34];
    ele[27][32] != ele[27][35];
    ele[27][32] != ele[28][30];
    ele[27][32] != ele[28][31];
    ele[27][32] != ele[28][32];
    ele[27][32] != ele[28][33];
    ele[27][32] != ele[28][34];
    ele[27][32] != ele[28][35];
    ele[27][32] != ele[29][30];
    ele[27][32] != ele[29][31];
    ele[27][32] != ele[29][32];
    ele[27][32] != ele[29][33];
    ele[27][32] != ele[29][34];
    ele[27][32] != ele[29][35];
    ele[27][32] != ele[30][32];
    ele[27][32] != ele[31][32];
    ele[27][32] != ele[32][32];
    ele[27][32] != ele[33][32];
    ele[27][32] != ele[34][32];
    ele[27][32] != ele[35][32];
    ele[27][33] != ele[27][34];
    ele[27][33] != ele[27][35];
    ele[27][33] != ele[28][30];
    ele[27][33] != ele[28][31];
    ele[27][33] != ele[28][32];
    ele[27][33] != ele[28][33];
    ele[27][33] != ele[28][34];
    ele[27][33] != ele[28][35];
    ele[27][33] != ele[29][30];
    ele[27][33] != ele[29][31];
    ele[27][33] != ele[29][32];
    ele[27][33] != ele[29][33];
    ele[27][33] != ele[29][34];
    ele[27][33] != ele[29][35];
    ele[27][33] != ele[30][33];
    ele[27][33] != ele[31][33];
    ele[27][33] != ele[32][33];
    ele[27][33] != ele[33][33];
    ele[27][33] != ele[34][33];
    ele[27][33] != ele[35][33];
    ele[27][34] != ele[27][35];
    ele[27][34] != ele[28][30];
    ele[27][34] != ele[28][31];
    ele[27][34] != ele[28][32];
    ele[27][34] != ele[28][33];
    ele[27][34] != ele[28][34];
    ele[27][34] != ele[28][35];
    ele[27][34] != ele[29][30];
    ele[27][34] != ele[29][31];
    ele[27][34] != ele[29][32];
    ele[27][34] != ele[29][33];
    ele[27][34] != ele[29][34];
    ele[27][34] != ele[29][35];
    ele[27][34] != ele[30][34];
    ele[27][34] != ele[31][34];
    ele[27][34] != ele[32][34];
    ele[27][34] != ele[33][34];
    ele[27][34] != ele[34][34];
    ele[27][34] != ele[35][34];
    ele[27][35] != ele[28][30];
    ele[27][35] != ele[28][31];
    ele[27][35] != ele[28][32];
    ele[27][35] != ele[28][33];
    ele[27][35] != ele[28][34];
    ele[27][35] != ele[28][35];
    ele[27][35] != ele[29][30];
    ele[27][35] != ele[29][31];
    ele[27][35] != ele[29][32];
    ele[27][35] != ele[29][33];
    ele[27][35] != ele[29][34];
    ele[27][35] != ele[29][35];
    ele[27][35] != ele[30][35];
    ele[27][35] != ele[31][35];
    ele[27][35] != ele[32][35];
    ele[27][35] != ele[33][35];
    ele[27][35] != ele[34][35];
    ele[27][35] != ele[35][35];
    ele[27][4] != ele[27][10];
    ele[27][4] != ele[27][11];
    ele[27][4] != ele[27][12];
    ele[27][4] != ele[27][13];
    ele[27][4] != ele[27][14];
    ele[27][4] != ele[27][15];
    ele[27][4] != ele[27][16];
    ele[27][4] != ele[27][17];
    ele[27][4] != ele[27][18];
    ele[27][4] != ele[27][19];
    ele[27][4] != ele[27][20];
    ele[27][4] != ele[27][21];
    ele[27][4] != ele[27][22];
    ele[27][4] != ele[27][23];
    ele[27][4] != ele[27][24];
    ele[27][4] != ele[27][25];
    ele[27][4] != ele[27][26];
    ele[27][4] != ele[27][27];
    ele[27][4] != ele[27][28];
    ele[27][4] != ele[27][29];
    ele[27][4] != ele[27][30];
    ele[27][4] != ele[27][31];
    ele[27][4] != ele[27][32];
    ele[27][4] != ele[27][33];
    ele[27][4] != ele[27][34];
    ele[27][4] != ele[27][35];
    ele[27][4] != ele[27][5];
    ele[27][4] != ele[27][6];
    ele[27][4] != ele[27][7];
    ele[27][4] != ele[27][8];
    ele[27][4] != ele[27][9];
    ele[27][4] != ele[28][0];
    ele[27][4] != ele[28][1];
    ele[27][4] != ele[28][2];
    ele[27][4] != ele[28][3];
    ele[27][4] != ele[28][4];
    ele[27][4] != ele[28][5];
    ele[27][4] != ele[29][0];
    ele[27][4] != ele[29][1];
    ele[27][4] != ele[29][2];
    ele[27][4] != ele[29][3];
    ele[27][4] != ele[29][4];
    ele[27][4] != ele[29][5];
    ele[27][4] != ele[30][4];
    ele[27][4] != ele[31][4];
    ele[27][4] != ele[32][4];
    ele[27][4] != ele[33][4];
    ele[27][4] != ele[34][4];
    ele[27][4] != ele[35][4];
    ele[27][5] != ele[27][10];
    ele[27][5] != ele[27][11];
    ele[27][5] != ele[27][12];
    ele[27][5] != ele[27][13];
    ele[27][5] != ele[27][14];
    ele[27][5] != ele[27][15];
    ele[27][5] != ele[27][16];
    ele[27][5] != ele[27][17];
    ele[27][5] != ele[27][18];
    ele[27][5] != ele[27][19];
    ele[27][5] != ele[27][20];
    ele[27][5] != ele[27][21];
    ele[27][5] != ele[27][22];
    ele[27][5] != ele[27][23];
    ele[27][5] != ele[27][24];
    ele[27][5] != ele[27][25];
    ele[27][5] != ele[27][26];
    ele[27][5] != ele[27][27];
    ele[27][5] != ele[27][28];
    ele[27][5] != ele[27][29];
    ele[27][5] != ele[27][30];
    ele[27][5] != ele[27][31];
    ele[27][5] != ele[27][32];
    ele[27][5] != ele[27][33];
    ele[27][5] != ele[27][34];
    ele[27][5] != ele[27][35];
    ele[27][5] != ele[27][6];
    ele[27][5] != ele[27][7];
    ele[27][5] != ele[27][8];
    ele[27][5] != ele[27][9];
    ele[27][5] != ele[28][0];
    ele[27][5] != ele[28][1];
    ele[27][5] != ele[28][2];
    ele[27][5] != ele[28][3];
    ele[27][5] != ele[28][4];
    ele[27][5] != ele[28][5];
    ele[27][5] != ele[29][0];
    ele[27][5] != ele[29][1];
    ele[27][5] != ele[29][2];
    ele[27][5] != ele[29][3];
    ele[27][5] != ele[29][4];
    ele[27][5] != ele[29][5];
    ele[27][5] != ele[30][5];
    ele[27][5] != ele[31][5];
    ele[27][5] != ele[32][5];
    ele[27][5] != ele[33][5];
    ele[27][5] != ele[34][5];
    ele[27][5] != ele[35][5];
    ele[27][6] != ele[27][10];
    ele[27][6] != ele[27][11];
    ele[27][6] != ele[27][12];
    ele[27][6] != ele[27][13];
    ele[27][6] != ele[27][14];
    ele[27][6] != ele[27][15];
    ele[27][6] != ele[27][16];
    ele[27][6] != ele[27][17];
    ele[27][6] != ele[27][18];
    ele[27][6] != ele[27][19];
    ele[27][6] != ele[27][20];
    ele[27][6] != ele[27][21];
    ele[27][6] != ele[27][22];
    ele[27][6] != ele[27][23];
    ele[27][6] != ele[27][24];
    ele[27][6] != ele[27][25];
    ele[27][6] != ele[27][26];
    ele[27][6] != ele[27][27];
    ele[27][6] != ele[27][28];
    ele[27][6] != ele[27][29];
    ele[27][6] != ele[27][30];
    ele[27][6] != ele[27][31];
    ele[27][6] != ele[27][32];
    ele[27][6] != ele[27][33];
    ele[27][6] != ele[27][34];
    ele[27][6] != ele[27][35];
    ele[27][6] != ele[27][7];
    ele[27][6] != ele[27][8];
    ele[27][6] != ele[27][9];
    ele[27][6] != ele[28][10];
    ele[27][6] != ele[28][11];
    ele[27][6] != ele[28][6];
    ele[27][6] != ele[28][7];
    ele[27][6] != ele[28][8];
    ele[27][6] != ele[28][9];
    ele[27][6] != ele[29][10];
    ele[27][6] != ele[29][11];
    ele[27][6] != ele[29][6];
    ele[27][6] != ele[29][7];
    ele[27][6] != ele[29][8];
    ele[27][6] != ele[29][9];
    ele[27][6] != ele[30][6];
    ele[27][6] != ele[31][6];
    ele[27][6] != ele[32][6];
    ele[27][6] != ele[33][6];
    ele[27][6] != ele[34][6];
    ele[27][6] != ele[35][6];
    ele[27][7] != ele[27][10];
    ele[27][7] != ele[27][11];
    ele[27][7] != ele[27][12];
    ele[27][7] != ele[27][13];
    ele[27][7] != ele[27][14];
    ele[27][7] != ele[27][15];
    ele[27][7] != ele[27][16];
    ele[27][7] != ele[27][17];
    ele[27][7] != ele[27][18];
    ele[27][7] != ele[27][19];
    ele[27][7] != ele[27][20];
    ele[27][7] != ele[27][21];
    ele[27][7] != ele[27][22];
    ele[27][7] != ele[27][23];
    ele[27][7] != ele[27][24];
    ele[27][7] != ele[27][25];
    ele[27][7] != ele[27][26];
    ele[27][7] != ele[27][27];
    ele[27][7] != ele[27][28];
    ele[27][7] != ele[27][29];
    ele[27][7] != ele[27][30];
    ele[27][7] != ele[27][31];
    ele[27][7] != ele[27][32];
    ele[27][7] != ele[27][33];
    ele[27][7] != ele[27][34];
    ele[27][7] != ele[27][35];
    ele[27][7] != ele[27][8];
    ele[27][7] != ele[27][9];
    ele[27][7] != ele[28][10];
    ele[27][7] != ele[28][11];
    ele[27][7] != ele[28][6];
    ele[27][7] != ele[28][7];
    ele[27][7] != ele[28][8];
    ele[27][7] != ele[28][9];
    ele[27][7] != ele[29][10];
    ele[27][7] != ele[29][11];
    ele[27][7] != ele[29][6];
    ele[27][7] != ele[29][7];
    ele[27][7] != ele[29][8];
    ele[27][7] != ele[29][9];
    ele[27][7] != ele[30][7];
    ele[27][7] != ele[31][7];
    ele[27][7] != ele[32][7];
    ele[27][7] != ele[33][7];
    ele[27][7] != ele[34][7];
    ele[27][7] != ele[35][7];
    ele[27][8] != ele[27][10];
    ele[27][8] != ele[27][11];
    ele[27][8] != ele[27][12];
    ele[27][8] != ele[27][13];
    ele[27][8] != ele[27][14];
    ele[27][8] != ele[27][15];
    ele[27][8] != ele[27][16];
    ele[27][8] != ele[27][17];
    ele[27][8] != ele[27][18];
    ele[27][8] != ele[27][19];
    ele[27][8] != ele[27][20];
    ele[27][8] != ele[27][21];
    ele[27][8] != ele[27][22];
    ele[27][8] != ele[27][23];
    ele[27][8] != ele[27][24];
    ele[27][8] != ele[27][25];
    ele[27][8] != ele[27][26];
    ele[27][8] != ele[27][27];
    ele[27][8] != ele[27][28];
    ele[27][8] != ele[27][29];
    ele[27][8] != ele[27][30];
    ele[27][8] != ele[27][31];
    ele[27][8] != ele[27][32];
    ele[27][8] != ele[27][33];
    ele[27][8] != ele[27][34];
    ele[27][8] != ele[27][35];
    ele[27][8] != ele[27][9];
    ele[27][8] != ele[28][10];
    ele[27][8] != ele[28][11];
    ele[27][8] != ele[28][6];
    ele[27][8] != ele[28][7];
    ele[27][8] != ele[28][8];
    ele[27][8] != ele[28][9];
    ele[27][8] != ele[29][10];
    ele[27][8] != ele[29][11];
    ele[27][8] != ele[29][6];
    ele[27][8] != ele[29][7];
    ele[27][8] != ele[29][8];
    ele[27][8] != ele[29][9];
    ele[27][8] != ele[30][8];
    ele[27][8] != ele[31][8];
    ele[27][8] != ele[32][8];
    ele[27][8] != ele[33][8];
    ele[27][8] != ele[34][8];
    ele[27][8] != ele[35][8];
    ele[27][9] != ele[27][10];
    ele[27][9] != ele[27][11];
    ele[27][9] != ele[27][12];
    ele[27][9] != ele[27][13];
    ele[27][9] != ele[27][14];
    ele[27][9] != ele[27][15];
    ele[27][9] != ele[27][16];
    ele[27][9] != ele[27][17];
    ele[27][9] != ele[27][18];
    ele[27][9] != ele[27][19];
    ele[27][9] != ele[27][20];
    ele[27][9] != ele[27][21];
    ele[27][9] != ele[27][22];
    ele[27][9] != ele[27][23];
    ele[27][9] != ele[27][24];
    ele[27][9] != ele[27][25];
    ele[27][9] != ele[27][26];
    ele[27][9] != ele[27][27];
    ele[27][9] != ele[27][28];
    ele[27][9] != ele[27][29];
    ele[27][9] != ele[27][30];
    ele[27][9] != ele[27][31];
    ele[27][9] != ele[27][32];
    ele[27][9] != ele[27][33];
    ele[27][9] != ele[27][34];
    ele[27][9] != ele[27][35];
    ele[27][9] != ele[28][10];
    ele[27][9] != ele[28][11];
    ele[27][9] != ele[28][6];
    ele[27][9] != ele[28][7];
    ele[27][9] != ele[28][8];
    ele[27][9] != ele[28][9];
    ele[27][9] != ele[29][10];
    ele[27][9] != ele[29][11];
    ele[27][9] != ele[29][6];
    ele[27][9] != ele[29][7];
    ele[27][9] != ele[29][8];
    ele[27][9] != ele[29][9];
    ele[27][9] != ele[30][9];
    ele[27][9] != ele[31][9];
    ele[27][9] != ele[32][9];
    ele[27][9] != ele[33][9];
    ele[27][9] != ele[34][9];
    ele[27][9] != ele[35][9];
    ele[28][0] != ele[28][1];
    ele[28][0] != ele[28][10];
    ele[28][0] != ele[28][11];
    ele[28][0] != ele[28][12];
    ele[28][0] != ele[28][13];
    ele[28][0] != ele[28][14];
    ele[28][0] != ele[28][15];
    ele[28][0] != ele[28][16];
    ele[28][0] != ele[28][17];
    ele[28][0] != ele[28][18];
    ele[28][0] != ele[28][19];
    ele[28][0] != ele[28][2];
    ele[28][0] != ele[28][20];
    ele[28][0] != ele[28][21];
    ele[28][0] != ele[28][22];
    ele[28][0] != ele[28][23];
    ele[28][0] != ele[28][24];
    ele[28][0] != ele[28][25];
    ele[28][0] != ele[28][26];
    ele[28][0] != ele[28][27];
    ele[28][0] != ele[28][28];
    ele[28][0] != ele[28][29];
    ele[28][0] != ele[28][3];
    ele[28][0] != ele[28][30];
    ele[28][0] != ele[28][31];
    ele[28][0] != ele[28][32];
    ele[28][0] != ele[28][33];
    ele[28][0] != ele[28][34];
    ele[28][0] != ele[28][35];
    ele[28][0] != ele[28][4];
    ele[28][0] != ele[28][5];
    ele[28][0] != ele[28][6];
    ele[28][0] != ele[28][7];
    ele[28][0] != ele[28][8];
    ele[28][0] != ele[28][9];
    ele[28][0] != ele[29][0];
    ele[28][0] != ele[29][1];
    ele[28][0] != ele[29][2];
    ele[28][0] != ele[29][3];
    ele[28][0] != ele[29][4];
    ele[28][0] != ele[29][5];
    ele[28][0] != ele[30][0];
    ele[28][0] != ele[31][0];
    ele[28][0] != ele[32][0];
    ele[28][0] != ele[33][0];
    ele[28][0] != ele[34][0];
    ele[28][0] != ele[35][0];
    ele[28][1] != ele[28][10];
    ele[28][1] != ele[28][11];
    ele[28][1] != ele[28][12];
    ele[28][1] != ele[28][13];
    ele[28][1] != ele[28][14];
    ele[28][1] != ele[28][15];
    ele[28][1] != ele[28][16];
    ele[28][1] != ele[28][17];
    ele[28][1] != ele[28][18];
    ele[28][1] != ele[28][19];
    ele[28][1] != ele[28][2];
    ele[28][1] != ele[28][20];
    ele[28][1] != ele[28][21];
    ele[28][1] != ele[28][22];
    ele[28][1] != ele[28][23];
    ele[28][1] != ele[28][24];
    ele[28][1] != ele[28][25];
    ele[28][1] != ele[28][26];
    ele[28][1] != ele[28][27];
    ele[28][1] != ele[28][28];
    ele[28][1] != ele[28][29];
    ele[28][1] != ele[28][3];
    ele[28][1] != ele[28][30];
    ele[28][1] != ele[28][31];
    ele[28][1] != ele[28][32];
    ele[28][1] != ele[28][33];
    ele[28][1] != ele[28][34];
    ele[28][1] != ele[28][35];
    ele[28][1] != ele[28][4];
    ele[28][1] != ele[28][5];
    ele[28][1] != ele[28][6];
    ele[28][1] != ele[28][7];
    ele[28][1] != ele[28][8];
    ele[28][1] != ele[28][9];
    ele[28][1] != ele[29][0];
    ele[28][1] != ele[29][1];
    ele[28][1] != ele[29][2];
    ele[28][1] != ele[29][3];
    ele[28][1] != ele[29][4];
    ele[28][1] != ele[29][5];
    ele[28][1] != ele[30][1];
    ele[28][1] != ele[31][1];
    ele[28][1] != ele[32][1];
    ele[28][1] != ele[33][1];
    ele[28][1] != ele[34][1];
    ele[28][1] != ele[35][1];
    ele[28][10] != ele[28][11];
    ele[28][10] != ele[28][12];
    ele[28][10] != ele[28][13];
    ele[28][10] != ele[28][14];
    ele[28][10] != ele[28][15];
    ele[28][10] != ele[28][16];
    ele[28][10] != ele[28][17];
    ele[28][10] != ele[28][18];
    ele[28][10] != ele[28][19];
    ele[28][10] != ele[28][20];
    ele[28][10] != ele[28][21];
    ele[28][10] != ele[28][22];
    ele[28][10] != ele[28][23];
    ele[28][10] != ele[28][24];
    ele[28][10] != ele[28][25];
    ele[28][10] != ele[28][26];
    ele[28][10] != ele[28][27];
    ele[28][10] != ele[28][28];
    ele[28][10] != ele[28][29];
    ele[28][10] != ele[28][30];
    ele[28][10] != ele[28][31];
    ele[28][10] != ele[28][32];
    ele[28][10] != ele[28][33];
    ele[28][10] != ele[28][34];
    ele[28][10] != ele[28][35];
    ele[28][10] != ele[29][10];
    ele[28][10] != ele[29][11];
    ele[28][10] != ele[29][6];
    ele[28][10] != ele[29][7];
    ele[28][10] != ele[29][8];
    ele[28][10] != ele[29][9];
    ele[28][10] != ele[30][10];
    ele[28][10] != ele[31][10];
    ele[28][10] != ele[32][10];
    ele[28][10] != ele[33][10];
    ele[28][10] != ele[34][10];
    ele[28][10] != ele[35][10];
    ele[28][11] != ele[28][12];
    ele[28][11] != ele[28][13];
    ele[28][11] != ele[28][14];
    ele[28][11] != ele[28][15];
    ele[28][11] != ele[28][16];
    ele[28][11] != ele[28][17];
    ele[28][11] != ele[28][18];
    ele[28][11] != ele[28][19];
    ele[28][11] != ele[28][20];
    ele[28][11] != ele[28][21];
    ele[28][11] != ele[28][22];
    ele[28][11] != ele[28][23];
    ele[28][11] != ele[28][24];
    ele[28][11] != ele[28][25];
    ele[28][11] != ele[28][26];
    ele[28][11] != ele[28][27];
    ele[28][11] != ele[28][28];
    ele[28][11] != ele[28][29];
    ele[28][11] != ele[28][30];
    ele[28][11] != ele[28][31];
    ele[28][11] != ele[28][32];
    ele[28][11] != ele[28][33];
    ele[28][11] != ele[28][34];
    ele[28][11] != ele[28][35];
    ele[28][11] != ele[29][10];
    ele[28][11] != ele[29][11];
    ele[28][11] != ele[29][6];
    ele[28][11] != ele[29][7];
    ele[28][11] != ele[29][8];
    ele[28][11] != ele[29][9];
    ele[28][11] != ele[30][11];
    ele[28][11] != ele[31][11];
    ele[28][11] != ele[32][11];
    ele[28][11] != ele[33][11];
    ele[28][11] != ele[34][11];
    ele[28][11] != ele[35][11];
    ele[28][12] != ele[28][13];
    ele[28][12] != ele[28][14];
    ele[28][12] != ele[28][15];
    ele[28][12] != ele[28][16];
    ele[28][12] != ele[28][17];
    ele[28][12] != ele[28][18];
    ele[28][12] != ele[28][19];
    ele[28][12] != ele[28][20];
    ele[28][12] != ele[28][21];
    ele[28][12] != ele[28][22];
    ele[28][12] != ele[28][23];
    ele[28][12] != ele[28][24];
    ele[28][12] != ele[28][25];
    ele[28][12] != ele[28][26];
    ele[28][12] != ele[28][27];
    ele[28][12] != ele[28][28];
    ele[28][12] != ele[28][29];
    ele[28][12] != ele[28][30];
    ele[28][12] != ele[28][31];
    ele[28][12] != ele[28][32];
    ele[28][12] != ele[28][33];
    ele[28][12] != ele[28][34];
    ele[28][12] != ele[28][35];
    ele[28][12] != ele[29][12];
    ele[28][12] != ele[29][13];
    ele[28][12] != ele[29][14];
    ele[28][12] != ele[29][15];
    ele[28][12] != ele[29][16];
    ele[28][12] != ele[29][17];
    ele[28][12] != ele[30][12];
    ele[28][12] != ele[31][12];
    ele[28][12] != ele[32][12];
    ele[28][12] != ele[33][12];
    ele[28][12] != ele[34][12];
    ele[28][12] != ele[35][12];
    ele[28][13] != ele[28][14];
    ele[28][13] != ele[28][15];
    ele[28][13] != ele[28][16];
    ele[28][13] != ele[28][17];
    ele[28][13] != ele[28][18];
    ele[28][13] != ele[28][19];
    ele[28][13] != ele[28][20];
    ele[28][13] != ele[28][21];
    ele[28][13] != ele[28][22];
    ele[28][13] != ele[28][23];
    ele[28][13] != ele[28][24];
    ele[28][13] != ele[28][25];
    ele[28][13] != ele[28][26];
    ele[28][13] != ele[28][27];
    ele[28][13] != ele[28][28];
    ele[28][13] != ele[28][29];
    ele[28][13] != ele[28][30];
    ele[28][13] != ele[28][31];
    ele[28][13] != ele[28][32];
    ele[28][13] != ele[28][33];
    ele[28][13] != ele[28][34];
    ele[28][13] != ele[28][35];
    ele[28][13] != ele[29][12];
    ele[28][13] != ele[29][13];
    ele[28][13] != ele[29][14];
    ele[28][13] != ele[29][15];
    ele[28][13] != ele[29][16];
    ele[28][13] != ele[29][17];
    ele[28][13] != ele[30][13];
    ele[28][13] != ele[31][13];
    ele[28][13] != ele[32][13];
    ele[28][13] != ele[33][13];
    ele[28][13] != ele[34][13];
    ele[28][13] != ele[35][13];
    ele[28][14] != ele[28][15];
    ele[28][14] != ele[28][16];
    ele[28][14] != ele[28][17];
    ele[28][14] != ele[28][18];
    ele[28][14] != ele[28][19];
    ele[28][14] != ele[28][20];
    ele[28][14] != ele[28][21];
    ele[28][14] != ele[28][22];
    ele[28][14] != ele[28][23];
    ele[28][14] != ele[28][24];
    ele[28][14] != ele[28][25];
    ele[28][14] != ele[28][26];
    ele[28][14] != ele[28][27];
    ele[28][14] != ele[28][28];
    ele[28][14] != ele[28][29];
    ele[28][14] != ele[28][30];
    ele[28][14] != ele[28][31];
    ele[28][14] != ele[28][32];
    ele[28][14] != ele[28][33];
    ele[28][14] != ele[28][34];
    ele[28][14] != ele[28][35];
    ele[28][14] != ele[29][12];
    ele[28][14] != ele[29][13];
    ele[28][14] != ele[29][14];
    ele[28][14] != ele[29][15];
    ele[28][14] != ele[29][16];
    ele[28][14] != ele[29][17];
    ele[28][14] != ele[30][14];
    ele[28][14] != ele[31][14];
    ele[28][14] != ele[32][14];
    ele[28][14] != ele[33][14];
    ele[28][14] != ele[34][14];
    ele[28][14] != ele[35][14];
    ele[28][15] != ele[28][16];
    ele[28][15] != ele[28][17];
    ele[28][15] != ele[28][18];
    ele[28][15] != ele[28][19];
    ele[28][15] != ele[28][20];
    ele[28][15] != ele[28][21];
    ele[28][15] != ele[28][22];
    ele[28][15] != ele[28][23];
    ele[28][15] != ele[28][24];
    ele[28][15] != ele[28][25];
    ele[28][15] != ele[28][26];
    ele[28][15] != ele[28][27];
    ele[28][15] != ele[28][28];
    ele[28][15] != ele[28][29];
    ele[28][15] != ele[28][30];
    ele[28][15] != ele[28][31];
    ele[28][15] != ele[28][32];
    ele[28][15] != ele[28][33];
    ele[28][15] != ele[28][34];
    ele[28][15] != ele[28][35];
    ele[28][15] != ele[29][12];
    ele[28][15] != ele[29][13];
    ele[28][15] != ele[29][14];
    ele[28][15] != ele[29][15];
    ele[28][15] != ele[29][16];
    ele[28][15] != ele[29][17];
    ele[28][15] != ele[30][15];
    ele[28][15] != ele[31][15];
    ele[28][15] != ele[32][15];
    ele[28][15] != ele[33][15];
    ele[28][15] != ele[34][15];
    ele[28][15] != ele[35][15];
    ele[28][16] != ele[28][17];
    ele[28][16] != ele[28][18];
    ele[28][16] != ele[28][19];
    ele[28][16] != ele[28][20];
    ele[28][16] != ele[28][21];
    ele[28][16] != ele[28][22];
    ele[28][16] != ele[28][23];
    ele[28][16] != ele[28][24];
    ele[28][16] != ele[28][25];
    ele[28][16] != ele[28][26];
    ele[28][16] != ele[28][27];
    ele[28][16] != ele[28][28];
    ele[28][16] != ele[28][29];
    ele[28][16] != ele[28][30];
    ele[28][16] != ele[28][31];
    ele[28][16] != ele[28][32];
    ele[28][16] != ele[28][33];
    ele[28][16] != ele[28][34];
    ele[28][16] != ele[28][35];
    ele[28][16] != ele[29][12];
    ele[28][16] != ele[29][13];
    ele[28][16] != ele[29][14];
    ele[28][16] != ele[29][15];
    ele[28][16] != ele[29][16];
    ele[28][16] != ele[29][17];
    ele[28][16] != ele[30][16];
    ele[28][16] != ele[31][16];
    ele[28][16] != ele[32][16];
    ele[28][16] != ele[33][16];
    ele[28][16] != ele[34][16];
    ele[28][16] != ele[35][16];
    ele[28][17] != ele[28][18];
    ele[28][17] != ele[28][19];
    ele[28][17] != ele[28][20];
    ele[28][17] != ele[28][21];
    ele[28][17] != ele[28][22];
    ele[28][17] != ele[28][23];
    ele[28][17] != ele[28][24];
    ele[28][17] != ele[28][25];
    ele[28][17] != ele[28][26];
    ele[28][17] != ele[28][27];
    ele[28][17] != ele[28][28];
    ele[28][17] != ele[28][29];
    ele[28][17] != ele[28][30];
    ele[28][17] != ele[28][31];
    ele[28][17] != ele[28][32];
    ele[28][17] != ele[28][33];
    ele[28][17] != ele[28][34];
    ele[28][17] != ele[28][35];
    ele[28][17] != ele[29][12];
    ele[28][17] != ele[29][13];
    ele[28][17] != ele[29][14];
    ele[28][17] != ele[29][15];
    ele[28][17] != ele[29][16];
    ele[28][17] != ele[29][17];
    ele[28][17] != ele[30][17];
    ele[28][17] != ele[31][17];
    ele[28][17] != ele[32][17];
    ele[28][17] != ele[33][17];
    ele[28][17] != ele[34][17];
    ele[28][17] != ele[35][17];
    ele[28][18] != ele[28][19];
    ele[28][18] != ele[28][20];
    ele[28][18] != ele[28][21];
    ele[28][18] != ele[28][22];
    ele[28][18] != ele[28][23];
    ele[28][18] != ele[28][24];
    ele[28][18] != ele[28][25];
    ele[28][18] != ele[28][26];
    ele[28][18] != ele[28][27];
    ele[28][18] != ele[28][28];
    ele[28][18] != ele[28][29];
    ele[28][18] != ele[28][30];
    ele[28][18] != ele[28][31];
    ele[28][18] != ele[28][32];
    ele[28][18] != ele[28][33];
    ele[28][18] != ele[28][34];
    ele[28][18] != ele[28][35];
    ele[28][18] != ele[29][18];
    ele[28][18] != ele[29][19];
    ele[28][18] != ele[29][20];
    ele[28][18] != ele[29][21];
    ele[28][18] != ele[29][22];
    ele[28][18] != ele[29][23];
    ele[28][18] != ele[30][18];
    ele[28][18] != ele[31][18];
    ele[28][18] != ele[32][18];
    ele[28][18] != ele[33][18];
    ele[28][18] != ele[34][18];
    ele[28][18] != ele[35][18];
    ele[28][19] != ele[28][20];
    ele[28][19] != ele[28][21];
    ele[28][19] != ele[28][22];
    ele[28][19] != ele[28][23];
    ele[28][19] != ele[28][24];
    ele[28][19] != ele[28][25];
    ele[28][19] != ele[28][26];
    ele[28][19] != ele[28][27];
    ele[28][19] != ele[28][28];
    ele[28][19] != ele[28][29];
    ele[28][19] != ele[28][30];
    ele[28][19] != ele[28][31];
    ele[28][19] != ele[28][32];
    ele[28][19] != ele[28][33];
    ele[28][19] != ele[28][34];
    ele[28][19] != ele[28][35];
    ele[28][19] != ele[29][18];
    ele[28][19] != ele[29][19];
    ele[28][19] != ele[29][20];
    ele[28][19] != ele[29][21];
    ele[28][19] != ele[29][22];
    ele[28][19] != ele[29][23];
    ele[28][19] != ele[30][19];
    ele[28][19] != ele[31][19];
    ele[28][19] != ele[32][19];
    ele[28][19] != ele[33][19];
    ele[28][19] != ele[34][19];
    ele[28][19] != ele[35][19];
    ele[28][2] != ele[28][10];
    ele[28][2] != ele[28][11];
    ele[28][2] != ele[28][12];
    ele[28][2] != ele[28][13];
    ele[28][2] != ele[28][14];
    ele[28][2] != ele[28][15];
    ele[28][2] != ele[28][16];
    ele[28][2] != ele[28][17];
    ele[28][2] != ele[28][18];
    ele[28][2] != ele[28][19];
    ele[28][2] != ele[28][20];
    ele[28][2] != ele[28][21];
    ele[28][2] != ele[28][22];
    ele[28][2] != ele[28][23];
    ele[28][2] != ele[28][24];
    ele[28][2] != ele[28][25];
    ele[28][2] != ele[28][26];
    ele[28][2] != ele[28][27];
    ele[28][2] != ele[28][28];
    ele[28][2] != ele[28][29];
    ele[28][2] != ele[28][3];
    ele[28][2] != ele[28][30];
    ele[28][2] != ele[28][31];
    ele[28][2] != ele[28][32];
    ele[28][2] != ele[28][33];
    ele[28][2] != ele[28][34];
    ele[28][2] != ele[28][35];
    ele[28][2] != ele[28][4];
    ele[28][2] != ele[28][5];
    ele[28][2] != ele[28][6];
    ele[28][2] != ele[28][7];
    ele[28][2] != ele[28][8];
    ele[28][2] != ele[28][9];
    ele[28][2] != ele[29][0];
    ele[28][2] != ele[29][1];
    ele[28][2] != ele[29][2];
    ele[28][2] != ele[29][3];
    ele[28][2] != ele[29][4];
    ele[28][2] != ele[29][5];
    ele[28][2] != ele[30][2];
    ele[28][2] != ele[31][2];
    ele[28][2] != ele[32][2];
    ele[28][2] != ele[33][2];
    ele[28][2] != ele[34][2];
    ele[28][2] != ele[35][2];
    ele[28][20] != ele[28][21];
    ele[28][20] != ele[28][22];
    ele[28][20] != ele[28][23];
    ele[28][20] != ele[28][24];
    ele[28][20] != ele[28][25];
    ele[28][20] != ele[28][26];
    ele[28][20] != ele[28][27];
    ele[28][20] != ele[28][28];
    ele[28][20] != ele[28][29];
    ele[28][20] != ele[28][30];
    ele[28][20] != ele[28][31];
    ele[28][20] != ele[28][32];
    ele[28][20] != ele[28][33];
    ele[28][20] != ele[28][34];
    ele[28][20] != ele[28][35];
    ele[28][20] != ele[29][18];
    ele[28][20] != ele[29][19];
    ele[28][20] != ele[29][20];
    ele[28][20] != ele[29][21];
    ele[28][20] != ele[29][22];
    ele[28][20] != ele[29][23];
    ele[28][20] != ele[30][20];
    ele[28][20] != ele[31][20];
    ele[28][20] != ele[32][20];
    ele[28][20] != ele[33][20];
    ele[28][20] != ele[34][20];
    ele[28][20] != ele[35][20];
    ele[28][21] != ele[28][22];
    ele[28][21] != ele[28][23];
    ele[28][21] != ele[28][24];
    ele[28][21] != ele[28][25];
    ele[28][21] != ele[28][26];
    ele[28][21] != ele[28][27];
    ele[28][21] != ele[28][28];
    ele[28][21] != ele[28][29];
    ele[28][21] != ele[28][30];
    ele[28][21] != ele[28][31];
    ele[28][21] != ele[28][32];
    ele[28][21] != ele[28][33];
    ele[28][21] != ele[28][34];
    ele[28][21] != ele[28][35];
    ele[28][21] != ele[29][18];
    ele[28][21] != ele[29][19];
    ele[28][21] != ele[29][20];
    ele[28][21] != ele[29][21];
    ele[28][21] != ele[29][22];
    ele[28][21] != ele[29][23];
    ele[28][21] != ele[30][21];
    ele[28][21] != ele[31][21];
    ele[28][21] != ele[32][21];
    ele[28][21] != ele[33][21];
    ele[28][21] != ele[34][21];
    ele[28][21] != ele[35][21];
    ele[28][22] != ele[28][23];
    ele[28][22] != ele[28][24];
    ele[28][22] != ele[28][25];
    ele[28][22] != ele[28][26];
    ele[28][22] != ele[28][27];
    ele[28][22] != ele[28][28];
    ele[28][22] != ele[28][29];
    ele[28][22] != ele[28][30];
    ele[28][22] != ele[28][31];
    ele[28][22] != ele[28][32];
    ele[28][22] != ele[28][33];
    ele[28][22] != ele[28][34];
    ele[28][22] != ele[28][35];
    ele[28][22] != ele[29][18];
    ele[28][22] != ele[29][19];
    ele[28][22] != ele[29][20];
    ele[28][22] != ele[29][21];
    ele[28][22] != ele[29][22];
    ele[28][22] != ele[29][23];
    ele[28][22] != ele[30][22];
    ele[28][22] != ele[31][22];
    ele[28][22] != ele[32][22];
    ele[28][22] != ele[33][22];
    ele[28][22] != ele[34][22];
    ele[28][22] != ele[35][22];
    ele[28][23] != ele[28][24];
    ele[28][23] != ele[28][25];
    ele[28][23] != ele[28][26];
    ele[28][23] != ele[28][27];
    ele[28][23] != ele[28][28];
    ele[28][23] != ele[28][29];
    ele[28][23] != ele[28][30];
    ele[28][23] != ele[28][31];
    ele[28][23] != ele[28][32];
    ele[28][23] != ele[28][33];
    ele[28][23] != ele[28][34];
    ele[28][23] != ele[28][35];
    ele[28][23] != ele[29][18];
    ele[28][23] != ele[29][19];
    ele[28][23] != ele[29][20];
    ele[28][23] != ele[29][21];
    ele[28][23] != ele[29][22];
    ele[28][23] != ele[29][23];
    ele[28][23] != ele[30][23];
    ele[28][23] != ele[31][23];
    ele[28][23] != ele[32][23];
    ele[28][23] != ele[33][23];
    ele[28][23] != ele[34][23];
    ele[28][23] != ele[35][23];
    ele[28][24] != ele[28][25];
    ele[28][24] != ele[28][26];
    ele[28][24] != ele[28][27];
    ele[28][24] != ele[28][28];
    ele[28][24] != ele[28][29];
    ele[28][24] != ele[28][30];
    ele[28][24] != ele[28][31];
    ele[28][24] != ele[28][32];
    ele[28][24] != ele[28][33];
    ele[28][24] != ele[28][34];
    ele[28][24] != ele[28][35];
    ele[28][24] != ele[29][24];
    ele[28][24] != ele[29][25];
    ele[28][24] != ele[29][26];
    ele[28][24] != ele[29][27];
    ele[28][24] != ele[29][28];
    ele[28][24] != ele[29][29];
    ele[28][24] != ele[30][24];
    ele[28][24] != ele[31][24];
    ele[28][24] != ele[32][24];
    ele[28][24] != ele[33][24];
    ele[28][24] != ele[34][24];
    ele[28][24] != ele[35][24];
    ele[28][25] != ele[28][26];
    ele[28][25] != ele[28][27];
    ele[28][25] != ele[28][28];
    ele[28][25] != ele[28][29];
    ele[28][25] != ele[28][30];
    ele[28][25] != ele[28][31];
    ele[28][25] != ele[28][32];
    ele[28][25] != ele[28][33];
    ele[28][25] != ele[28][34];
    ele[28][25] != ele[28][35];
    ele[28][25] != ele[29][24];
    ele[28][25] != ele[29][25];
    ele[28][25] != ele[29][26];
    ele[28][25] != ele[29][27];
    ele[28][25] != ele[29][28];
    ele[28][25] != ele[29][29];
    ele[28][25] != ele[30][25];
    ele[28][25] != ele[31][25];
    ele[28][25] != ele[32][25];
    ele[28][25] != ele[33][25];
    ele[28][25] != ele[34][25];
    ele[28][25] != ele[35][25];
    ele[28][26] != ele[28][27];
    ele[28][26] != ele[28][28];
    ele[28][26] != ele[28][29];
    ele[28][26] != ele[28][30];
    ele[28][26] != ele[28][31];
    ele[28][26] != ele[28][32];
    ele[28][26] != ele[28][33];
    ele[28][26] != ele[28][34];
    ele[28][26] != ele[28][35];
    ele[28][26] != ele[29][24];
    ele[28][26] != ele[29][25];
    ele[28][26] != ele[29][26];
    ele[28][26] != ele[29][27];
    ele[28][26] != ele[29][28];
    ele[28][26] != ele[29][29];
    ele[28][26] != ele[30][26];
    ele[28][26] != ele[31][26];
    ele[28][26] != ele[32][26];
    ele[28][26] != ele[33][26];
    ele[28][26] != ele[34][26];
    ele[28][26] != ele[35][26];
    ele[28][27] != ele[28][28];
    ele[28][27] != ele[28][29];
    ele[28][27] != ele[28][30];
    ele[28][27] != ele[28][31];
    ele[28][27] != ele[28][32];
    ele[28][27] != ele[28][33];
    ele[28][27] != ele[28][34];
    ele[28][27] != ele[28][35];
    ele[28][27] != ele[29][24];
    ele[28][27] != ele[29][25];
    ele[28][27] != ele[29][26];
    ele[28][27] != ele[29][27];
    ele[28][27] != ele[29][28];
    ele[28][27] != ele[29][29];
    ele[28][27] != ele[30][27];
    ele[28][27] != ele[31][27];
    ele[28][27] != ele[32][27];
    ele[28][27] != ele[33][27];
    ele[28][27] != ele[34][27];
    ele[28][27] != ele[35][27];
    ele[28][28] != ele[28][29];
    ele[28][28] != ele[28][30];
    ele[28][28] != ele[28][31];
    ele[28][28] != ele[28][32];
    ele[28][28] != ele[28][33];
    ele[28][28] != ele[28][34];
    ele[28][28] != ele[28][35];
    ele[28][28] != ele[29][24];
    ele[28][28] != ele[29][25];
    ele[28][28] != ele[29][26];
    ele[28][28] != ele[29][27];
    ele[28][28] != ele[29][28];
    ele[28][28] != ele[29][29];
    ele[28][28] != ele[30][28];
    ele[28][28] != ele[31][28];
    ele[28][28] != ele[32][28];
    ele[28][28] != ele[33][28];
    ele[28][28] != ele[34][28];
    ele[28][28] != ele[35][28];
    ele[28][29] != ele[28][30];
    ele[28][29] != ele[28][31];
    ele[28][29] != ele[28][32];
    ele[28][29] != ele[28][33];
    ele[28][29] != ele[28][34];
    ele[28][29] != ele[28][35];
    ele[28][29] != ele[29][24];
    ele[28][29] != ele[29][25];
    ele[28][29] != ele[29][26];
    ele[28][29] != ele[29][27];
    ele[28][29] != ele[29][28];
    ele[28][29] != ele[29][29];
    ele[28][29] != ele[30][29];
    ele[28][29] != ele[31][29];
    ele[28][29] != ele[32][29];
    ele[28][29] != ele[33][29];
    ele[28][29] != ele[34][29];
    ele[28][29] != ele[35][29];
    ele[28][3] != ele[28][10];
    ele[28][3] != ele[28][11];
    ele[28][3] != ele[28][12];
    ele[28][3] != ele[28][13];
    ele[28][3] != ele[28][14];
    ele[28][3] != ele[28][15];
    ele[28][3] != ele[28][16];
    ele[28][3] != ele[28][17];
    ele[28][3] != ele[28][18];
    ele[28][3] != ele[28][19];
    ele[28][3] != ele[28][20];
    ele[28][3] != ele[28][21];
    ele[28][3] != ele[28][22];
    ele[28][3] != ele[28][23];
    ele[28][3] != ele[28][24];
    ele[28][3] != ele[28][25];
    ele[28][3] != ele[28][26];
    ele[28][3] != ele[28][27];
    ele[28][3] != ele[28][28];
    ele[28][3] != ele[28][29];
    ele[28][3] != ele[28][30];
    ele[28][3] != ele[28][31];
    ele[28][3] != ele[28][32];
    ele[28][3] != ele[28][33];
    ele[28][3] != ele[28][34];
    ele[28][3] != ele[28][35];
    ele[28][3] != ele[28][4];
    ele[28][3] != ele[28][5];
    ele[28][3] != ele[28][6];
    ele[28][3] != ele[28][7];
    ele[28][3] != ele[28][8];
    ele[28][3] != ele[28][9];
    ele[28][3] != ele[29][0];
    ele[28][3] != ele[29][1];
    ele[28][3] != ele[29][2];
    ele[28][3] != ele[29][3];
    ele[28][3] != ele[29][4];
    ele[28][3] != ele[29][5];
    ele[28][3] != ele[30][3];
    ele[28][3] != ele[31][3];
    ele[28][3] != ele[32][3];
    ele[28][3] != ele[33][3];
    ele[28][3] != ele[34][3];
    ele[28][3] != ele[35][3];
    ele[28][30] != ele[28][31];
    ele[28][30] != ele[28][32];
    ele[28][30] != ele[28][33];
    ele[28][30] != ele[28][34];
    ele[28][30] != ele[28][35];
    ele[28][30] != ele[29][30];
    ele[28][30] != ele[29][31];
    ele[28][30] != ele[29][32];
    ele[28][30] != ele[29][33];
    ele[28][30] != ele[29][34];
    ele[28][30] != ele[29][35];
    ele[28][30] != ele[30][30];
    ele[28][30] != ele[31][30];
    ele[28][30] != ele[32][30];
    ele[28][30] != ele[33][30];
    ele[28][30] != ele[34][30];
    ele[28][30] != ele[35][30];
    ele[28][31] != ele[28][32];
    ele[28][31] != ele[28][33];
    ele[28][31] != ele[28][34];
    ele[28][31] != ele[28][35];
    ele[28][31] != ele[29][30];
    ele[28][31] != ele[29][31];
    ele[28][31] != ele[29][32];
    ele[28][31] != ele[29][33];
    ele[28][31] != ele[29][34];
    ele[28][31] != ele[29][35];
    ele[28][31] != ele[30][31];
    ele[28][31] != ele[31][31];
    ele[28][31] != ele[32][31];
    ele[28][31] != ele[33][31];
    ele[28][31] != ele[34][31];
    ele[28][31] != ele[35][31];
    ele[28][32] != ele[28][33];
    ele[28][32] != ele[28][34];
    ele[28][32] != ele[28][35];
    ele[28][32] != ele[29][30];
    ele[28][32] != ele[29][31];
    ele[28][32] != ele[29][32];
    ele[28][32] != ele[29][33];
    ele[28][32] != ele[29][34];
    ele[28][32] != ele[29][35];
    ele[28][32] != ele[30][32];
    ele[28][32] != ele[31][32];
    ele[28][32] != ele[32][32];
    ele[28][32] != ele[33][32];
    ele[28][32] != ele[34][32];
    ele[28][32] != ele[35][32];
    ele[28][33] != ele[28][34];
    ele[28][33] != ele[28][35];
    ele[28][33] != ele[29][30];
    ele[28][33] != ele[29][31];
    ele[28][33] != ele[29][32];
    ele[28][33] != ele[29][33];
    ele[28][33] != ele[29][34];
    ele[28][33] != ele[29][35];
    ele[28][33] != ele[30][33];
    ele[28][33] != ele[31][33];
    ele[28][33] != ele[32][33];
    ele[28][33] != ele[33][33];
    ele[28][33] != ele[34][33];
    ele[28][33] != ele[35][33];
    ele[28][34] != ele[28][35];
    ele[28][34] != ele[29][30];
    ele[28][34] != ele[29][31];
    ele[28][34] != ele[29][32];
    ele[28][34] != ele[29][33];
    ele[28][34] != ele[29][34];
    ele[28][34] != ele[29][35];
    ele[28][34] != ele[30][34];
    ele[28][34] != ele[31][34];
    ele[28][34] != ele[32][34];
    ele[28][34] != ele[33][34];
    ele[28][34] != ele[34][34];
    ele[28][34] != ele[35][34];
    ele[28][35] != ele[29][30];
    ele[28][35] != ele[29][31];
    ele[28][35] != ele[29][32];
    ele[28][35] != ele[29][33];
    ele[28][35] != ele[29][34];
    ele[28][35] != ele[29][35];
    ele[28][35] != ele[30][35];
    ele[28][35] != ele[31][35];
    ele[28][35] != ele[32][35];
    ele[28][35] != ele[33][35];
    ele[28][35] != ele[34][35];
    ele[28][35] != ele[35][35];
    ele[28][4] != ele[28][10];
    ele[28][4] != ele[28][11];
    ele[28][4] != ele[28][12];
    ele[28][4] != ele[28][13];
    ele[28][4] != ele[28][14];
    ele[28][4] != ele[28][15];
    ele[28][4] != ele[28][16];
    ele[28][4] != ele[28][17];
    ele[28][4] != ele[28][18];
    ele[28][4] != ele[28][19];
    ele[28][4] != ele[28][20];
    ele[28][4] != ele[28][21];
    ele[28][4] != ele[28][22];
    ele[28][4] != ele[28][23];
    ele[28][4] != ele[28][24];
    ele[28][4] != ele[28][25];
    ele[28][4] != ele[28][26];
    ele[28][4] != ele[28][27];
    ele[28][4] != ele[28][28];
    ele[28][4] != ele[28][29];
    ele[28][4] != ele[28][30];
    ele[28][4] != ele[28][31];
    ele[28][4] != ele[28][32];
    ele[28][4] != ele[28][33];
    ele[28][4] != ele[28][34];
    ele[28][4] != ele[28][35];
    ele[28][4] != ele[28][5];
    ele[28][4] != ele[28][6];
    ele[28][4] != ele[28][7];
    ele[28][4] != ele[28][8];
    ele[28][4] != ele[28][9];
    ele[28][4] != ele[29][0];
    ele[28][4] != ele[29][1];
    ele[28][4] != ele[29][2];
    ele[28][4] != ele[29][3];
    ele[28][4] != ele[29][4];
    ele[28][4] != ele[29][5];
    ele[28][4] != ele[30][4];
    ele[28][4] != ele[31][4];
    ele[28][4] != ele[32][4];
    ele[28][4] != ele[33][4];
    ele[28][4] != ele[34][4];
    ele[28][4] != ele[35][4];
    ele[28][5] != ele[28][10];
    ele[28][5] != ele[28][11];
    ele[28][5] != ele[28][12];
    ele[28][5] != ele[28][13];
    ele[28][5] != ele[28][14];
    ele[28][5] != ele[28][15];
    ele[28][5] != ele[28][16];
    ele[28][5] != ele[28][17];
    ele[28][5] != ele[28][18];
    ele[28][5] != ele[28][19];
    ele[28][5] != ele[28][20];
    ele[28][5] != ele[28][21];
    ele[28][5] != ele[28][22];
    ele[28][5] != ele[28][23];
    ele[28][5] != ele[28][24];
    ele[28][5] != ele[28][25];
    ele[28][5] != ele[28][26];
    ele[28][5] != ele[28][27];
    ele[28][5] != ele[28][28];
    ele[28][5] != ele[28][29];
    ele[28][5] != ele[28][30];
    ele[28][5] != ele[28][31];
    ele[28][5] != ele[28][32];
    ele[28][5] != ele[28][33];
    ele[28][5] != ele[28][34];
    ele[28][5] != ele[28][35];
    ele[28][5] != ele[28][6];
    ele[28][5] != ele[28][7];
    ele[28][5] != ele[28][8];
    ele[28][5] != ele[28][9];
    ele[28][5] != ele[29][0];
    ele[28][5] != ele[29][1];
    ele[28][5] != ele[29][2];
    ele[28][5] != ele[29][3];
    ele[28][5] != ele[29][4];
    ele[28][5] != ele[29][5];
    ele[28][5] != ele[30][5];
    ele[28][5] != ele[31][5];
    ele[28][5] != ele[32][5];
    ele[28][5] != ele[33][5];
    ele[28][5] != ele[34][5];
    ele[28][5] != ele[35][5];
    ele[28][6] != ele[28][10];
    ele[28][6] != ele[28][11];
    ele[28][6] != ele[28][12];
    ele[28][6] != ele[28][13];
    ele[28][6] != ele[28][14];
    ele[28][6] != ele[28][15];
    ele[28][6] != ele[28][16];
    ele[28][6] != ele[28][17];
    ele[28][6] != ele[28][18];
    ele[28][6] != ele[28][19];
    ele[28][6] != ele[28][20];
    ele[28][6] != ele[28][21];
    ele[28][6] != ele[28][22];
    ele[28][6] != ele[28][23];
    ele[28][6] != ele[28][24];
    ele[28][6] != ele[28][25];
    ele[28][6] != ele[28][26];
    ele[28][6] != ele[28][27];
    ele[28][6] != ele[28][28];
    ele[28][6] != ele[28][29];
    ele[28][6] != ele[28][30];
    ele[28][6] != ele[28][31];
    ele[28][6] != ele[28][32];
    ele[28][6] != ele[28][33];
    ele[28][6] != ele[28][34];
    ele[28][6] != ele[28][35];
    ele[28][6] != ele[28][7];
    ele[28][6] != ele[28][8];
    ele[28][6] != ele[28][9];
    ele[28][6] != ele[29][10];
    ele[28][6] != ele[29][11];
    ele[28][6] != ele[29][6];
    ele[28][6] != ele[29][7];
    ele[28][6] != ele[29][8];
    ele[28][6] != ele[29][9];
    ele[28][6] != ele[30][6];
    ele[28][6] != ele[31][6];
    ele[28][6] != ele[32][6];
    ele[28][6] != ele[33][6];
    ele[28][6] != ele[34][6];
    ele[28][6] != ele[35][6];
    ele[28][7] != ele[28][10];
    ele[28][7] != ele[28][11];
    ele[28][7] != ele[28][12];
    ele[28][7] != ele[28][13];
    ele[28][7] != ele[28][14];
    ele[28][7] != ele[28][15];
    ele[28][7] != ele[28][16];
    ele[28][7] != ele[28][17];
    ele[28][7] != ele[28][18];
    ele[28][7] != ele[28][19];
    ele[28][7] != ele[28][20];
    ele[28][7] != ele[28][21];
    ele[28][7] != ele[28][22];
    ele[28][7] != ele[28][23];
    ele[28][7] != ele[28][24];
    ele[28][7] != ele[28][25];
    ele[28][7] != ele[28][26];
    ele[28][7] != ele[28][27];
    ele[28][7] != ele[28][28];
    ele[28][7] != ele[28][29];
    ele[28][7] != ele[28][30];
    ele[28][7] != ele[28][31];
    ele[28][7] != ele[28][32];
    ele[28][7] != ele[28][33];
    ele[28][7] != ele[28][34];
    ele[28][7] != ele[28][35];
    ele[28][7] != ele[28][8];
    ele[28][7] != ele[28][9];
    ele[28][7] != ele[29][10];
    ele[28][7] != ele[29][11];
    ele[28][7] != ele[29][6];
    ele[28][7] != ele[29][7];
    ele[28][7] != ele[29][8];
    ele[28][7] != ele[29][9];
    ele[28][7] != ele[30][7];
    ele[28][7] != ele[31][7];
    ele[28][7] != ele[32][7];
    ele[28][7] != ele[33][7];
    ele[28][7] != ele[34][7];
    ele[28][7] != ele[35][7];
    ele[28][8] != ele[28][10];
    ele[28][8] != ele[28][11];
    ele[28][8] != ele[28][12];
    ele[28][8] != ele[28][13];
    ele[28][8] != ele[28][14];
    ele[28][8] != ele[28][15];
    ele[28][8] != ele[28][16];
    ele[28][8] != ele[28][17];
    ele[28][8] != ele[28][18];
    ele[28][8] != ele[28][19];
    ele[28][8] != ele[28][20];
    ele[28][8] != ele[28][21];
    ele[28][8] != ele[28][22];
    ele[28][8] != ele[28][23];
    ele[28][8] != ele[28][24];
    ele[28][8] != ele[28][25];
    ele[28][8] != ele[28][26];
    ele[28][8] != ele[28][27];
    ele[28][8] != ele[28][28];
    ele[28][8] != ele[28][29];
    ele[28][8] != ele[28][30];
    ele[28][8] != ele[28][31];
    ele[28][8] != ele[28][32];
    ele[28][8] != ele[28][33];
    ele[28][8] != ele[28][34];
    ele[28][8] != ele[28][35];
    ele[28][8] != ele[28][9];
    ele[28][8] != ele[29][10];
    ele[28][8] != ele[29][11];
    ele[28][8] != ele[29][6];
    ele[28][8] != ele[29][7];
    ele[28][8] != ele[29][8];
    ele[28][8] != ele[29][9];
    ele[28][8] != ele[30][8];
    ele[28][8] != ele[31][8];
    ele[28][8] != ele[32][8];
    ele[28][8] != ele[33][8];
    ele[28][8] != ele[34][8];
    ele[28][8] != ele[35][8];
    ele[28][9] != ele[28][10];
    ele[28][9] != ele[28][11];
    ele[28][9] != ele[28][12];
    ele[28][9] != ele[28][13];
    ele[28][9] != ele[28][14];
    ele[28][9] != ele[28][15];
    ele[28][9] != ele[28][16];
    ele[28][9] != ele[28][17];
    ele[28][9] != ele[28][18];
    ele[28][9] != ele[28][19];
    ele[28][9] != ele[28][20];
    ele[28][9] != ele[28][21];
    ele[28][9] != ele[28][22];
    ele[28][9] != ele[28][23];
    ele[28][9] != ele[28][24];
    ele[28][9] != ele[28][25];
    ele[28][9] != ele[28][26];
    ele[28][9] != ele[28][27];
    ele[28][9] != ele[28][28];
    ele[28][9] != ele[28][29];
    ele[28][9] != ele[28][30];
    ele[28][9] != ele[28][31];
    ele[28][9] != ele[28][32];
    ele[28][9] != ele[28][33];
    ele[28][9] != ele[28][34];
    ele[28][9] != ele[28][35];
    ele[28][9] != ele[29][10];
    ele[28][9] != ele[29][11];
    ele[28][9] != ele[29][6];
    ele[28][9] != ele[29][7];
    ele[28][9] != ele[29][8];
    ele[28][9] != ele[29][9];
    ele[28][9] != ele[30][9];
    ele[28][9] != ele[31][9];
    ele[28][9] != ele[32][9];
    ele[28][9] != ele[33][9];
    ele[28][9] != ele[34][9];
    ele[28][9] != ele[35][9];
    ele[29][0] != ele[29][1];
    ele[29][0] != ele[29][10];
    ele[29][0] != ele[29][11];
    ele[29][0] != ele[29][12];
    ele[29][0] != ele[29][13];
    ele[29][0] != ele[29][14];
    ele[29][0] != ele[29][15];
    ele[29][0] != ele[29][16];
    ele[29][0] != ele[29][17];
    ele[29][0] != ele[29][18];
    ele[29][0] != ele[29][19];
    ele[29][0] != ele[29][2];
    ele[29][0] != ele[29][20];
    ele[29][0] != ele[29][21];
    ele[29][0] != ele[29][22];
    ele[29][0] != ele[29][23];
    ele[29][0] != ele[29][24];
    ele[29][0] != ele[29][25];
    ele[29][0] != ele[29][26];
    ele[29][0] != ele[29][27];
    ele[29][0] != ele[29][28];
    ele[29][0] != ele[29][29];
    ele[29][0] != ele[29][3];
    ele[29][0] != ele[29][30];
    ele[29][0] != ele[29][31];
    ele[29][0] != ele[29][32];
    ele[29][0] != ele[29][33];
    ele[29][0] != ele[29][34];
    ele[29][0] != ele[29][35];
    ele[29][0] != ele[29][4];
    ele[29][0] != ele[29][5];
    ele[29][0] != ele[29][6];
    ele[29][0] != ele[29][7];
    ele[29][0] != ele[29][8];
    ele[29][0] != ele[29][9];
    ele[29][0] != ele[30][0];
    ele[29][0] != ele[31][0];
    ele[29][0] != ele[32][0];
    ele[29][0] != ele[33][0];
    ele[29][0] != ele[34][0];
    ele[29][0] != ele[35][0];
    ele[29][1] != ele[29][10];
    ele[29][1] != ele[29][11];
    ele[29][1] != ele[29][12];
    ele[29][1] != ele[29][13];
    ele[29][1] != ele[29][14];
    ele[29][1] != ele[29][15];
    ele[29][1] != ele[29][16];
    ele[29][1] != ele[29][17];
    ele[29][1] != ele[29][18];
    ele[29][1] != ele[29][19];
    ele[29][1] != ele[29][2];
    ele[29][1] != ele[29][20];
    ele[29][1] != ele[29][21];
    ele[29][1] != ele[29][22];
    ele[29][1] != ele[29][23];
    ele[29][1] != ele[29][24];
    ele[29][1] != ele[29][25];
    ele[29][1] != ele[29][26];
    ele[29][1] != ele[29][27];
    ele[29][1] != ele[29][28];
    ele[29][1] != ele[29][29];
    ele[29][1] != ele[29][3];
    ele[29][1] != ele[29][30];
    ele[29][1] != ele[29][31];
    ele[29][1] != ele[29][32];
    ele[29][1] != ele[29][33];
    ele[29][1] != ele[29][34];
    ele[29][1] != ele[29][35];
    ele[29][1] != ele[29][4];
    ele[29][1] != ele[29][5];
    ele[29][1] != ele[29][6];
    ele[29][1] != ele[29][7];
    ele[29][1] != ele[29][8];
    ele[29][1] != ele[29][9];
    ele[29][1] != ele[30][1];
    ele[29][1] != ele[31][1];
    ele[29][1] != ele[32][1];
    ele[29][1] != ele[33][1];
    ele[29][1] != ele[34][1];
    ele[29][1] != ele[35][1];
    ele[29][10] != ele[29][11];
    ele[29][10] != ele[29][12];
    ele[29][10] != ele[29][13];
    ele[29][10] != ele[29][14];
    ele[29][10] != ele[29][15];
    ele[29][10] != ele[29][16];
    ele[29][10] != ele[29][17];
    ele[29][10] != ele[29][18];
    ele[29][10] != ele[29][19];
    ele[29][10] != ele[29][20];
    ele[29][10] != ele[29][21];
    ele[29][10] != ele[29][22];
    ele[29][10] != ele[29][23];
    ele[29][10] != ele[29][24];
    ele[29][10] != ele[29][25];
    ele[29][10] != ele[29][26];
    ele[29][10] != ele[29][27];
    ele[29][10] != ele[29][28];
    ele[29][10] != ele[29][29];
    ele[29][10] != ele[29][30];
    ele[29][10] != ele[29][31];
    ele[29][10] != ele[29][32];
    ele[29][10] != ele[29][33];
    ele[29][10] != ele[29][34];
    ele[29][10] != ele[29][35];
    ele[29][10] != ele[30][10];
    ele[29][10] != ele[31][10];
    ele[29][10] != ele[32][10];
    ele[29][10] != ele[33][10];
    ele[29][10] != ele[34][10];
    ele[29][10] != ele[35][10];
    ele[29][11] != ele[29][12];
    ele[29][11] != ele[29][13];
    ele[29][11] != ele[29][14];
    ele[29][11] != ele[29][15];
    ele[29][11] != ele[29][16];
    ele[29][11] != ele[29][17];
    ele[29][11] != ele[29][18];
    ele[29][11] != ele[29][19];
    ele[29][11] != ele[29][20];
    ele[29][11] != ele[29][21];
    ele[29][11] != ele[29][22];
    ele[29][11] != ele[29][23];
    ele[29][11] != ele[29][24];
    ele[29][11] != ele[29][25];
    ele[29][11] != ele[29][26];
    ele[29][11] != ele[29][27];
    ele[29][11] != ele[29][28];
    ele[29][11] != ele[29][29];
    ele[29][11] != ele[29][30];
    ele[29][11] != ele[29][31];
    ele[29][11] != ele[29][32];
    ele[29][11] != ele[29][33];
    ele[29][11] != ele[29][34];
    ele[29][11] != ele[29][35];
    ele[29][11] != ele[30][11];
    ele[29][11] != ele[31][11];
    ele[29][11] != ele[32][11];
    ele[29][11] != ele[33][11];
    ele[29][11] != ele[34][11];
    ele[29][11] != ele[35][11];
    ele[29][12] != ele[29][13];
    ele[29][12] != ele[29][14];
    ele[29][12] != ele[29][15];
    ele[29][12] != ele[29][16];
    ele[29][12] != ele[29][17];
    ele[29][12] != ele[29][18];
    ele[29][12] != ele[29][19];
    ele[29][12] != ele[29][20];
    ele[29][12] != ele[29][21];
    ele[29][12] != ele[29][22];
    ele[29][12] != ele[29][23];
    ele[29][12] != ele[29][24];
    ele[29][12] != ele[29][25];
    ele[29][12] != ele[29][26];
    ele[29][12] != ele[29][27];
    ele[29][12] != ele[29][28];
    ele[29][12] != ele[29][29];
    ele[29][12] != ele[29][30];
    ele[29][12] != ele[29][31];
    ele[29][12] != ele[29][32];
    ele[29][12] != ele[29][33];
    ele[29][12] != ele[29][34];
    ele[29][12] != ele[29][35];
    ele[29][12] != ele[30][12];
    ele[29][12] != ele[31][12];
    ele[29][12] != ele[32][12];
    ele[29][12] != ele[33][12];
    ele[29][12] != ele[34][12];
    ele[29][12] != ele[35][12];
    ele[29][13] != ele[29][14];
    ele[29][13] != ele[29][15];
    ele[29][13] != ele[29][16];
    ele[29][13] != ele[29][17];
    ele[29][13] != ele[29][18];
    ele[29][13] != ele[29][19];
    ele[29][13] != ele[29][20];
    ele[29][13] != ele[29][21];
    ele[29][13] != ele[29][22];
    ele[29][13] != ele[29][23];
    ele[29][13] != ele[29][24];
    ele[29][13] != ele[29][25];
    ele[29][13] != ele[29][26];
    ele[29][13] != ele[29][27];
    ele[29][13] != ele[29][28];
    ele[29][13] != ele[29][29];
    ele[29][13] != ele[29][30];
    ele[29][13] != ele[29][31];
    ele[29][13] != ele[29][32];
    ele[29][13] != ele[29][33];
    ele[29][13] != ele[29][34];
    ele[29][13] != ele[29][35];
    ele[29][13] != ele[30][13];
    ele[29][13] != ele[31][13];
    ele[29][13] != ele[32][13];
    ele[29][13] != ele[33][13];
    ele[29][13] != ele[34][13];
    ele[29][13] != ele[35][13];
    ele[29][14] != ele[29][15];
    ele[29][14] != ele[29][16];
    ele[29][14] != ele[29][17];
    ele[29][14] != ele[29][18];
    ele[29][14] != ele[29][19];
    ele[29][14] != ele[29][20];
    ele[29][14] != ele[29][21];
    ele[29][14] != ele[29][22];
    ele[29][14] != ele[29][23];
    ele[29][14] != ele[29][24];
    ele[29][14] != ele[29][25];
    ele[29][14] != ele[29][26];
    ele[29][14] != ele[29][27];
    ele[29][14] != ele[29][28];
    ele[29][14] != ele[29][29];
    ele[29][14] != ele[29][30];
    ele[29][14] != ele[29][31];
    ele[29][14] != ele[29][32];
    ele[29][14] != ele[29][33];
    ele[29][14] != ele[29][34];
    ele[29][14] != ele[29][35];
    ele[29][14] != ele[30][14];
    ele[29][14] != ele[31][14];
    ele[29][14] != ele[32][14];
    ele[29][14] != ele[33][14];
    ele[29][14] != ele[34][14];
    ele[29][14] != ele[35][14];
    ele[29][15] != ele[29][16];
    ele[29][15] != ele[29][17];
    ele[29][15] != ele[29][18];
    ele[29][15] != ele[29][19];
    ele[29][15] != ele[29][20];
    ele[29][15] != ele[29][21];
    ele[29][15] != ele[29][22];
    ele[29][15] != ele[29][23];
    ele[29][15] != ele[29][24];
    ele[29][15] != ele[29][25];
    ele[29][15] != ele[29][26];
    ele[29][15] != ele[29][27];
    ele[29][15] != ele[29][28];
    ele[29][15] != ele[29][29];
    ele[29][15] != ele[29][30];
    ele[29][15] != ele[29][31];
    ele[29][15] != ele[29][32];
    ele[29][15] != ele[29][33];
    ele[29][15] != ele[29][34];
    ele[29][15] != ele[29][35];
    ele[29][15] != ele[30][15];
    ele[29][15] != ele[31][15];
    ele[29][15] != ele[32][15];
    ele[29][15] != ele[33][15];
    ele[29][15] != ele[34][15];
    ele[29][15] != ele[35][15];
    ele[29][16] != ele[29][17];
    ele[29][16] != ele[29][18];
    ele[29][16] != ele[29][19];
    ele[29][16] != ele[29][20];
    ele[29][16] != ele[29][21];
    ele[29][16] != ele[29][22];
    ele[29][16] != ele[29][23];
    ele[29][16] != ele[29][24];
    ele[29][16] != ele[29][25];
    ele[29][16] != ele[29][26];
    ele[29][16] != ele[29][27];
    ele[29][16] != ele[29][28];
    ele[29][16] != ele[29][29];
    ele[29][16] != ele[29][30];
    ele[29][16] != ele[29][31];
    ele[29][16] != ele[29][32];
    ele[29][16] != ele[29][33];
    ele[29][16] != ele[29][34];
    ele[29][16] != ele[29][35];
    ele[29][16] != ele[30][16];
    ele[29][16] != ele[31][16];
    ele[29][16] != ele[32][16];
    ele[29][16] != ele[33][16];
    ele[29][16] != ele[34][16];
    ele[29][16] != ele[35][16];
    ele[29][17] != ele[29][18];
    ele[29][17] != ele[29][19];
    ele[29][17] != ele[29][20];
    ele[29][17] != ele[29][21];
    ele[29][17] != ele[29][22];
    ele[29][17] != ele[29][23];
    ele[29][17] != ele[29][24];
    ele[29][17] != ele[29][25];
    ele[29][17] != ele[29][26];
    ele[29][17] != ele[29][27];
    ele[29][17] != ele[29][28];
    ele[29][17] != ele[29][29];
    ele[29][17] != ele[29][30];
    ele[29][17] != ele[29][31];
    ele[29][17] != ele[29][32];
    ele[29][17] != ele[29][33];
    ele[29][17] != ele[29][34];
    ele[29][17] != ele[29][35];
    ele[29][17] != ele[30][17];
    ele[29][17] != ele[31][17];
    ele[29][17] != ele[32][17];
    ele[29][17] != ele[33][17];
    ele[29][17] != ele[34][17];
    ele[29][17] != ele[35][17];
    ele[29][18] != ele[29][19];
    ele[29][18] != ele[29][20];
    ele[29][18] != ele[29][21];
    ele[29][18] != ele[29][22];
    ele[29][18] != ele[29][23];
    ele[29][18] != ele[29][24];
    ele[29][18] != ele[29][25];
    ele[29][18] != ele[29][26];
    ele[29][18] != ele[29][27];
    ele[29][18] != ele[29][28];
    ele[29][18] != ele[29][29];
    ele[29][18] != ele[29][30];
    ele[29][18] != ele[29][31];
    ele[29][18] != ele[29][32];
    ele[29][18] != ele[29][33];
    ele[29][18] != ele[29][34];
    ele[29][18] != ele[29][35];
    ele[29][18] != ele[30][18];
    ele[29][18] != ele[31][18];
    ele[29][18] != ele[32][18];
    ele[29][18] != ele[33][18];
    ele[29][18] != ele[34][18];
    ele[29][18] != ele[35][18];
    ele[29][19] != ele[29][20];
    ele[29][19] != ele[29][21];
    ele[29][19] != ele[29][22];
    ele[29][19] != ele[29][23];
    ele[29][19] != ele[29][24];
    ele[29][19] != ele[29][25];
    ele[29][19] != ele[29][26];
    ele[29][19] != ele[29][27];
    ele[29][19] != ele[29][28];
    ele[29][19] != ele[29][29];
    ele[29][19] != ele[29][30];
    ele[29][19] != ele[29][31];
    ele[29][19] != ele[29][32];
    ele[29][19] != ele[29][33];
    ele[29][19] != ele[29][34];
    ele[29][19] != ele[29][35];
    ele[29][19] != ele[30][19];
    ele[29][19] != ele[31][19];
    ele[29][19] != ele[32][19];
    ele[29][19] != ele[33][19];
    ele[29][19] != ele[34][19];
    ele[29][19] != ele[35][19];
    ele[29][2] != ele[29][10];
    ele[29][2] != ele[29][11];
    ele[29][2] != ele[29][12];
    ele[29][2] != ele[29][13];
    ele[29][2] != ele[29][14];
    ele[29][2] != ele[29][15];
    ele[29][2] != ele[29][16];
    ele[29][2] != ele[29][17];
    ele[29][2] != ele[29][18];
    ele[29][2] != ele[29][19];
    ele[29][2] != ele[29][20];
    ele[29][2] != ele[29][21];
    ele[29][2] != ele[29][22];
    ele[29][2] != ele[29][23];
    ele[29][2] != ele[29][24];
    ele[29][2] != ele[29][25];
    ele[29][2] != ele[29][26];
    ele[29][2] != ele[29][27];
    ele[29][2] != ele[29][28];
    ele[29][2] != ele[29][29];
    ele[29][2] != ele[29][3];
    ele[29][2] != ele[29][30];
    ele[29][2] != ele[29][31];
    ele[29][2] != ele[29][32];
    ele[29][2] != ele[29][33];
    ele[29][2] != ele[29][34];
    ele[29][2] != ele[29][35];
    ele[29][2] != ele[29][4];
    ele[29][2] != ele[29][5];
    ele[29][2] != ele[29][6];
    ele[29][2] != ele[29][7];
    ele[29][2] != ele[29][8];
    ele[29][2] != ele[29][9];
    ele[29][2] != ele[30][2];
    ele[29][2] != ele[31][2];
    ele[29][2] != ele[32][2];
    ele[29][2] != ele[33][2];
    ele[29][2] != ele[34][2];
    ele[29][2] != ele[35][2];
    ele[29][20] != ele[29][21];
    ele[29][20] != ele[29][22];
    ele[29][20] != ele[29][23];
    ele[29][20] != ele[29][24];
    ele[29][20] != ele[29][25];
    ele[29][20] != ele[29][26];
    ele[29][20] != ele[29][27];
    ele[29][20] != ele[29][28];
    ele[29][20] != ele[29][29];
    ele[29][20] != ele[29][30];
    ele[29][20] != ele[29][31];
    ele[29][20] != ele[29][32];
    ele[29][20] != ele[29][33];
    ele[29][20] != ele[29][34];
    ele[29][20] != ele[29][35];
    ele[29][20] != ele[30][20];
    ele[29][20] != ele[31][20];
    ele[29][20] != ele[32][20];
    ele[29][20] != ele[33][20];
    ele[29][20] != ele[34][20];
    ele[29][20] != ele[35][20];
    ele[29][21] != ele[29][22];
    ele[29][21] != ele[29][23];
    ele[29][21] != ele[29][24];
    ele[29][21] != ele[29][25];
    ele[29][21] != ele[29][26];
    ele[29][21] != ele[29][27];
    ele[29][21] != ele[29][28];
    ele[29][21] != ele[29][29];
    ele[29][21] != ele[29][30];
    ele[29][21] != ele[29][31];
    ele[29][21] != ele[29][32];
    ele[29][21] != ele[29][33];
    ele[29][21] != ele[29][34];
    ele[29][21] != ele[29][35];
    ele[29][21] != ele[30][21];
    ele[29][21] != ele[31][21];
    ele[29][21] != ele[32][21];
    ele[29][21] != ele[33][21];
    ele[29][21] != ele[34][21];
    ele[29][21] != ele[35][21];
    ele[29][22] != ele[29][23];
    ele[29][22] != ele[29][24];
    ele[29][22] != ele[29][25];
    ele[29][22] != ele[29][26];
    ele[29][22] != ele[29][27];
    ele[29][22] != ele[29][28];
    ele[29][22] != ele[29][29];
    ele[29][22] != ele[29][30];
    ele[29][22] != ele[29][31];
    ele[29][22] != ele[29][32];
    ele[29][22] != ele[29][33];
    ele[29][22] != ele[29][34];
    ele[29][22] != ele[29][35];
    ele[29][22] != ele[30][22];
    ele[29][22] != ele[31][22];
    ele[29][22] != ele[32][22];
    ele[29][22] != ele[33][22];
    ele[29][22] != ele[34][22];
    ele[29][22] != ele[35][22];
    ele[29][23] != ele[29][24];
    ele[29][23] != ele[29][25];
    ele[29][23] != ele[29][26];
    ele[29][23] != ele[29][27];
    ele[29][23] != ele[29][28];
    ele[29][23] != ele[29][29];
    ele[29][23] != ele[29][30];
    ele[29][23] != ele[29][31];
    ele[29][23] != ele[29][32];
    ele[29][23] != ele[29][33];
    ele[29][23] != ele[29][34];
    ele[29][23] != ele[29][35];
    ele[29][23] != ele[30][23];
    ele[29][23] != ele[31][23];
    ele[29][23] != ele[32][23];
    ele[29][23] != ele[33][23];
    ele[29][23] != ele[34][23];
    ele[29][23] != ele[35][23];
    ele[29][24] != ele[29][25];
    ele[29][24] != ele[29][26];
    ele[29][24] != ele[29][27];
    ele[29][24] != ele[29][28];
    ele[29][24] != ele[29][29];
    ele[29][24] != ele[29][30];
    ele[29][24] != ele[29][31];
    ele[29][24] != ele[29][32];
    ele[29][24] != ele[29][33];
    ele[29][24] != ele[29][34];
    ele[29][24] != ele[29][35];
    ele[29][24] != ele[30][24];
    ele[29][24] != ele[31][24];
    ele[29][24] != ele[32][24];
    ele[29][24] != ele[33][24];
    ele[29][24] != ele[34][24];
    ele[29][24] != ele[35][24];
    ele[29][25] != ele[29][26];
    ele[29][25] != ele[29][27];
    ele[29][25] != ele[29][28];
    ele[29][25] != ele[29][29];
    ele[29][25] != ele[29][30];
    ele[29][25] != ele[29][31];
    ele[29][25] != ele[29][32];
    ele[29][25] != ele[29][33];
    ele[29][25] != ele[29][34];
    ele[29][25] != ele[29][35];
    ele[29][25] != ele[30][25];
    ele[29][25] != ele[31][25];
    ele[29][25] != ele[32][25];
    ele[29][25] != ele[33][25];
    ele[29][25] != ele[34][25];
    ele[29][25] != ele[35][25];
    ele[29][26] != ele[29][27];
    ele[29][26] != ele[29][28];
    ele[29][26] != ele[29][29];
    ele[29][26] != ele[29][30];
    ele[29][26] != ele[29][31];
    ele[29][26] != ele[29][32];
    ele[29][26] != ele[29][33];
    ele[29][26] != ele[29][34];
    ele[29][26] != ele[29][35];
    ele[29][26] != ele[30][26];
    ele[29][26] != ele[31][26];
    ele[29][26] != ele[32][26];
    ele[29][26] != ele[33][26];
    ele[29][26] != ele[34][26];
    ele[29][26] != ele[35][26];
    ele[29][27] != ele[29][28];
    ele[29][27] != ele[29][29];
    ele[29][27] != ele[29][30];
    ele[29][27] != ele[29][31];
    ele[29][27] != ele[29][32];
    ele[29][27] != ele[29][33];
    ele[29][27] != ele[29][34];
    ele[29][27] != ele[29][35];
    ele[29][27] != ele[30][27];
    ele[29][27] != ele[31][27];
    ele[29][27] != ele[32][27];
    ele[29][27] != ele[33][27];
    ele[29][27] != ele[34][27];
    ele[29][27] != ele[35][27];
    ele[29][28] != ele[29][29];
    ele[29][28] != ele[29][30];
    ele[29][28] != ele[29][31];
    ele[29][28] != ele[29][32];
    ele[29][28] != ele[29][33];
    ele[29][28] != ele[29][34];
    ele[29][28] != ele[29][35];
    ele[29][28] != ele[30][28];
    ele[29][28] != ele[31][28];
    ele[29][28] != ele[32][28];
    ele[29][28] != ele[33][28];
    ele[29][28] != ele[34][28];
    ele[29][28] != ele[35][28];
    ele[29][29] != ele[29][30];
    ele[29][29] != ele[29][31];
    ele[29][29] != ele[29][32];
    ele[29][29] != ele[29][33];
    ele[29][29] != ele[29][34];
    ele[29][29] != ele[29][35];
    ele[29][29] != ele[30][29];
    ele[29][29] != ele[31][29];
    ele[29][29] != ele[32][29];
    ele[29][29] != ele[33][29];
    ele[29][29] != ele[34][29];
    ele[29][29] != ele[35][29];
    ele[29][3] != ele[29][10];
    ele[29][3] != ele[29][11];
    ele[29][3] != ele[29][12];
    ele[29][3] != ele[29][13];
    ele[29][3] != ele[29][14];
    ele[29][3] != ele[29][15];
    ele[29][3] != ele[29][16];
    ele[29][3] != ele[29][17];
    ele[29][3] != ele[29][18];
    ele[29][3] != ele[29][19];
    ele[29][3] != ele[29][20];
    ele[29][3] != ele[29][21];
    ele[29][3] != ele[29][22];
    ele[29][3] != ele[29][23];
    ele[29][3] != ele[29][24];
    ele[29][3] != ele[29][25];
    ele[29][3] != ele[29][26];
    ele[29][3] != ele[29][27];
    ele[29][3] != ele[29][28];
    ele[29][3] != ele[29][29];
    ele[29][3] != ele[29][30];
    ele[29][3] != ele[29][31];
    ele[29][3] != ele[29][32];
    ele[29][3] != ele[29][33];
    ele[29][3] != ele[29][34];
    ele[29][3] != ele[29][35];
    ele[29][3] != ele[29][4];
    ele[29][3] != ele[29][5];
    ele[29][3] != ele[29][6];
    ele[29][3] != ele[29][7];
    ele[29][3] != ele[29][8];
    ele[29][3] != ele[29][9];
    ele[29][3] != ele[30][3];
    ele[29][3] != ele[31][3];
    ele[29][3] != ele[32][3];
    ele[29][3] != ele[33][3];
    ele[29][3] != ele[34][3];
    ele[29][3] != ele[35][3];
    ele[29][30] != ele[29][31];
    ele[29][30] != ele[29][32];
    ele[29][30] != ele[29][33];
    ele[29][30] != ele[29][34];
    ele[29][30] != ele[29][35];
    ele[29][30] != ele[30][30];
    ele[29][30] != ele[31][30];
    ele[29][30] != ele[32][30];
    ele[29][30] != ele[33][30];
    ele[29][30] != ele[34][30];
    ele[29][30] != ele[35][30];
    ele[29][31] != ele[29][32];
    ele[29][31] != ele[29][33];
    ele[29][31] != ele[29][34];
    ele[29][31] != ele[29][35];
    ele[29][31] != ele[30][31];
    ele[29][31] != ele[31][31];
    ele[29][31] != ele[32][31];
    ele[29][31] != ele[33][31];
    ele[29][31] != ele[34][31];
    ele[29][31] != ele[35][31];
    ele[29][32] != ele[29][33];
    ele[29][32] != ele[29][34];
    ele[29][32] != ele[29][35];
    ele[29][32] != ele[30][32];
    ele[29][32] != ele[31][32];
    ele[29][32] != ele[32][32];
    ele[29][32] != ele[33][32];
    ele[29][32] != ele[34][32];
    ele[29][32] != ele[35][32];
    ele[29][33] != ele[29][34];
    ele[29][33] != ele[29][35];
    ele[29][33] != ele[30][33];
    ele[29][33] != ele[31][33];
    ele[29][33] != ele[32][33];
    ele[29][33] != ele[33][33];
    ele[29][33] != ele[34][33];
    ele[29][33] != ele[35][33];
    ele[29][34] != ele[29][35];
    ele[29][34] != ele[30][34];
    ele[29][34] != ele[31][34];
    ele[29][34] != ele[32][34];
    ele[29][34] != ele[33][34];
    ele[29][34] != ele[34][34];
    ele[29][34] != ele[35][34];
    ele[29][35] != ele[30][35];
    ele[29][35] != ele[31][35];
    ele[29][35] != ele[32][35];
    ele[29][35] != ele[33][35];
    ele[29][35] != ele[34][35];
    ele[29][35] != ele[35][35];
    ele[29][4] != ele[29][10];
    ele[29][4] != ele[29][11];
    ele[29][4] != ele[29][12];
    ele[29][4] != ele[29][13];
    ele[29][4] != ele[29][14];
    ele[29][4] != ele[29][15];
    ele[29][4] != ele[29][16];
    ele[29][4] != ele[29][17];
    ele[29][4] != ele[29][18];
    ele[29][4] != ele[29][19];
    ele[29][4] != ele[29][20];
    ele[29][4] != ele[29][21];
    ele[29][4] != ele[29][22];
    ele[29][4] != ele[29][23];
    ele[29][4] != ele[29][24];
    ele[29][4] != ele[29][25];
    ele[29][4] != ele[29][26];
    ele[29][4] != ele[29][27];
    ele[29][4] != ele[29][28];
    ele[29][4] != ele[29][29];
    ele[29][4] != ele[29][30];
    ele[29][4] != ele[29][31];
    ele[29][4] != ele[29][32];
    ele[29][4] != ele[29][33];
    ele[29][4] != ele[29][34];
    ele[29][4] != ele[29][35];
    ele[29][4] != ele[29][5];
    ele[29][4] != ele[29][6];
    ele[29][4] != ele[29][7];
    ele[29][4] != ele[29][8];
    ele[29][4] != ele[29][9];
    ele[29][4] != ele[30][4];
    ele[29][4] != ele[31][4];
    ele[29][4] != ele[32][4];
    ele[29][4] != ele[33][4];
    ele[29][4] != ele[34][4];
    ele[29][4] != ele[35][4];
    ele[29][5] != ele[29][10];
    ele[29][5] != ele[29][11];
    ele[29][5] != ele[29][12];
    ele[29][5] != ele[29][13];
    ele[29][5] != ele[29][14];
    ele[29][5] != ele[29][15];
    ele[29][5] != ele[29][16];
    ele[29][5] != ele[29][17];
    ele[29][5] != ele[29][18];
    ele[29][5] != ele[29][19];
    ele[29][5] != ele[29][20];
    ele[29][5] != ele[29][21];
    ele[29][5] != ele[29][22];
    ele[29][5] != ele[29][23];
    ele[29][5] != ele[29][24];
    ele[29][5] != ele[29][25];
    ele[29][5] != ele[29][26];
    ele[29][5] != ele[29][27];
    ele[29][5] != ele[29][28];
    ele[29][5] != ele[29][29];
    ele[29][5] != ele[29][30];
    ele[29][5] != ele[29][31];
    ele[29][5] != ele[29][32];
    ele[29][5] != ele[29][33];
    ele[29][5] != ele[29][34];
    ele[29][5] != ele[29][35];
    ele[29][5] != ele[29][6];
    ele[29][5] != ele[29][7];
    ele[29][5] != ele[29][8];
    ele[29][5] != ele[29][9];
    ele[29][5] != ele[30][5];
    ele[29][5] != ele[31][5];
    ele[29][5] != ele[32][5];
    ele[29][5] != ele[33][5];
    ele[29][5] != ele[34][5];
    ele[29][5] != ele[35][5];
    ele[29][6] != ele[29][10];
    ele[29][6] != ele[29][11];
    ele[29][6] != ele[29][12];
    ele[29][6] != ele[29][13];
    ele[29][6] != ele[29][14];
    ele[29][6] != ele[29][15];
    ele[29][6] != ele[29][16];
    ele[29][6] != ele[29][17];
    ele[29][6] != ele[29][18];
    ele[29][6] != ele[29][19];
    ele[29][6] != ele[29][20];
    ele[29][6] != ele[29][21];
    ele[29][6] != ele[29][22];
    ele[29][6] != ele[29][23];
    ele[29][6] != ele[29][24];
    ele[29][6] != ele[29][25];
    ele[29][6] != ele[29][26];
    ele[29][6] != ele[29][27];
    ele[29][6] != ele[29][28];
    ele[29][6] != ele[29][29];
    ele[29][6] != ele[29][30];
    ele[29][6] != ele[29][31];
    ele[29][6] != ele[29][32];
    ele[29][6] != ele[29][33];
    ele[29][6] != ele[29][34];
    ele[29][6] != ele[29][35];
    ele[29][6] != ele[29][7];
    ele[29][6] != ele[29][8];
    ele[29][6] != ele[29][9];
    ele[29][6] != ele[30][6];
    ele[29][6] != ele[31][6];
    ele[29][6] != ele[32][6];
    ele[29][6] != ele[33][6];
    ele[29][6] != ele[34][6];
    ele[29][6] != ele[35][6];
    ele[29][7] != ele[29][10];
    ele[29][7] != ele[29][11];
    ele[29][7] != ele[29][12];
    ele[29][7] != ele[29][13];
    ele[29][7] != ele[29][14];
    ele[29][7] != ele[29][15];
    ele[29][7] != ele[29][16];
    ele[29][7] != ele[29][17];
    ele[29][7] != ele[29][18];
    ele[29][7] != ele[29][19];
    ele[29][7] != ele[29][20];
    ele[29][7] != ele[29][21];
    ele[29][7] != ele[29][22];
    ele[29][7] != ele[29][23];
    ele[29][7] != ele[29][24];
    ele[29][7] != ele[29][25];
    ele[29][7] != ele[29][26];
    ele[29][7] != ele[29][27];
    ele[29][7] != ele[29][28];
    ele[29][7] != ele[29][29];
    ele[29][7] != ele[29][30];
    ele[29][7] != ele[29][31];
    ele[29][7] != ele[29][32];
    ele[29][7] != ele[29][33];
    ele[29][7] != ele[29][34];
    ele[29][7] != ele[29][35];
    ele[29][7] != ele[29][8];
    ele[29][7] != ele[29][9];
    ele[29][7] != ele[30][7];
    ele[29][7] != ele[31][7];
    ele[29][7] != ele[32][7];
    ele[29][7] != ele[33][7];
    ele[29][7] != ele[34][7];
    ele[29][7] != ele[35][7];
    ele[29][8] != ele[29][10];
    ele[29][8] != ele[29][11];
    ele[29][8] != ele[29][12];
    ele[29][8] != ele[29][13];
    ele[29][8] != ele[29][14];
    ele[29][8] != ele[29][15];
    ele[29][8] != ele[29][16];
    ele[29][8] != ele[29][17];
    ele[29][8] != ele[29][18];
    ele[29][8] != ele[29][19];
    ele[29][8] != ele[29][20];
    ele[29][8] != ele[29][21];
    ele[29][8] != ele[29][22];
    ele[29][8] != ele[29][23];
    ele[29][8] != ele[29][24];
    ele[29][8] != ele[29][25];
    ele[29][8] != ele[29][26];
    ele[29][8] != ele[29][27];
    ele[29][8] != ele[29][28];
    ele[29][8] != ele[29][29];
    ele[29][8] != ele[29][30];
    ele[29][8] != ele[29][31];
    ele[29][8] != ele[29][32];
    ele[29][8] != ele[29][33];
    ele[29][8] != ele[29][34];
    ele[29][8] != ele[29][35];
    ele[29][8] != ele[29][9];
    ele[29][8] != ele[30][8];
    ele[29][8] != ele[31][8];
    ele[29][8] != ele[32][8];
    ele[29][8] != ele[33][8];
    ele[29][8] != ele[34][8];
    ele[29][8] != ele[35][8];
    ele[29][9] != ele[29][10];
    ele[29][9] != ele[29][11];
    ele[29][9] != ele[29][12];
    ele[29][9] != ele[29][13];
    ele[29][9] != ele[29][14];
    ele[29][9] != ele[29][15];
    ele[29][9] != ele[29][16];
    ele[29][9] != ele[29][17];
    ele[29][9] != ele[29][18];
    ele[29][9] != ele[29][19];
    ele[29][9] != ele[29][20];
    ele[29][9] != ele[29][21];
    ele[29][9] != ele[29][22];
    ele[29][9] != ele[29][23];
    ele[29][9] != ele[29][24];
    ele[29][9] != ele[29][25];
    ele[29][9] != ele[29][26];
    ele[29][9] != ele[29][27];
    ele[29][9] != ele[29][28];
    ele[29][9] != ele[29][29];
    ele[29][9] != ele[29][30];
    ele[29][9] != ele[29][31];
    ele[29][9] != ele[29][32];
    ele[29][9] != ele[29][33];
    ele[29][9] != ele[29][34];
    ele[29][9] != ele[29][35];
    ele[29][9] != ele[30][9];
    ele[29][9] != ele[31][9];
    ele[29][9] != ele[32][9];
    ele[29][9] != ele[33][9];
    ele[29][9] != ele[34][9];
    ele[29][9] != ele[35][9];
    ele[3][0] != ele[10][0];
    ele[3][0] != ele[11][0];
    ele[3][0] != ele[12][0];
    ele[3][0] != ele[13][0];
    ele[3][0] != ele[14][0];
    ele[3][0] != ele[15][0];
    ele[3][0] != ele[16][0];
    ele[3][0] != ele[17][0];
    ele[3][0] != ele[18][0];
    ele[3][0] != ele[19][0];
    ele[3][0] != ele[20][0];
    ele[3][0] != ele[21][0];
    ele[3][0] != ele[22][0];
    ele[3][0] != ele[23][0];
    ele[3][0] != ele[24][0];
    ele[3][0] != ele[25][0];
    ele[3][0] != ele[26][0];
    ele[3][0] != ele[27][0];
    ele[3][0] != ele[28][0];
    ele[3][0] != ele[29][0];
    ele[3][0] != ele[3][1];
    ele[3][0] != ele[3][10];
    ele[3][0] != ele[3][11];
    ele[3][0] != ele[3][12];
    ele[3][0] != ele[3][13];
    ele[3][0] != ele[3][14];
    ele[3][0] != ele[3][15];
    ele[3][0] != ele[3][16];
    ele[3][0] != ele[3][17];
    ele[3][0] != ele[3][18];
    ele[3][0] != ele[3][19];
    ele[3][0] != ele[3][2];
    ele[3][0] != ele[3][20];
    ele[3][0] != ele[3][21];
    ele[3][0] != ele[3][22];
    ele[3][0] != ele[3][23];
    ele[3][0] != ele[3][24];
    ele[3][0] != ele[3][25];
    ele[3][0] != ele[3][26];
    ele[3][0] != ele[3][27];
    ele[3][0] != ele[3][28];
    ele[3][0] != ele[3][29];
    ele[3][0] != ele[3][3];
    ele[3][0] != ele[3][30];
    ele[3][0] != ele[3][31];
    ele[3][0] != ele[3][32];
    ele[3][0] != ele[3][33];
    ele[3][0] != ele[3][34];
    ele[3][0] != ele[3][35];
    ele[3][0] != ele[3][4];
    ele[3][0] != ele[3][5];
    ele[3][0] != ele[3][6];
    ele[3][0] != ele[3][7];
    ele[3][0] != ele[3][8];
    ele[3][0] != ele[3][9];
    ele[3][0] != ele[30][0];
    ele[3][0] != ele[31][0];
    ele[3][0] != ele[32][0];
    ele[3][0] != ele[33][0];
    ele[3][0] != ele[34][0];
    ele[3][0] != ele[35][0];
    ele[3][0] != ele[4][0];
    ele[3][0] != ele[4][1];
    ele[3][0] != ele[4][2];
    ele[3][0] != ele[4][3];
    ele[3][0] != ele[4][4];
    ele[3][0] != ele[4][5];
    ele[3][0] != ele[5][0];
    ele[3][0] != ele[5][1];
    ele[3][0] != ele[5][2];
    ele[3][0] != ele[5][3];
    ele[3][0] != ele[5][4];
    ele[3][0] != ele[5][5];
    ele[3][0] != ele[6][0];
    ele[3][0] != ele[7][0];
    ele[3][0] != ele[8][0];
    ele[3][0] != ele[9][0];
    ele[3][1] != ele[10][1];
    ele[3][1] != ele[11][1];
    ele[3][1] != ele[12][1];
    ele[3][1] != ele[13][1];
    ele[3][1] != ele[14][1];
    ele[3][1] != ele[15][1];
    ele[3][1] != ele[16][1];
    ele[3][1] != ele[17][1];
    ele[3][1] != ele[18][1];
    ele[3][1] != ele[19][1];
    ele[3][1] != ele[20][1];
    ele[3][1] != ele[21][1];
    ele[3][1] != ele[22][1];
    ele[3][1] != ele[23][1];
    ele[3][1] != ele[24][1];
    ele[3][1] != ele[25][1];
    ele[3][1] != ele[26][1];
    ele[3][1] != ele[27][1];
    ele[3][1] != ele[28][1];
    ele[3][1] != ele[29][1];
    ele[3][1] != ele[3][10];
    ele[3][1] != ele[3][11];
    ele[3][1] != ele[3][12];
    ele[3][1] != ele[3][13];
    ele[3][1] != ele[3][14];
    ele[3][1] != ele[3][15];
    ele[3][1] != ele[3][16];
    ele[3][1] != ele[3][17];
    ele[3][1] != ele[3][18];
    ele[3][1] != ele[3][19];
    ele[3][1] != ele[3][2];
    ele[3][1] != ele[3][20];
    ele[3][1] != ele[3][21];
    ele[3][1] != ele[3][22];
    ele[3][1] != ele[3][23];
    ele[3][1] != ele[3][24];
    ele[3][1] != ele[3][25];
    ele[3][1] != ele[3][26];
    ele[3][1] != ele[3][27];
    ele[3][1] != ele[3][28];
    ele[3][1] != ele[3][29];
    ele[3][1] != ele[3][3];
    ele[3][1] != ele[3][30];
    ele[3][1] != ele[3][31];
    ele[3][1] != ele[3][32];
    ele[3][1] != ele[3][33];
    ele[3][1] != ele[3][34];
    ele[3][1] != ele[3][35];
    ele[3][1] != ele[3][4];
    ele[3][1] != ele[3][5];
    ele[3][1] != ele[3][6];
    ele[3][1] != ele[3][7];
    ele[3][1] != ele[3][8];
    ele[3][1] != ele[3][9];
    ele[3][1] != ele[30][1];
    ele[3][1] != ele[31][1];
    ele[3][1] != ele[32][1];
    ele[3][1] != ele[33][1];
    ele[3][1] != ele[34][1];
    ele[3][1] != ele[35][1];
    ele[3][1] != ele[4][0];
    ele[3][1] != ele[4][1];
    ele[3][1] != ele[4][2];
    ele[3][1] != ele[4][3];
    ele[3][1] != ele[4][4];
    ele[3][1] != ele[4][5];
    ele[3][1] != ele[5][0];
    ele[3][1] != ele[5][1];
    ele[3][1] != ele[5][2];
    ele[3][1] != ele[5][3];
    ele[3][1] != ele[5][4];
    ele[3][1] != ele[5][5];
    ele[3][1] != ele[6][1];
    ele[3][1] != ele[7][1];
    ele[3][1] != ele[8][1];
    ele[3][1] != ele[9][1];
    ele[3][10] != ele[10][10];
    ele[3][10] != ele[11][10];
    ele[3][10] != ele[12][10];
    ele[3][10] != ele[13][10];
    ele[3][10] != ele[14][10];
    ele[3][10] != ele[15][10];
    ele[3][10] != ele[16][10];
    ele[3][10] != ele[17][10];
    ele[3][10] != ele[18][10];
    ele[3][10] != ele[19][10];
    ele[3][10] != ele[20][10];
    ele[3][10] != ele[21][10];
    ele[3][10] != ele[22][10];
    ele[3][10] != ele[23][10];
    ele[3][10] != ele[24][10];
    ele[3][10] != ele[25][10];
    ele[3][10] != ele[26][10];
    ele[3][10] != ele[27][10];
    ele[3][10] != ele[28][10];
    ele[3][10] != ele[29][10];
    ele[3][10] != ele[3][11];
    ele[3][10] != ele[3][12];
    ele[3][10] != ele[3][13];
    ele[3][10] != ele[3][14];
    ele[3][10] != ele[3][15];
    ele[3][10] != ele[3][16];
    ele[3][10] != ele[3][17];
    ele[3][10] != ele[3][18];
    ele[3][10] != ele[3][19];
    ele[3][10] != ele[3][20];
    ele[3][10] != ele[3][21];
    ele[3][10] != ele[3][22];
    ele[3][10] != ele[3][23];
    ele[3][10] != ele[3][24];
    ele[3][10] != ele[3][25];
    ele[3][10] != ele[3][26];
    ele[3][10] != ele[3][27];
    ele[3][10] != ele[3][28];
    ele[3][10] != ele[3][29];
    ele[3][10] != ele[3][30];
    ele[3][10] != ele[3][31];
    ele[3][10] != ele[3][32];
    ele[3][10] != ele[3][33];
    ele[3][10] != ele[3][34];
    ele[3][10] != ele[3][35];
    ele[3][10] != ele[30][10];
    ele[3][10] != ele[31][10];
    ele[3][10] != ele[32][10];
    ele[3][10] != ele[33][10];
    ele[3][10] != ele[34][10];
    ele[3][10] != ele[35][10];
    ele[3][10] != ele[4][10];
    ele[3][10] != ele[4][11];
    ele[3][10] != ele[4][6];
    ele[3][10] != ele[4][7];
    ele[3][10] != ele[4][8];
    ele[3][10] != ele[4][9];
    ele[3][10] != ele[5][10];
    ele[3][10] != ele[5][11];
    ele[3][10] != ele[5][6];
    ele[3][10] != ele[5][7];
    ele[3][10] != ele[5][8];
    ele[3][10] != ele[5][9];
    ele[3][10] != ele[6][10];
    ele[3][10] != ele[7][10];
    ele[3][10] != ele[8][10];
    ele[3][10] != ele[9][10];
    ele[3][11] != ele[10][11];
    ele[3][11] != ele[11][11];
    ele[3][11] != ele[12][11];
    ele[3][11] != ele[13][11];
    ele[3][11] != ele[14][11];
    ele[3][11] != ele[15][11];
    ele[3][11] != ele[16][11];
    ele[3][11] != ele[17][11];
    ele[3][11] != ele[18][11];
    ele[3][11] != ele[19][11];
    ele[3][11] != ele[20][11];
    ele[3][11] != ele[21][11];
    ele[3][11] != ele[22][11];
    ele[3][11] != ele[23][11];
    ele[3][11] != ele[24][11];
    ele[3][11] != ele[25][11];
    ele[3][11] != ele[26][11];
    ele[3][11] != ele[27][11];
    ele[3][11] != ele[28][11];
    ele[3][11] != ele[29][11];
    ele[3][11] != ele[3][12];
    ele[3][11] != ele[3][13];
    ele[3][11] != ele[3][14];
    ele[3][11] != ele[3][15];
    ele[3][11] != ele[3][16];
    ele[3][11] != ele[3][17];
    ele[3][11] != ele[3][18];
    ele[3][11] != ele[3][19];
    ele[3][11] != ele[3][20];
    ele[3][11] != ele[3][21];
    ele[3][11] != ele[3][22];
    ele[3][11] != ele[3][23];
    ele[3][11] != ele[3][24];
    ele[3][11] != ele[3][25];
    ele[3][11] != ele[3][26];
    ele[3][11] != ele[3][27];
    ele[3][11] != ele[3][28];
    ele[3][11] != ele[3][29];
    ele[3][11] != ele[3][30];
    ele[3][11] != ele[3][31];
    ele[3][11] != ele[3][32];
    ele[3][11] != ele[3][33];
    ele[3][11] != ele[3][34];
    ele[3][11] != ele[3][35];
    ele[3][11] != ele[30][11];
    ele[3][11] != ele[31][11];
    ele[3][11] != ele[32][11];
    ele[3][11] != ele[33][11];
    ele[3][11] != ele[34][11];
    ele[3][11] != ele[35][11];
    ele[3][11] != ele[4][10];
    ele[3][11] != ele[4][11];
    ele[3][11] != ele[4][6];
    ele[3][11] != ele[4][7];
    ele[3][11] != ele[4][8];
    ele[3][11] != ele[4][9];
    ele[3][11] != ele[5][10];
    ele[3][11] != ele[5][11];
    ele[3][11] != ele[5][6];
    ele[3][11] != ele[5][7];
    ele[3][11] != ele[5][8];
    ele[3][11] != ele[5][9];
    ele[3][11] != ele[6][11];
    ele[3][11] != ele[7][11];
    ele[3][11] != ele[8][11];
    ele[3][11] != ele[9][11];
    ele[3][12] != ele[10][12];
    ele[3][12] != ele[11][12];
    ele[3][12] != ele[12][12];
    ele[3][12] != ele[13][12];
    ele[3][12] != ele[14][12];
    ele[3][12] != ele[15][12];
    ele[3][12] != ele[16][12];
    ele[3][12] != ele[17][12];
    ele[3][12] != ele[18][12];
    ele[3][12] != ele[19][12];
    ele[3][12] != ele[20][12];
    ele[3][12] != ele[21][12];
    ele[3][12] != ele[22][12];
    ele[3][12] != ele[23][12];
    ele[3][12] != ele[24][12];
    ele[3][12] != ele[25][12];
    ele[3][12] != ele[26][12];
    ele[3][12] != ele[27][12];
    ele[3][12] != ele[28][12];
    ele[3][12] != ele[29][12];
    ele[3][12] != ele[3][13];
    ele[3][12] != ele[3][14];
    ele[3][12] != ele[3][15];
    ele[3][12] != ele[3][16];
    ele[3][12] != ele[3][17];
    ele[3][12] != ele[3][18];
    ele[3][12] != ele[3][19];
    ele[3][12] != ele[3][20];
    ele[3][12] != ele[3][21];
    ele[3][12] != ele[3][22];
    ele[3][12] != ele[3][23];
    ele[3][12] != ele[3][24];
    ele[3][12] != ele[3][25];
    ele[3][12] != ele[3][26];
    ele[3][12] != ele[3][27];
    ele[3][12] != ele[3][28];
    ele[3][12] != ele[3][29];
    ele[3][12] != ele[3][30];
    ele[3][12] != ele[3][31];
    ele[3][12] != ele[3][32];
    ele[3][12] != ele[3][33];
    ele[3][12] != ele[3][34];
    ele[3][12] != ele[3][35];
    ele[3][12] != ele[30][12];
    ele[3][12] != ele[31][12];
    ele[3][12] != ele[32][12];
    ele[3][12] != ele[33][12];
    ele[3][12] != ele[34][12];
    ele[3][12] != ele[35][12];
    ele[3][12] != ele[4][12];
    ele[3][12] != ele[4][13];
    ele[3][12] != ele[4][14];
    ele[3][12] != ele[4][15];
    ele[3][12] != ele[4][16];
    ele[3][12] != ele[4][17];
    ele[3][12] != ele[5][12];
    ele[3][12] != ele[5][13];
    ele[3][12] != ele[5][14];
    ele[3][12] != ele[5][15];
    ele[3][12] != ele[5][16];
    ele[3][12] != ele[5][17];
    ele[3][12] != ele[6][12];
    ele[3][12] != ele[7][12];
    ele[3][12] != ele[8][12];
    ele[3][12] != ele[9][12];
    ele[3][13] != ele[10][13];
    ele[3][13] != ele[11][13];
    ele[3][13] != ele[12][13];
    ele[3][13] != ele[13][13];
    ele[3][13] != ele[14][13];
    ele[3][13] != ele[15][13];
    ele[3][13] != ele[16][13];
    ele[3][13] != ele[17][13];
    ele[3][13] != ele[18][13];
    ele[3][13] != ele[19][13];
    ele[3][13] != ele[20][13];
    ele[3][13] != ele[21][13];
    ele[3][13] != ele[22][13];
    ele[3][13] != ele[23][13];
    ele[3][13] != ele[24][13];
    ele[3][13] != ele[25][13];
    ele[3][13] != ele[26][13];
    ele[3][13] != ele[27][13];
    ele[3][13] != ele[28][13];
    ele[3][13] != ele[29][13];
    ele[3][13] != ele[3][14];
    ele[3][13] != ele[3][15];
    ele[3][13] != ele[3][16];
    ele[3][13] != ele[3][17];
    ele[3][13] != ele[3][18];
    ele[3][13] != ele[3][19];
    ele[3][13] != ele[3][20];
    ele[3][13] != ele[3][21];
    ele[3][13] != ele[3][22];
    ele[3][13] != ele[3][23];
    ele[3][13] != ele[3][24];
    ele[3][13] != ele[3][25];
    ele[3][13] != ele[3][26];
    ele[3][13] != ele[3][27];
    ele[3][13] != ele[3][28];
    ele[3][13] != ele[3][29];
    ele[3][13] != ele[3][30];
    ele[3][13] != ele[3][31];
    ele[3][13] != ele[3][32];
    ele[3][13] != ele[3][33];
    ele[3][13] != ele[3][34];
    ele[3][13] != ele[3][35];
    ele[3][13] != ele[30][13];
    ele[3][13] != ele[31][13];
    ele[3][13] != ele[32][13];
    ele[3][13] != ele[33][13];
    ele[3][13] != ele[34][13];
    ele[3][13] != ele[35][13];
    ele[3][13] != ele[4][12];
    ele[3][13] != ele[4][13];
    ele[3][13] != ele[4][14];
    ele[3][13] != ele[4][15];
    ele[3][13] != ele[4][16];
    ele[3][13] != ele[4][17];
    ele[3][13] != ele[5][12];
    ele[3][13] != ele[5][13];
    ele[3][13] != ele[5][14];
    ele[3][13] != ele[5][15];
    ele[3][13] != ele[5][16];
    ele[3][13] != ele[5][17];
    ele[3][13] != ele[6][13];
    ele[3][13] != ele[7][13];
    ele[3][13] != ele[8][13];
    ele[3][13] != ele[9][13];
    ele[3][14] != ele[10][14];
    ele[3][14] != ele[11][14];
    ele[3][14] != ele[12][14];
    ele[3][14] != ele[13][14];
    ele[3][14] != ele[14][14];
    ele[3][14] != ele[15][14];
    ele[3][14] != ele[16][14];
    ele[3][14] != ele[17][14];
    ele[3][14] != ele[18][14];
    ele[3][14] != ele[19][14];
    ele[3][14] != ele[20][14];
    ele[3][14] != ele[21][14];
    ele[3][14] != ele[22][14];
    ele[3][14] != ele[23][14];
    ele[3][14] != ele[24][14];
    ele[3][14] != ele[25][14];
    ele[3][14] != ele[26][14];
    ele[3][14] != ele[27][14];
    ele[3][14] != ele[28][14];
    ele[3][14] != ele[29][14];
    ele[3][14] != ele[3][15];
    ele[3][14] != ele[3][16];
    ele[3][14] != ele[3][17];
    ele[3][14] != ele[3][18];
    ele[3][14] != ele[3][19];
    ele[3][14] != ele[3][20];
    ele[3][14] != ele[3][21];
    ele[3][14] != ele[3][22];
    ele[3][14] != ele[3][23];
    ele[3][14] != ele[3][24];
    ele[3][14] != ele[3][25];
    ele[3][14] != ele[3][26];
    ele[3][14] != ele[3][27];
    ele[3][14] != ele[3][28];
    ele[3][14] != ele[3][29];
    ele[3][14] != ele[3][30];
    ele[3][14] != ele[3][31];
    ele[3][14] != ele[3][32];
    ele[3][14] != ele[3][33];
    ele[3][14] != ele[3][34];
    ele[3][14] != ele[3][35];
    ele[3][14] != ele[30][14];
    ele[3][14] != ele[31][14];
    ele[3][14] != ele[32][14];
    ele[3][14] != ele[33][14];
    ele[3][14] != ele[34][14];
    ele[3][14] != ele[35][14];
    ele[3][14] != ele[4][12];
    ele[3][14] != ele[4][13];
    ele[3][14] != ele[4][14];
    ele[3][14] != ele[4][15];
    ele[3][14] != ele[4][16];
    ele[3][14] != ele[4][17];
    ele[3][14] != ele[5][12];
    ele[3][14] != ele[5][13];
    ele[3][14] != ele[5][14];
    ele[3][14] != ele[5][15];
    ele[3][14] != ele[5][16];
    ele[3][14] != ele[5][17];
    ele[3][14] != ele[6][14];
    ele[3][14] != ele[7][14];
    ele[3][14] != ele[8][14];
    ele[3][14] != ele[9][14];
    ele[3][15] != ele[10][15];
    ele[3][15] != ele[11][15];
    ele[3][15] != ele[12][15];
    ele[3][15] != ele[13][15];
    ele[3][15] != ele[14][15];
    ele[3][15] != ele[15][15];
    ele[3][15] != ele[16][15];
    ele[3][15] != ele[17][15];
    ele[3][15] != ele[18][15];
    ele[3][15] != ele[19][15];
    ele[3][15] != ele[20][15];
    ele[3][15] != ele[21][15];
    ele[3][15] != ele[22][15];
    ele[3][15] != ele[23][15];
    ele[3][15] != ele[24][15];
    ele[3][15] != ele[25][15];
    ele[3][15] != ele[26][15];
    ele[3][15] != ele[27][15];
    ele[3][15] != ele[28][15];
    ele[3][15] != ele[29][15];
    ele[3][15] != ele[3][16];
    ele[3][15] != ele[3][17];
    ele[3][15] != ele[3][18];
    ele[3][15] != ele[3][19];
    ele[3][15] != ele[3][20];
    ele[3][15] != ele[3][21];
    ele[3][15] != ele[3][22];
    ele[3][15] != ele[3][23];
    ele[3][15] != ele[3][24];
    ele[3][15] != ele[3][25];
    ele[3][15] != ele[3][26];
    ele[3][15] != ele[3][27];
    ele[3][15] != ele[3][28];
    ele[3][15] != ele[3][29];
    ele[3][15] != ele[3][30];
    ele[3][15] != ele[3][31];
    ele[3][15] != ele[3][32];
    ele[3][15] != ele[3][33];
    ele[3][15] != ele[3][34];
    ele[3][15] != ele[3][35];
    ele[3][15] != ele[30][15];
    ele[3][15] != ele[31][15];
    ele[3][15] != ele[32][15];
    ele[3][15] != ele[33][15];
    ele[3][15] != ele[34][15];
    ele[3][15] != ele[35][15];
    ele[3][15] != ele[4][12];
    ele[3][15] != ele[4][13];
    ele[3][15] != ele[4][14];
    ele[3][15] != ele[4][15];
    ele[3][15] != ele[4][16];
    ele[3][15] != ele[4][17];
    ele[3][15] != ele[5][12];
    ele[3][15] != ele[5][13];
    ele[3][15] != ele[5][14];
    ele[3][15] != ele[5][15];
    ele[3][15] != ele[5][16];
    ele[3][15] != ele[5][17];
    ele[3][15] != ele[6][15];
    ele[3][15] != ele[7][15];
    ele[3][15] != ele[8][15];
    ele[3][15] != ele[9][15];
    ele[3][16] != ele[10][16];
    ele[3][16] != ele[11][16];
    ele[3][16] != ele[12][16];
    ele[3][16] != ele[13][16];
    ele[3][16] != ele[14][16];
    ele[3][16] != ele[15][16];
    ele[3][16] != ele[16][16];
    ele[3][16] != ele[17][16];
    ele[3][16] != ele[18][16];
    ele[3][16] != ele[19][16];
    ele[3][16] != ele[20][16];
    ele[3][16] != ele[21][16];
    ele[3][16] != ele[22][16];
    ele[3][16] != ele[23][16];
    ele[3][16] != ele[24][16];
    ele[3][16] != ele[25][16];
    ele[3][16] != ele[26][16];
    ele[3][16] != ele[27][16];
    ele[3][16] != ele[28][16];
    ele[3][16] != ele[29][16];
    ele[3][16] != ele[3][17];
    ele[3][16] != ele[3][18];
    ele[3][16] != ele[3][19];
    ele[3][16] != ele[3][20];
    ele[3][16] != ele[3][21];
    ele[3][16] != ele[3][22];
    ele[3][16] != ele[3][23];
    ele[3][16] != ele[3][24];
    ele[3][16] != ele[3][25];
    ele[3][16] != ele[3][26];
    ele[3][16] != ele[3][27];
    ele[3][16] != ele[3][28];
    ele[3][16] != ele[3][29];
    ele[3][16] != ele[3][30];
    ele[3][16] != ele[3][31];
    ele[3][16] != ele[3][32];
    ele[3][16] != ele[3][33];
    ele[3][16] != ele[3][34];
    ele[3][16] != ele[3][35];
    ele[3][16] != ele[30][16];
    ele[3][16] != ele[31][16];
    ele[3][16] != ele[32][16];
    ele[3][16] != ele[33][16];
    ele[3][16] != ele[34][16];
    ele[3][16] != ele[35][16];
    ele[3][16] != ele[4][12];
    ele[3][16] != ele[4][13];
    ele[3][16] != ele[4][14];
    ele[3][16] != ele[4][15];
    ele[3][16] != ele[4][16];
    ele[3][16] != ele[4][17];
    ele[3][16] != ele[5][12];
    ele[3][16] != ele[5][13];
    ele[3][16] != ele[5][14];
    ele[3][16] != ele[5][15];
    ele[3][16] != ele[5][16];
    ele[3][16] != ele[5][17];
    ele[3][16] != ele[6][16];
    ele[3][16] != ele[7][16];
    ele[3][16] != ele[8][16];
    ele[3][16] != ele[9][16];
    ele[3][17] != ele[10][17];
    ele[3][17] != ele[11][17];
    ele[3][17] != ele[12][17];
    ele[3][17] != ele[13][17];
    ele[3][17] != ele[14][17];
    ele[3][17] != ele[15][17];
    ele[3][17] != ele[16][17];
    ele[3][17] != ele[17][17];
    ele[3][17] != ele[18][17];
    ele[3][17] != ele[19][17];
    ele[3][17] != ele[20][17];
    ele[3][17] != ele[21][17];
    ele[3][17] != ele[22][17];
    ele[3][17] != ele[23][17];
    ele[3][17] != ele[24][17];
    ele[3][17] != ele[25][17];
    ele[3][17] != ele[26][17];
    ele[3][17] != ele[27][17];
    ele[3][17] != ele[28][17];
    ele[3][17] != ele[29][17];
    ele[3][17] != ele[3][18];
    ele[3][17] != ele[3][19];
    ele[3][17] != ele[3][20];
    ele[3][17] != ele[3][21];
    ele[3][17] != ele[3][22];
    ele[3][17] != ele[3][23];
    ele[3][17] != ele[3][24];
    ele[3][17] != ele[3][25];
    ele[3][17] != ele[3][26];
    ele[3][17] != ele[3][27];
    ele[3][17] != ele[3][28];
    ele[3][17] != ele[3][29];
    ele[3][17] != ele[3][30];
    ele[3][17] != ele[3][31];
    ele[3][17] != ele[3][32];
    ele[3][17] != ele[3][33];
    ele[3][17] != ele[3][34];
    ele[3][17] != ele[3][35];
    ele[3][17] != ele[30][17];
    ele[3][17] != ele[31][17];
    ele[3][17] != ele[32][17];
    ele[3][17] != ele[33][17];
    ele[3][17] != ele[34][17];
    ele[3][17] != ele[35][17];
    ele[3][17] != ele[4][12];
    ele[3][17] != ele[4][13];
    ele[3][17] != ele[4][14];
    ele[3][17] != ele[4][15];
    ele[3][17] != ele[4][16];
    ele[3][17] != ele[4][17];
    ele[3][17] != ele[5][12];
    ele[3][17] != ele[5][13];
    ele[3][17] != ele[5][14];
    ele[3][17] != ele[5][15];
    ele[3][17] != ele[5][16];
    ele[3][17] != ele[5][17];
    ele[3][17] != ele[6][17];
    ele[3][17] != ele[7][17];
    ele[3][17] != ele[8][17];
    ele[3][17] != ele[9][17];
    ele[3][18] != ele[10][18];
    ele[3][18] != ele[11][18];
    ele[3][18] != ele[12][18];
    ele[3][18] != ele[13][18];
    ele[3][18] != ele[14][18];
    ele[3][18] != ele[15][18];
    ele[3][18] != ele[16][18];
    ele[3][18] != ele[17][18];
    ele[3][18] != ele[18][18];
    ele[3][18] != ele[19][18];
    ele[3][18] != ele[20][18];
    ele[3][18] != ele[21][18];
    ele[3][18] != ele[22][18];
    ele[3][18] != ele[23][18];
    ele[3][18] != ele[24][18];
    ele[3][18] != ele[25][18];
    ele[3][18] != ele[26][18];
    ele[3][18] != ele[27][18];
    ele[3][18] != ele[28][18];
    ele[3][18] != ele[29][18];
    ele[3][18] != ele[3][19];
    ele[3][18] != ele[3][20];
    ele[3][18] != ele[3][21];
    ele[3][18] != ele[3][22];
    ele[3][18] != ele[3][23];
    ele[3][18] != ele[3][24];
    ele[3][18] != ele[3][25];
    ele[3][18] != ele[3][26];
    ele[3][18] != ele[3][27];
    ele[3][18] != ele[3][28];
    ele[3][18] != ele[3][29];
    ele[3][18] != ele[3][30];
    ele[3][18] != ele[3][31];
    ele[3][18] != ele[3][32];
    ele[3][18] != ele[3][33];
    ele[3][18] != ele[3][34];
    ele[3][18] != ele[3][35];
    ele[3][18] != ele[30][18];
    ele[3][18] != ele[31][18];
    ele[3][18] != ele[32][18];
    ele[3][18] != ele[33][18];
    ele[3][18] != ele[34][18];
    ele[3][18] != ele[35][18];
    ele[3][18] != ele[4][18];
    ele[3][18] != ele[4][19];
    ele[3][18] != ele[4][20];
    ele[3][18] != ele[4][21];
    ele[3][18] != ele[4][22];
    ele[3][18] != ele[4][23];
    ele[3][18] != ele[5][18];
    ele[3][18] != ele[5][19];
    ele[3][18] != ele[5][20];
    ele[3][18] != ele[5][21];
    ele[3][18] != ele[5][22];
    ele[3][18] != ele[5][23];
    ele[3][18] != ele[6][18];
    ele[3][18] != ele[7][18];
    ele[3][18] != ele[8][18];
    ele[3][18] != ele[9][18];
    ele[3][19] != ele[10][19];
    ele[3][19] != ele[11][19];
    ele[3][19] != ele[12][19];
    ele[3][19] != ele[13][19];
    ele[3][19] != ele[14][19];
    ele[3][19] != ele[15][19];
    ele[3][19] != ele[16][19];
    ele[3][19] != ele[17][19];
    ele[3][19] != ele[18][19];
    ele[3][19] != ele[19][19];
    ele[3][19] != ele[20][19];
    ele[3][19] != ele[21][19];
    ele[3][19] != ele[22][19];
    ele[3][19] != ele[23][19];
    ele[3][19] != ele[24][19];
    ele[3][19] != ele[25][19];
    ele[3][19] != ele[26][19];
    ele[3][19] != ele[27][19];
    ele[3][19] != ele[28][19];
    ele[3][19] != ele[29][19];
    ele[3][19] != ele[3][20];
    ele[3][19] != ele[3][21];
    ele[3][19] != ele[3][22];
    ele[3][19] != ele[3][23];
    ele[3][19] != ele[3][24];
    ele[3][19] != ele[3][25];
    ele[3][19] != ele[3][26];
    ele[3][19] != ele[3][27];
    ele[3][19] != ele[3][28];
    ele[3][19] != ele[3][29];
    ele[3][19] != ele[3][30];
    ele[3][19] != ele[3][31];
    ele[3][19] != ele[3][32];
    ele[3][19] != ele[3][33];
    ele[3][19] != ele[3][34];
    ele[3][19] != ele[3][35];
    ele[3][19] != ele[30][19];
    ele[3][19] != ele[31][19];
    ele[3][19] != ele[32][19];
    ele[3][19] != ele[33][19];
    ele[3][19] != ele[34][19];
    ele[3][19] != ele[35][19];
    ele[3][19] != ele[4][18];
    ele[3][19] != ele[4][19];
    ele[3][19] != ele[4][20];
    ele[3][19] != ele[4][21];
    ele[3][19] != ele[4][22];
    ele[3][19] != ele[4][23];
    ele[3][19] != ele[5][18];
    ele[3][19] != ele[5][19];
    ele[3][19] != ele[5][20];
    ele[3][19] != ele[5][21];
    ele[3][19] != ele[5][22];
    ele[3][19] != ele[5][23];
    ele[3][19] != ele[6][19];
    ele[3][19] != ele[7][19];
    ele[3][19] != ele[8][19];
    ele[3][19] != ele[9][19];
    ele[3][2] != ele[10][2];
    ele[3][2] != ele[11][2];
    ele[3][2] != ele[12][2];
    ele[3][2] != ele[13][2];
    ele[3][2] != ele[14][2];
    ele[3][2] != ele[15][2];
    ele[3][2] != ele[16][2];
    ele[3][2] != ele[17][2];
    ele[3][2] != ele[18][2];
    ele[3][2] != ele[19][2];
    ele[3][2] != ele[20][2];
    ele[3][2] != ele[21][2];
    ele[3][2] != ele[22][2];
    ele[3][2] != ele[23][2];
    ele[3][2] != ele[24][2];
    ele[3][2] != ele[25][2];
    ele[3][2] != ele[26][2];
    ele[3][2] != ele[27][2];
    ele[3][2] != ele[28][2];
    ele[3][2] != ele[29][2];
    ele[3][2] != ele[3][10];
    ele[3][2] != ele[3][11];
    ele[3][2] != ele[3][12];
    ele[3][2] != ele[3][13];
    ele[3][2] != ele[3][14];
    ele[3][2] != ele[3][15];
    ele[3][2] != ele[3][16];
    ele[3][2] != ele[3][17];
    ele[3][2] != ele[3][18];
    ele[3][2] != ele[3][19];
    ele[3][2] != ele[3][20];
    ele[3][2] != ele[3][21];
    ele[3][2] != ele[3][22];
    ele[3][2] != ele[3][23];
    ele[3][2] != ele[3][24];
    ele[3][2] != ele[3][25];
    ele[3][2] != ele[3][26];
    ele[3][2] != ele[3][27];
    ele[3][2] != ele[3][28];
    ele[3][2] != ele[3][29];
    ele[3][2] != ele[3][3];
    ele[3][2] != ele[3][30];
    ele[3][2] != ele[3][31];
    ele[3][2] != ele[3][32];
    ele[3][2] != ele[3][33];
    ele[3][2] != ele[3][34];
    ele[3][2] != ele[3][35];
    ele[3][2] != ele[3][4];
    ele[3][2] != ele[3][5];
    ele[3][2] != ele[3][6];
    ele[3][2] != ele[3][7];
    ele[3][2] != ele[3][8];
    ele[3][2] != ele[3][9];
    ele[3][2] != ele[30][2];
    ele[3][2] != ele[31][2];
    ele[3][2] != ele[32][2];
    ele[3][2] != ele[33][2];
    ele[3][2] != ele[34][2];
    ele[3][2] != ele[35][2];
    ele[3][2] != ele[4][0];
    ele[3][2] != ele[4][1];
    ele[3][2] != ele[4][2];
    ele[3][2] != ele[4][3];
    ele[3][2] != ele[4][4];
    ele[3][2] != ele[4][5];
    ele[3][2] != ele[5][0];
    ele[3][2] != ele[5][1];
    ele[3][2] != ele[5][2];
    ele[3][2] != ele[5][3];
    ele[3][2] != ele[5][4];
    ele[3][2] != ele[5][5];
    ele[3][2] != ele[6][2];
    ele[3][2] != ele[7][2];
    ele[3][2] != ele[8][2];
    ele[3][2] != ele[9][2];
    ele[3][20] != ele[10][20];
    ele[3][20] != ele[11][20];
    ele[3][20] != ele[12][20];
    ele[3][20] != ele[13][20];
    ele[3][20] != ele[14][20];
    ele[3][20] != ele[15][20];
    ele[3][20] != ele[16][20];
    ele[3][20] != ele[17][20];
    ele[3][20] != ele[18][20];
    ele[3][20] != ele[19][20];
    ele[3][20] != ele[20][20];
    ele[3][20] != ele[21][20];
    ele[3][20] != ele[22][20];
    ele[3][20] != ele[23][20];
    ele[3][20] != ele[24][20];
    ele[3][20] != ele[25][20];
    ele[3][20] != ele[26][20];
    ele[3][20] != ele[27][20];
    ele[3][20] != ele[28][20];
    ele[3][20] != ele[29][20];
    ele[3][20] != ele[3][21];
    ele[3][20] != ele[3][22];
    ele[3][20] != ele[3][23];
    ele[3][20] != ele[3][24];
    ele[3][20] != ele[3][25];
    ele[3][20] != ele[3][26];
    ele[3][20] != ele[3][27];
    ele[3][20] != ele[3][28];
    ele[3][20] != ele[3][29];
    ele[3][20] != ele[3][30];
    ele[3][20] != ele[3][31];
    ele[3][20] != ele[3][32];
    ele[3][20] != ele[3][33];
    ele[3][20] != ele[3][34];
    ele[3][20] != ele[3][35];
    ele[3][20] != ele[30][20];
    ele[3][20] != ele[31][20];
    ele[3][20] != ele[32][20];
    ele[3][20] != ele[33][20];
    ele[3][20] != ele[34][20];
    ele[3][20] != ele[35][20];
    ele[3][20] != ele[4][18];
    ele[3][20] != ele[4][19];
    ele[3][20] != ele[4][20];
    ele[3][20] != ele[4][21];
    ele[3][20] != ele[4][22];
    ele[3][20] != ele[4][23];
    ele[3][20] != ele[5][18];
    ele[3][20] != ele[5][19];
    ele[3][20] != ele[5][20];
    ele[3][20] != ele[5][21];
    ele[3][20] != ele[5][22];
    ele[3][20] != ele[5][23];
    ele[3][20] != ele[6][20];
    ele[3][20] != ele[7][20];
    ele[3][20] != ele[8][20];
    ele[3][20] != ele[9][20];
    ele[3][21] != ele[10][21];
    ele[3][21] != ele[11][21];
    ele[3][21] != ele[12][21];
    ele[3][21] != ele[13][21];
    ele[3][21] != ele[14][21];
    ele[3][21] != ele[15][21];
    ele[3][21] != ele[16][21];
    ele[3][21] != ele[17][21];
    ele[3][21] != ele[18][21];
    ele[3][21] != ele[19][21];
    ele[3][21] != ele[20][21];
    ele[3][21] != ele[21][21];
    ele[3][21] != ele[22][21];
    ele[3][21] != ele[23][21];
    ele[3][21] != ele[24][21];
    ele[3][21] != ele[25][21];
    ele[3][21] != ele[26][21];
    ele[3][21] != ele[27][21];
    ele[3][21] != ele[28][21];
    ele[3][21] != ele[29][21];
    ele[3][21] != ele[3][22];
    ele[3][21] != ele[3][23];
    ele[3][21] != ele[3][24];
    ele[3][21] != ele[3][25];
    ele[3][21] != ele[3][26];
    ele[3][21] != ele[3][27];
    ele[3][21] != ele[3][28];
    ele[3][21] != ele[3][29];
    ele[3][21] != ele[3][30];
    ele[3][21] != ele[3][31];
    ele[3][21] != ele[3][32];
    ele[3][21] != ele[3][33];
    ele[3][21] != ele[3][34];
    ele[3][21] != ele[3][35];
    ele[3][21] != ele[30][21];
    ele[3][21] != ele[31][21];
    ele[3][21] != ele[32][21];
    ele[3][21] != ele[33][21];
    ele[3][21] != ele[34][21];
    ele[3][21] != ele[35][21];
    ele[3][21] != ele[4][18];
    ele[3][21] != ele[4][19];
    ele[3][21] != ele[4][20];
    ele[3][21] != ele[4][21];
    ele[3][21] != ele[4][22];
    ele[3][21] != ele[4][23];
    ele[3][21] != ele[5][18];
    ele[3][21] != ele[5][19];
    ele[3][21] != ele[5][20];
    ele[3][21] != ele[5][21];
    ele[3][21] != ele[5][22];
    ele[3][21] != ele[5][23];
    ele[3][21] != ele[6][21];
    ele[3][21] != ele[7][21];
    ele[3][21] != ele[8][21];
    ele[3][21] != ele[9][21];
    ele[3][22] != ele[10][22];
    ele[3][22] != ele[11][22];
    ele[3][22] != ele[12][22];
    ele[3][22] != ele[13][22];
    ele[3][22] != ele[14][22];
    ele[3][22] != ele[15][22];
    ele[3][22] != ele[16][22];
    ele[3][22] != ele[17][22];
    ele[3][22] != ele[18][22];
    ele[3][22] != ele[19][22];
    ele[3][22] != ele[20][22];
    ele[3][22] != ele[21][22];
    ele[3][22] != ele[22][22];
    ele[3][22] != ele[23][22];
    ele[3][22] != ele[24][22];
    ele[3][22] != ele[25][22];
    ele[3][22] != ele[26][22];
    ele[3][22] != ele[27][22];
    ele[3][22] != ele[28][22];
    ele[3][22] != ele[29][22];
    ele[3][22] != ele[3][23];
    ele[3][22] != ele[3][24];
    ele[3][22] != ele[3][25];
    ele[3][22] != ele[3][26];
    ele[3][22] != ele[3][27];
    ele[3][22] != ele[3][28];
    ele[3][22] != ele[3][29];
    ele[3][22] != ele[3][30];
    ele[3][22] != ele[3][31];
    ele[3][22] != ele[3][32];
    ele[3][22] != ele[3][33];
    ele[3][22] != ele[3][34];
    ele[3][22] != ele[3][35];
    ele[3][22] != ele[30][22];
    ele[3][22] != ele[31][22];
    ele[3][22] != ele[32][22];
    ele[3][22] != ele[33][22];
    ele[3][22] != ele[34][22];
    ele[3][22] != ele[35][22];
    ele[3][22] != ele[4][18];
    ele[3][22] != ele[4][19];
    ele[3][22] != ele[4][20];
    ele[3][22] != ele[4][21];
    ele[3][22] != ele[4][22];
    ele[3][22] != ele[4][23];
    ele[3][22] != ele[5][18];
    ele[3][22] != ele[5][19];
    ele[3][22] != ele[5][20];
    ele[3][22] != ele[5][21];
    ele[3][22] != ele[5][22];
    ele[3][22] != ele[5][23];
    ele[3][22] != ele[6][22];
    ele[3][22] != ele[7][22];
    ele[3][22] != ele[8][22];
    ele[3][22] != ele[9][22];
    ele[3][23] != ele[10][23];
    ele[3][23] != ele[11][23];
    ele[3][23] != ele[12][23];
    ele[3][23] != ele[13][23];
    ele[3][23] != ele[14][23];
    ele[3][23] != ele[15][23];
    ele[3][23] != ele[16][23];
    ele[3][23] != ele[17][23];
    ele[3][23] != ele[18][23];
    ele[3][23] != ele[19][23];
    ele[3][23] != ele[20][23];
    ele[3][23] != ele[21][23];
    ele[3][23] != ele[22][23];
    ele[3][23] != ele[23][23];
    ele[3][23] != ele[24][23];
    ele[3][23] != ele[25][23];
    ele[3][23] != ele[26][23];
    ele[3][23] != ele[27][23];
    ele[3][23] != ele[28][23];
    ele[3][23] != ele[29][23];
    ele[3][23] != ele[3][24];
    ele[3][23] != ele[3][25];
    ele[3][23] != ele[3][26];
    ele[3][23] != ele[3][27];
    ele[3][23] != ele[3][28];
    ele[3][23] != ele[3][29];
    ele[3][23] != ele[3][30];
    ele[3][23] != ele[3][31];
    ele[3][23] != ele[3][32];
    ele[3][23] != ele[3][33];
    ele[3][23] != ele[3][34];
    ele[3][23] != ele[3][35];
    ele[3][23] != ele[30][23];
    ele[3][23] != ele[31][23];
    ele[3][23] != ele[32][23];
    ele[3][23] != ele[33][23];
    ele[3][23] != ele[34][23];
    ele[3][23] != ele[35][23];
    ele[3][23] != ele[4][18];
    ele[3][23] != ele[4][19];
    ele[3][23] != ele[4][20];
    ele[3][23] != ele[4][21];
    ele[3][23] != ele[4][22];
    ele[3][23] != ele[4][23];
    ele[3][23] != ele[5][18];
    ele[3][23] != ele[5][19];
    ele[3][23] != ele[5][20];
    ele[3][23] != ele[5][21];
    ele[3][23] != ele[5][22];
    ele[3][23] != ele[5][23];
    ele[3][23] != ele[6][23];
    ele[3][23] != ele[7][23];
    ele[3][23] != ele[8][23];
    ele[3][23] != ele[9][23];
    ele[3][24] != ele[10][24];
    ele[3][24] != ele[11][24];
    ele[3][24] != ele[12][24];
    ele[3][24] != ele[13][24];
    ele[3][24] != ele[14][24];
    ele[3][24] != ele[15][24];
    ele[3][24] != ele[16][24];
    ele[3][24] != ele[17][24];
    ele[3][24] != ele[18][24];
    ele[3][24] != ele[19][24];
    ele[3][24] != ele[20][24];
    ele[3][24] != ele[21][24];
    ele[3][24] != ele[22][24];
    ele[3][24] != ele[23][24];
    ele[3][24] != ele[24][24];
    ele[3][24] != ele[25][24];
    ele[3][24] != ele[26][24];
    ele[3][24] != ele[27][24];
    ele[3][24] != ele[28][24];
    ele[3][24] != ele[29][24];
    ele[3][24] != ele[3][25];
    ele[3][24] != ele[3][26];
    ele[3][24] != ele[3][27];
    ele[3][24] != ele[3][28];
    ele[3][24] != ele[3][29];
    ele[3][24] != ele[3][30];
    ele[3][24] != ele[3][31];
    ele[3][24] != ele[3][32];
    ele[3][24] != ele[3][33];
    ele[3][24] != ele[3][34];
    ele[3][24] != ele[3][35];
    ele[3][24] != ele[30][24];
    ele[3][24] != ele[31][24];
    ele[3][24] != ele[32][24];
    ele[3][24] != ele[33][24];
    ele[3][24] != ele[34][24];
    ele[3][24] != ele[35][24];
    ele[3][24] != ele[4][24];
    ele[3][24] != ele[4][25];
    ele[3][24] != ele[4][26];
    ele[3][24] != ele[4][27];
    ele[3][24] != ele[4][28];
    ele[3][24] != ele[4][29];
    ele[3][24] != ele[5][24];
    ele[3][24] != ele[5][25];
    ele[3][24] != ele[5][26];
    ele[3][24] != ele[5][27];
    ele[3][24] != ele[5][28];
    ele[3][24] != ele[5][29];
    ele[3][24] != ele[6][24];
    ele[3][24] != ele[7][24];
    ele[3][24] != ele[8][24];
    ele[3][24] != ele[9][24];
    ele[3][25] != ele[10][25];
    ele[3][25] != ele[11][25];
    ele[3][25] != ele[12][25];
    ele[3][25] != ele[13][25];
    ele[3][25] != ele[14][25];
    ele[3][25] != ele[15][25];
    ele[3][25] != ele[16][25];
    ele[3][25] != ele[17][25];
    ele[3][25] != ele[18][25];
    ele[3][25] != ele[19][25];
    ele[3][25] != ele[20][25];
    ele[3][25] != ele[21][25];
    ele[3][25] != ele[22][25];
    ele[3][25] != ele[23][25];
    ele[3][25] != ele[24][25];
    ele[3][25] != ele[25][25];
    ele[3][25] != ele[26][25];
    ele[3][25] != ele[27][25];
    ele[3][25] != ele[28][25];
    ele[3][25] != ele[29][25];
    ele[3][25] != ele[3][26];
    ele[3][25] != ele[3][27];
    ele[3][25] != ele[3][28];
    ele[3][25] != ele[3][29];
    ele[3][25] != ele[3][30];
    ele[3][25] != ele[3][31];
    ele[3][25] != ele[3][32];
    ele[3][25] != ele[3][33];
    ele[3][25] != ele[3][34];
    ele[3][25] != ele[3][35];
    ele[3][25] != ele[30][25];
    ele[3][25] != ele[31][25];
    ele[3][25] != ele[32][25];
    ele[3][25] != ele[33][25];
    ele[3][25] != ele[34][25];
    ele[3][25] != ele[35][25];
    ele[3][25] != ele[4][24];
    ele[3][25] != ele[4][25];
    ele[3][25] != ele[4][26];
    ele[3][25] != ele[4][27];
    ele[3][25] != ele[4][28];
    ele[3][25] != ele[4][29];
    ele[3][25] != ele[5][24];
    ele[3][25] != ele[5][25];
    ele[3][25] != ele[5][26];
    ele[3][25] != ele[5][27];
    ele[3][25] != ele[5][28];
    ele[3][25] != ele[5][29];
    ele[3][25] != ele[6][25];
    ele[3][25] != ele[7][25];
    ele[3][25] != ele[8][25];
    ele[3][25] != ele[9][25];
    ele[3][26] != ele[10][26];
    ele[3][26] != ele[11][26];
    ele[3][26] != ele[12][26];
    ele[3][26] != ele[13][26];
    ele[3][26] != ele[14][26];
    ele[3][26] != ele[15][26];
    ele[3][26] != ele[16][26];
    ele[3][26] != ele[17][26];
    ele[3][26] != ele[18][26];
    ele[3][26] != ele[19][26];
    ele[3][26] != ele[20][26];
    ele[3][26] != ele[21][26];
    ele[3][26] != ele[22][26];
    ele[3][26] != ele[23][26];
    ele[3][26] != ele[24][26];
    ele[3][26] != ele[25][26];
    ele[3][26] != ele[26][26];
    ele[3][26] != ele[27][26];
    ele[3][26] != ele[28][26];
    ele[3][26] != ele[29][26];
    ele[3][26] != ele[3][27];
    ele[3][26] != ele[3][28];
    ele[3][26] != ele[3][29];
    ele[3][26] != ele[3][30];
    ele[3][26] != ele[3][31];
    ele[3][26] != ele[3][32];
    ele[3][26] != ele[3][33];
    ele[3][26] != ele[3][34];
    ele[3][26] != ele[3][35];
    ele[3][26] != ele[30][26];
    ele[3][26] != ele[31][26];
    ele[3][26] != ele[32][26];
    ele[3][26] != ele[33][26];
    ele[3][26] != ele[34][26];
    ele[3][26] != ele[35][26];
    ele[3][26] != ele[4][24];
    ele[3][26] != ele[4][25];
    ele[3][26] != ele[4][26];
    ele[3][26] != ele[4][27];
    ele[3][26] != ele[4][28];
    ele[3][26] != ele[4][29];
    ele[3][26] != ele[5][24];
    ele[3][26] != ele[5][25];
    ele[3][26] != ele[5][26];
    ele[3][26] != ele[5][27];
    ele[3][26] != ele[5][28];
    ele[3][26] != ele[5][29];
    ele[3][26] != ele[6][26];
    ele[3][26] != ele[7][26];
    ele[3][26] != ele[8][26];
    ele[3][26] != ele[9][26];
    ele[3][27] != ele[10][27];
    ele[3][27] != ele[11][27];
    ele[3][27] != ele[12][27];
    ele[3][27] != ele[13][27];
    ele[3][27] != ele[14][27];
    ele[3][27] != ele[15][27];
    ele[3][27] != ele[16][27];
    ele[3][27] != ele[17][27];
    ele[3][27] != ele[18][27];
    ele[3][27] != ele[19][27];
    ele[3][27] != ele[20][27];
    ele[3][27] != ele[21][27];
    ele[3][27] != ele[22][27];
    ele[3][27] != ele[23][27];
    ele[3][27] != ele[24][27];
    ele[3][27] != ele[25][27];
    ele[3][27] != ele[26][27];
    ele[3][27] != ele[27][27];
    ele[3][27] != ele[28][27];
    ele[3][27] != ele[29][27];
    ele[3][27] != ele[3][28];
    ele[3][27] != ele[3][29];
    ele[3][27] != ele[3][30];
    ele[3][27] != ele[3][31];
    ele[3][27] != ele[3][32];
    ele[3][27] != ele[3][33];
    ele[3][27] != ele[3][34];
    ele[3][27] != ele[3][35];
    ele[3][27] != ele[30][27];
    ele[3][27] != ele[31][27];
    ele[3][27] != ele[32][27];
    ele[3][27] != ele[33][27];
    ele[3][27] != ele[34][27];
    ele[3][27] != ele[35][27];
    ele[3][27] != ele[4][24];
    ele[3][27] != ele[4][25];
    ele[3][27] != ele[4][26];
    ele[3][27] != ele[4][27];
    ele[3][27] != ele[4][28];
    ele[3][27] != ele[4][29];
    ele[3][27] != ele[5][24];
    ele[3][27] != ele[5][25];
    ele[3][27] != ele[5][26];
    ele[3][27] != ele[5][27];
    ele[3][27] != ele[5][28];
    ele[3][27] != ele[5][29];
    ele[3][27] != ele[6][27];
    ele[3][27] != ele[7][27];
    ele[3][27] != ele[8][27];
    ele[3][27] != ele[9][27];
    ele[3][28] != ele[10][28];
    ele[3][28] != ele[11][28];
    ele[3][28] != ele[12][28];
    ele[3][28] != ele[13][28];
    ele[3][28] != ele[14][28];
    ele[3][28] != ele[15][28];
    ele[3][28] != ele[16][28];
    ele[3][28] != ele[17][28];
    ele[3][28] != ele[18][28];
    ele[3][28] != ele[19][28];
    ele[3][28] != ele[20][28];
    ele[3][28] != ele[21][28];
    ele[3][28] != ele[22][28];
    ele[3][28] != ele[23][28];
    ele[3][28] != ele[24][28];
    ele[3][28] != ele[25][28];
    ele[3][28] != ele[26][28];
    ele[3][28] != ele[27][28];
    ele[3][28] != ele[28][28];
    ele[3][28] != ele[29][28];
    ele[3][28] != ele[3][29];
    ele[3][28] != ele[3][30];
    ele[3][28] != ele[3][31];
    ele[3][28] != ele[3][32];
    ele[3][28] != ele[3][33];
    ele[3][28] != ele[3][34];
    ele[3][28] != ele[3][35];
    ele[3][28] != ele[30][28];
    ele[3][28] != ele[31][28];
    ele[3][28] != ele[32][28];
    ele[3][28] != ele[33][28];
    ele[3][28] != ele[34][28];
    ele[3][28] != ele[35][28];
    ele[3][28] != ele[4][24];
    ele[3][28] != ele[4][25];
    ele[3][28] != ele[4][26];
    ele[3][28] != ele[4][27];
    ele[3][28] != ele[4][28];
    ele[3][28] != ele[4][29];
    ele[3][28] != ele[5][24];
    ele[3][28] != ele[5][25];
    ele[3][28] != ele[5][26];
    ele[3][28] != ele[5][27];
    ele[3][28] != ele[5][28];
    ele[3][28] != ele[5][29];
    ele[3][28] != ele[6][28];
    ele[3][28] != ele[7][28];
    ele[3][28] != ele[8][28];
    ele[3][28] != ele[9][28];
    ele[3][29] != ele[10][29];
    ele[3][29] != ele[11][29];
    ele[3][29] != ele[12][29];
    ele[3][29] != ele[13][29];
    ele[3][29] != ele[14][29];
    ele[3][29] != ele[15][29];
    ele[3][29] != ele[16][29];
    ele[3][29] != ele[17][29];
    ele[3][29] != ele[18][29];
    ele[3][29] != ele[19][29];
    ele[3][29] != ele[20][29];
    ele[3][29] != ele[21][29];
    ele[3][29] != ele[22][29];
    ele[3][29] != ele[23][29];
    ele[3][29] != ele[24][29];
    ele[3][29] != ele[25][29];
    ele[3][29] != ele[26][29];
    ele[3][29] != ele[27][29];
    ele[3][29] != ele[28][29];
    ele[3][29] != ele[29][29];
    ele[3][29] != ele[3][30];
    ele[3][29] != ele[3][31];
    ele[3][29] != ele[3][32];
    ele[3][29] != ele[3][33];
    ele[3][29] != ele[3][34];
    ele[3][29] != ele[3][35];
    ele[3][29] != ele[30][29];
    ele[3][29] != ele[31][29];
    ele[3][29] != ele[32][29];
    ele[3][29] != ele[33][29];
    ele[3][29] != ele[34][29];
    ele[3][29] != ele[35][29];
    ele[3][29] != ele[4][24];
    ele[3][29] != ele[4][25];
    ele[3][29] != ele[4][26];
    ele[3][29] != ele[4][27];
    ele[3][29] != ele[4][28];
    ele[3][29] != ele[4][29];
    ele[3][29] != ele[5][24];
    ele[3][29] != ele[5][25];
    ele[3][29] != ele[5][26];
    ele[3][29] != ele[5][27];
    ele[3][29] != ele[5][28];
    ele[3][29] != ele[5][29];
    ele[3][29] != ele[6][29];
    ele[3][29] != ele[7][29];
    ele[3][29] != ele[8][29];
    ele[3][29] != ele[9][29];
    ele[3][3] != ele[10][3];
    ele[3][3] != ele[11][3];
    ele[3][3] != ele[12][3];
    ele[3][3] != ele[13][3];
    ele[3][3] != ele[14][3];
    ele[3][3] != ele[15][3];
    ele[3][3] != ele[16][3];
    ele[3][3] != ele[17][3];
    ele[3][3] != ele[18][3];
    ele[3][3] != ele[19][3];
    ele[3][3] != ele[20][3];
    ele[3][3] != ele[21][3];
    ele[3][3] != ele[22][3];
    ele[3][3] != ele[23][3];
    ele[3][3] != ele[24][3];
    ele[3][3] != ele[25][3];
    ele[3][3] != ele[26][3];
    ele[3][3] != ele[27][3];
    ele[3][3] != ele[28][3];
    ele[3][3] != ele[29][3];
    ele[3][3] != ele[3][10];
    ele[3][3] != ele[3][11];
    ele[3][3] != ele[3][12];
    ele[3][3] != ele[3][13];
    ele[3][3] != ele[3][14];
    ele[3][3] != ele[3][15];
    ele[3][3] != ele[3][16];
    ele[3][3] != ele[3][17];
    ele[3][3] != ele[3][18];
    ele[3][3] != ele[3][19];
    ele[3][3] != ele[3][20];
    ele[3][3] != ele[3][21];
    ele[3][3] != ele[3][22];
    ele[3][3] != ele[3][23];
    ele[3][3] != ele[3][24];
    ele[3][3] != ele[3][25];
    ele[3][3] != ele[3][26];
    ele[3][3] != ele[3][27];
    ele[3][3] != ele[3][28];
    ele[3][3] != ele[3][29];
    ele[3][3] != ele[3][30];
    ele[3][3] != ele[3][31];
    ele[3][3] != ele[3][32];
    ele[3][3] != ele[3][33];
    ele[3][3] != ele[3][34];
    ele[3][3] != ele[3][35];
    ele[3][3] != ele[3][4];
    ele[3][3] != ele[3][5];
    ele[3][3] != ele[3][6];
    ele[3][3] != ele[3][7];
    ele[3][3] != ele[3][8];
    ele[3][3] != ele[3][9];
    ele[3][3] != ele[30][3];
    ele[3][3] != ele[31][3];
    ele[3][3] != ele[32][3];
    ele[3][3] != ele[33][3];
    ele[3][3] != ele[34][3];
    ele[3][3] != ele[35][3];
    ele[3][3] != ele[4][0];
    ele[3][3] != ele[4][1];
    ele[3][3] != ele[4][2];
    ele[3][3] != ele[4][3];
    ele[3][3] != ele[4][4];
    ele[3][3] != ele[4][5];
    ele[3][3] != ele[5][0];
    ele[3][3] != ele[5][1];
    ele[3][3] != ele[5][2];
    ele[3][3] != ele[5][3];
    ele[3][3] != ele[5][4];
    ele[3][3] != ele[5][5];
    ele[3][3] != ele[6][3];
    ele[3][3] != ele[7][3];
    ele[3][3] != ele[8][3];
    ele[3][3] != ele[9][3];
    ele[3][30] != ele[10][30];
    ele[3][30] != ele[11][30];
    ele[3][30] != ele[12][30];
    ele[3][30] != ele[13][30];
    ele[3][30] != ele[14][30];
    ele[3][30] != ele[15][30];
    ele[3][30] != ele[16][30];
    ele[3][30] != ele[17][30];
    ele[3][30] != ele[18][30];
    ele[3][30] != ele[19][30];
    ele[3][30] != ele[20][30];
    ele[3][30] != ele[21][30];
    ele[3][30] != ele[22][30];
    ele[3][30] != ele[23][30];
    ele[3][30] != ele[24][30];
    ele[3][30] != ele[25][30];
    ele[3][30] != ele[26][30];
    ele[3][30] != ele[27][30];
    ele[3][30] != ele[28][30];
    ele[3][30] != ele[29][30];
    ele[3][30] != ele[3][31];
    ele[3][30] != ele[3][32];
    ele[3][30] != ele[3][33];
    ele[3][30] != ele[3][34];
    ele[3][30] != ele[3][35];
    ele[3][30] != ele[30][30];
    ele[3][30] != ele[31][30];
    ele[3][30] != ele[32][30];
    ele[3][30] != ele[33][30];
    ele[3][30] != ele[34][30];
    ele[3][30] != ele[35][30];
    ele[3][30] != ele[4][30];
    ele[3][30] != ele[4][31];
    ele[3][30] != ele[4][32];
    ele[3][30] != ele[4][33];
    ele[3][30] != ele[4][34];
    ele[3][30] != ele[4][35];
    ele[3][30] != ele[5][30];
    ele[3][30] != ele[5][31];
    ele[3][30] != ele[5][32];
    ele[3][30] != ele[5][33];
    ele[3][30] != ele[5][34];
    ele[3][30] != ele[5][35];
    ele[3][30] != ele[6][30];
    ele[3][30] != ele[7][30];
    ele[3][30] != ele[8][30];
    ele[3][30] != ele[9][30];
    ele[3][31] != ele[10][31];
    ele[3][31] != ele[11][31];
    ele[3][31] != ele[12][31];
    ele[3][31] != ele[13][31];
    ele[3][31] != ele[14][31];
    ele[3][31] != ele[15][31];
    ele[3][31] != ele[16][31];
    ele[3][31] != ele[17][31];
    ele[3][31] != ele[18][31];
    ele[3][31] != ele[19][31];
    ele[3][31] != ele[20][31];
    ele[3][31] != ele[21][31];
    ele[3][31] != ele[22][31];
    ele[3][31] != ele[23][31];
    ele[3][31] != ele[24][31];
    ele[3][31] != ele[25][31];
    ele[3][31] != ele[26][31];
    ele[3][31] != ele[27][31];
    ele[3][31] != ele[28][31];
    ele[3][31] != ele[29][31];
    ele[3][31] != ele[3][32];
    ele[3][31] != ele[3][33];
    ele[3][31] != ele[3][34];
    ele[3][31] != ele[3][35];
    ele[3][31] != ele[30][31];
    ele[3][31] != ele[31][31];
    ele[3][31] != ele[32][31];
    ele[3][31] != ele[33][31];
    ele[3][31] != ele[34][31];
    ele[3][31] != ele[35][31];
    ele[3][31] != ele[4][30];
    ele[3][31] != ele[4][31];
    ele[3][31] != ele[4][32];
    ele[3][31] != ele[4][33];
    ele[3][31] != ele[4][34];
    ele[3][31] != ele[4][35];
    ele[3][31] != ele[5][30];
    ele[3][31] != ele[5][31];
    ele[3][31] != ele[5][32];
    ele[3][31] != ele[5][33];
    ele[3][31] != ele[5][34];
    ele[3][31] != ele[5][35];
    ele[3][31] != ele[6][31];
    ele[3][31] != ele[7][31];
    ele[3][31] != ele[8][31];
    ele[3][31] != ele[9][31];
    ele[3][32] != ele[10][32];
    ele[3][32] != ele[11][32];
    ele[3][32] != ele[12][32];
    ele[3][32] != ele[13][32];
    ele[3][32] != ele[14][32];
    ele[3][32] != ele[15][32];
    ele[3][32] != ele[16][32];
    ele[3][32] != ele[17][32];
    ele[3][32] != ele[18][32];
    ele[3][32] != ele[19][32];
    ele[3][32] != ele[20][32];
    ele[3][32] != ele[21][32];
    ele[3][32] != ele[22][32];
    ele[3][32] != ele[23][32];
    ele[3][32] != ele[24][32];
    ele[3][32] != ele[25][32];
    ele[3][32] != ele[26][32];
    ele[3][32] != ele[27][32];
    ele[3][32] != ele[28][32];
    ele[3][32] != ele[29][32];
    ele[3][32] != ele[3][33];
    ele[3][32] != ele[3][34];
    ele[3][32] != ele[3][35];
    ele[3][32] != ele[30][32];
    ele[3][32] != ele[31][32];
    ele[3][32] != ele[32][32];
    ele[3][32] != ele[33][32];
    ele[3][32] != ele[34][32];
    ele[3][32] != ele[35][32];
    ele[3][32] != ele[4][30];
    ele[3][32] != ele[4][31];
    ele[3][32] != ele[4][32];
    ele[3][32] != ele[4][33];
    ele[3][32] != ele[4][34];
    ele[3][32] != ele[4][35];
    ele[3][32] != ele[5][30];
    ele[3][32] != ele[5][31];
    ele[3][32] != ele[5][32];
    ele[3][32] != ele[5][33];
    ele[3][32] != ele[5][34];
    ele[3][32] != ele[5][35];
    ele[3][32] != ele[6][32];
    ele[3][32] != ele[7][32];
    ele[3][32] != ele[8][32];
    ele[3][32] != ele[9][32];
    ele[3][33] != ele[10][33];
    ele[3][33] != ele[11][33];
    ele[3][33] != ele[12][33];
    ele[3][33] != ele[13][33];
    ele[3][33] != ele[14][33];
    ele[3][33] != ele[15][33];
    ele[3][33] != ele[16][33];
    ele[3][33] != ele[17][33];
    ele[3][33] != ele[18][33];
    ele[3][33] != ele[19][33];
    ele[3][33] != ele[20][33];
    ele[3][33] != ele[21][33];
    ele[3][33] != ele[22][33];
    ele[3][33] != ele[23][33];
    ele[3][33] != ele[24][33];
    ele[3][33] != ele[25][33];
    ele[3][33] != ele[26][33];
    ele[3][33] != ele[27][33];
    ele[3][33] != ele[28][33];
    ele[3][33] != ele[29][33];
    ele[3][33] != ele[3][34];
    ele[3][33] != ele[3][35];
    ele[3][33] != ele[30][33];
    ele[3][33] != ele[31][33];
    ele[3][33] != ele[32][33];
    ele[3][33] != ele[33][33];
    ele[3][33] != ele[34][33];
    ele[3][33] != ele[35][33];
    ele[3][33] != ele[4][30];
    ele[3][33] != ele[4][31];
    ele[3][33] != ele[4][32];
    ele[3][33] != ele[4][33];
    ele[3][33] != ele[4][34];
    ele[3][33] != ele[4][35];
    ele[3][33] != ele[5][30];
    ele[3][33] != ele[5][31];
    ele[3][33] != ele[5][32];
    ele[3][33] != ele[5][33];
    ele[3][33] != ele[5][34];
    ele[3][33] != ele[5][35];
    ele[3][33] != ele[6][33];
    ele[3][33] != ele[7][33];
    ele[3][33] != ele[8][33];
    ele[3][33] != ele[9][33];
    ele[3][34] != ele[10][34];
    ele[3][34] != ele[11][34];
    ele[3][34] != ele[12][34];
    ele[3][34] != ele[13][34];
    ele[3][34] != ele[14][34];
    ele[3][34] != ele[15][34];
    ele[3][34] != ele[16][34];
    ele[3][34] != ele[17][34];
    ele[3][34] != ele[18][34];
    ele[3][34] != ele[19][34];
    ele[3][34] != ele[20][34];
    ele[3][34] != ele[21][34];
    ele[3][34] != ele[22][34];
    ele[3][34] != ele[23][34];
    ele[3][34] != ele[24][34];
    ele[3][34] != ele[25][34];
    ele[3][34] != ele[26][34];
    ele[3][34] != ele[27][34];
    ele[3][34] != ele[28][34];
    ele[3][34] != ele[29][34];
    ele[3][34] != ele[3][35];
    ele[3][34] != ele[30][34];
    ele[3][34] != ele[31][34];
    ele[3][34] != ele[32][34];
    ele[3][34] != ele[33][34];
    ele[3][34] != ele[34][34];
    ele[3][34] != ele[35][34];
    ele[3][34] != ele[4][30];
    ele[3][34] != ele[4][31];
    ele[3][34] != ele[4][32];
    ele[3][34] != ele[4][33];
    ele[3][34] != ele[4][34];
    ele[3][34] != ele[4][35];
    ele[3][34] != ele[5][30];
    ele[3][34] != ele[5][31];
    ele[3][34] != ele[5][32];
    ele[3][34] != ele[5][33];
    ele[3][34] != ele[5][34];
    ele[3][34] != ele[5][35];
    ele[3][34] != ele[6][34];
    ele[3][34] != ele[7][34];
    ele[3][34] != ele[8][34];
    ele[3][34] != ele[9][34];
    ele[3][35] != ele[10][35];
    ele[3][35] != ele[11][35];
    ele[3][35] != ele[12][35];
    ele[3][35] != ele[13][35];
    ele[3][35] != ele[14][35];
    ele[3][35] != ele[15][35];
    ele[3][35] != ele[16][35];
    ele[3][35] != ele[17][35];
    ele[3][35] != ele[18][35];
    ele[3][35] != ele[19][35];
    ele[3][35] != ele[20][35];
    ele[3][35] != ele[21][35];
    ele[3][35] != ele[22][35];
    ele[3][35] != ele[23][35];
    ele[3][35] != ele[24][35];
    ele[3][35] != ele[25][35];
    ele[3][35] != ele[26][35];
    ele[3][35] != ele[27][35];
    ele[3][35] != ele[28][35];
    ele[3][35] != ele[29][35];
    ele[3][35] != ele[30][35];
    ele[3][35] != ele[31][35];
    ele[3][35] != ele[32][35];
    ele[3][35] != ele[33][35];
    ele[3][35] != ele[34][35];
    ele[3][35] != ele[35][35];
    ele[3][35] != ele[4][30];
    ele[3][35] != ele[4][31];
    ele[3][35] != ele[4][32];
    ele[3][35] != ele[4][33];
    ele[3][35] != ele[4][34];
    ele[3][35] != ele[4][35];
    ele[3][35] != ele[5][30];
    ele[3][35] != ele[5][31];
    ele[3][35] != ele[5][32];
    ele[3][35] != ele[5][33];
    ele[3][35] != ele[5][34];
    ele[3][35] != ele[5][35];
    ele[3][35] != ele[6][35];
    ele[3][35] != ele[7][35];
    ele[3][35] != ele[8][35];
    ele[3][35] != ele[9][35];
    ele[3][4] != ele[10][4];
    ele[3][4] != ele[11][4];
    ele[3][4] != ele[12][4];
    ele[3][4] != ele[13][4];
    ele[3][4] != ele[14][4];
    ele[3][4] != ele[15][4];
    ele[3][4] != ele[16][4];
    ele[3][4] != ele[17][4];
    ele[3][4] != ele[18][4];
    ele[3][4] != ele[19][4];
    ele[3][4] != ele[20][4];
    ele[3][4] != ele[21][4];
    ele[3][4] != ele[22][4];
    ele[3][4] != ele[23][4];
    ele[3][4] != ele[24][4];
    ele[3][4] != ele[25][4];
    ele[3][4] != ele[26][4];
    ele[3][4] != ele[27][4];
    ele[3][4] != ele[28][4];
    ele[3][4] != ele[29][4];
    ele[3][4] != ele[3][10];
    ele[3][4] != ele[3][11];
    ele[3][4] != ele[3][12];
    ele[3][4] != ele[3][13];
    ele[3][4] != ele[3][14];
    ele[3][4] != ele[3][15];
    ele[3][4] != ele[3][16];
    ele[3][4] != ele[3][17];
    ele[3][4] != ele[3][18];
    ele[3][4] != ele[3][19];
    ele[3][4] != ele[3][20];
    ele[3][4] != ele[3][21];
    ele[3][4] != ele[3][22];
    ele[3][4] != ele[3][23];
    ele[3][4] != ele[3][24];
    ele[3][4] != ele[3][25];
    ele[3][4] != ele[3][26];
    ele[3][4] != ele[3][27];
    ele[3][4] != ele[3][28];
    ele[3][4] != ele[3][29];
    ele[3][4] != ele[3][30];
    ele[3][4] != ele[3][31];
    ele[3][4] != ele[3][32];
    ele[3][4] != ele[3][33];
    ele[3][4] != ele[3][34];
    ele[3][4] != ele[3][35];
    ele[3][4] != ele[3][5];
    ele[3][4] != ele[3][6];
    ele[3][4] != ele[3][7];
    ele[3][4] != ele[3][8];
    ele[3][4] != ele[3][9];
    ele[3][4] != ele[30][4];
    ele[3][4] != ele[31][4];
    ele[3][4] != ele[32][4];
    ele[3][4] != ele[33][4];
    ele[3][4] != ele[34][4];
    ele[3][4] != ele[35][4];
    ele[3][4] != ele[4][0];
    ele[3][4] != ele[4][1];
    ele[3][4] != ele[4][2];
    ele[3][4] != ele[4][3];
    ele[3][4] != ele[4][4];
    ele[3][4] != ele[4][5];
    ele[3][4] != ele[5][0];
    ele[3][4] != ele[5][1];
    ele[3][4] != ele[5][2];
    ele[3][4] != ele[5][3];
    ele[3][4] != ele[5][4];
    ele[3][4] != ele[5][5];
    ele[3][4] != ele[6][4];
    ele[3][4] != ele[7][4];
    ele[3][4] != ele[8][4];
    ele[3][4] != ele[9][4];
    ele[3][5] != ele[10][5];
    ele[3][5] != ele[11][5];
    ele[3][5] != ele[12][5];
    ele[3][5] != ele[13][5];
    ele[3][5] != ele[14][5];
    ele[3][5] != ele[15][5];
    ele[3][5] != ele[16][5];
    ele[3][5] != ele[17][5];
    ele[3][5] != ele[18][5];
    ele[3][5] != ele[19][5];
    ele[3][5] != ele[20][5];
    ele[3][5] != ele[21][5];
    ele[3][5] != ele[22][5];
    ele[3][5] != ele[23][5];
    ele[3][5] != ele[24][5];
    ele[3][5] != ele[25][5];
    ele[3][5] != ele[26][5];
    ele[3][5] != ele[27][5];
    ele[3][5] != ele[28][5];
    ele[3][5] != ele[29][5];
    ele[3][5] != ele[3][10];
    ele[3][5] != ele[3][11];
    ele[3][5] != ele[3][12];
    ele[3][5] != ele[3][13];
    ele[3][5] != ele[3][14];
    ele[3][5] != ele[3][15];
    ele[3][5] != ele[3][16];
    ele[3][5] != ele[3][17];
    ele[3][5] != ele[3][18];
    ele[3][5] != ele[3][19];
    ele[3][5] != ele[3][20];
    ele[3][5] != ele[3][21];
    ele[3][5] != ele[3][22];
    ele[3][5] != ele[3][23];
    ele[3][5] != ele[3][24];
    ele[3][5] != ele[3][25];
    ele[3][5] != ele[3][26];
    ele[3][5] != ele[3][27];
    ele[3][5] != ele[3][28];
    ele[3][5] != ele[3][29];
    ele[3][5] != ele[3][30];
    ele[3][5] != ele[3][31];
    ele[3][5] != ele[3][32];
    ele[3][5] != ele[3][33];
    ele[3][5] != ele[3][34];
    ele[3][5] != ele[3][35];
    ele[3][5] != ele[3][6];
    ele[3][5] != ele[3][7];
    ele[3][5] != ele[3][8];
    ele[3][5] != ele[3][9];
    ele[3][5] != ele[30][5];
    ele[3][5] != ele[31][5];
    ele[3][5] != ele[32][5];
    ele[3][5] != ele[33][5];
    ele[3][5] != ele[34][5];
    ele[3][5] != ele[35][5];
    ele[3][5] != ele[4][0];
    ele[3][5] != ele[4][1];
    ele[3][5] != ele[4][2];
    ele[3][5] != ele[4][3];
    ele[3][5] != ele[4][4];
    ele[3][5] != ele[4][5];
    ele[3][5] != ele[5][0];
    ele[3][5] != ele[5][1];
    ele[3][5] != ele[5][2];
    ele[3][5] != ele[5][3];
    ele[3][5] != ele[5][4];
    ele[3][5] != ele[5][5];
    ele[3][5] != ele[6][5];
    ele[3][5] != ele[7][5];
    ele[3][5] != ele[8][5];
    ele[3][5] != ele[9][5];
    ele[3][6] != ele[10][6];
    ele[3][6] != ele[11][6];
    ele[3][6] != ele[12][6];
    ele[3][6] != ele[13][6];
    ele[3][6] != ele[14][6];
    ele[3][6] != ele[15][6];
    ele[3][6] != ele[16][6];
    ele[3][6] != ele[17][6];
    ele[3][6] != ele[18][6];
    ele[3][6] != ele[19][6];
    ele[3][6] != ele[20][6];
    ele[3][6] != ele[21][6];
    ele[3][6] != ele[22][6];
    ele[3][6] != ele[23][6];
    ele[3][6] != ele[24][6];
    ele[3][6] != ele[25][6];
    ele[3][6] != ele[26][6];
    ele[3][6] != ele[27][6];
    ele[3][6] != ele[28][6];
    ele[3][6] != ele[29][6];
    ele[3][6] != ele[3][10];
    ele[3][6] != ele[3][11];
    ele[3][6] != ele[3][12];
    ele[3][6] != ele[3][13];
    ele[3][6] != ele[3][14];
    ele[3][6] != ele[3][15];
    ele[3][6] != ele[3][16];
    ele[3][6] != ele[3][17];
    ele[3][6] != ele[3][18];
    ele[3][6] != ele[3][19];
    ele[3][6] != ele[3][20];
    ele[3][6] != ele[3][21];
    ele[3][6] != ele[3][22];
    ele[3][6] != ele[3][23];
    ele[3][6] != ele[3][24];
    ele[3][6] != ele[3][25];
    ele[3][6] != ele[3][26];
    ele[3][6] != ele[3][27];
    ele[3][6] != ele[3][28];
    ele[3][6] != ele[3][29];
    ele[3][6] != ele[3][30];
    ele[3][6] != ele[3][31];
    ele[3][6] != ele[3][32];
    ele[3][6] != ele[3][33];
    ele[3][6] != ele[3][34];
    ele[3][6] != ele[3][35];
    ele[3][6] != ele[3][7];
    ele[3][6] != ele[3][8];
    ele[3][6] != ele[3][9];
    ele[3][6] != ele[30][6];
    ele[3][6] != ele[31][6];
    ele[3][6] != ele[32][6];
    ele[3][6] != ele[33][6];
    ele[3][6] != ele[34][6];
    ele[3][6] != ele[35][6];
    ele[3][6] != ele[4][10];
    ele[3][6] != ele[4][11];
    ele[3][6] != ele[4][6];
    ele[3][6] != ele[4][7];
    ele[3][6] != ele[4][8];
    ele[3][6] != ele[4][9];
    ele[3][6] != ele[5][10];
    ele[3][6] != ele[5][11];
    ele[3][6] != ele[5][6];
    ele[3][6] != ele[5][7];
    ele[3][6] != ele[5][8];
    ele[3][6] != ele[5][9];
    ele[3][6] != ele[6][6];
    ele[3][6] != ele[7][6];
    ele[3][6] != ele[8][6];
    ele[3][6] != ele[9][6];
    ele[3][7] != ele[10][7];
    ele[3][7] != ele[11][7];
    ele[3][7] != ele[12][7];
    ele[3][7] != ele[13][7];
    ele[3][7] != ele[14][7];
    ele[3][7] != ele[15][7];
    ele[3][7] != ele[16][7];
    ele[3][7] != ele[17][7];
    ele[3][7] != ele[18][7];
    ele[3][7] != ele[19][7];
    ele[3][7] != ele[20][7];
    ele[3][7] != ele[21][7];
    ele[3][7] != ele[22][7];
    ele[3][7] != ele[23][7];
    ele[3][7] != ele[24][7];
    ele[3][7] != ele[25][7];
    ele[3][7] != ele[26][7];
    ele[3][7] != ele[27][7];
    ele[3][7] != ele[28][7];
    ele[3][7] != ele[29][7];
    ele[3][7] != ele[3][10];
    ele[3][7] != ele[3][11];
    ele[3][7] != ele[3][12];
    ele[3][7] != ele[3][13];
    ele[3][7] != ele[3][14];
    ele[3][7] != ele[3][15];
    ele[3][7] != ele[3][16];
    ele[3][7] != ele[3][17];
    ele[3][7] != ele[3][18];
    ele[3][7] != ele[3][19];
    ele[3][7] != ele[3][20];
    ele[3][7] != ele[3][21];
    ele[3][7] != ele[3][22];
    ele[3][7] != ele[3][23];
    ele[3][7] != ele[3][24];
    ele[3][7] != ele[3][25];
    ele[3][7] != ele[3][26];
    ele[3][7] != ele[3][27];
    ele[3][7] != ele[3][28];
    ele[3][7] != ele[3][29];
    ele[3][7] != ele[3][30];
    ele[3][7] != ele[3][31];
    ele[3][7] != ele[3][32];
    ele[3][7] != ele[3][33];
    ele[3][7] != ele[3][34];
    ele[3][7] != ele[3][35];
    ele[3][7] != ele[3][8];
    ele[3][7] != ele[3][9];
    ele[3][7] != ele[30][7];
    ele[3][7] != ele[31][7];
    ele[3][7] != ele[32][7];
    ele[3][7] != ele[33][7];
    ele[3][7] != ele[34][7];
    ele[3][7] != ele[35][7];
    ele[3][7] != ele[4][10];
    ele[3][7] != ele[4][11];
    ele[3][7] != ele[4][6];
    ele[3][7] != ele[4][7];
    ele[3][7] != ele[4][8];
    ele[3][7] != ele[4][9];
    ele[3][7] != ele[5][10];
    ele[3][7] != ele[5][11];
    ele[3][7] != ele[5][6];
    ele[3][7] != ele[5][7];
    ele[3][7] != ele[5][8];
    ele[3][7] != ele[5][9];
    ele[3][7] != ele[6][7];
    ele[3][7] != ele[7][7];
    ele[3][7] != ele[8][7];
    ele[3][7] != ele[9][7];
    ele[3][8] != ele[10][8];
    ele[3][8] != ele[11][8];
    ele[3][8] != ele[12][8];
    ele[3][8] != ele[13][8];
    ele[3][8] != ele[14][8];
    ele[3][8] != ele[15][8];
    ele[3][8] != ele[16][8];
    ele[3][8] != ele[17][8];
    ele[3][8] != ele[18][8];
    ele[3][8] != ele[19][8];
    ele[3][8] != ele[20][8];
    ele[3][8] != ele[21][8];
    ele[3][8] != ele[22][8];
    ele[3][8] != ele[23][8];
    ele[3][8] != ele[24][8];
    ele[3][8] != ele[25][8];
    ele[3][8] != ele[26][8];
    ele[3][8] != ele[27][8];
    ele[3][8] != ele[28][8];
    ele[3][8] != ele[29][8];
    ele[3][8] != ele[3][10];
    ele[3][8] != ele[3][11];
    ele[3][8] != ele[3][12];
    ele[3][8] != ele[3][13];
    ele[3][8] != ele[3][14];
    ele[3][8] != ele[3][15];
    ele[3][8] != ele[3][16];
    ele[3][8] != ele[3][17];
    ele[3][8] != ele[3][18];
    ele[3][8] != ele[3][19];
    ele[3][8] != ele[3][20];
    ele[3][8] != ele[3][21];
    ele[3][8] != ele[3][22];
    ele[3][8] != ele[3][23];
    ele[3][8] != ele[3][24];
    ele[3][8] != ele[3][25];
    ele[3][8] != ele[3][26];
    ele[3][8] != ele[3][27];
    ele[3][8] != ele[3][28];
    ele[3][8] != ele[3][29];
    ele[3][8] != ele[3][30];
    ele[3][8] != ele[3][31];
    ele[3][8] != ele[3][32];
    ele[3][8] != ele[3][33];
    ele[3][8] != ele[3][34];
    ele[3][8] != ele[3][35];
    ele[3][8] != ele[3][9];
    ele[3][8] != ele[30][8];
    ele[3][8] != ele[31][8];
    ele[3][8] != ele[32][8];
    ele[3][8] != ele[33][8];
    ele[3][8] != ele[34][8];
    ele[3][8] != ele[35][8];
    ele[3][8] != ele[4][10];
    ele[3][8] != ele[4][11];
    ele[3][8] != ele[4][6];
    ele[3][8] != ele[4][7];
    ele[3][8] != ele[4][8];
    ele[3][8] != ele[4][9];
    ele[3][8] != ele[5][10];
    ele[3][8] != ele[5][11];
    ele[3][8] != ele[5][6];
    ele[3][8] != ele[5][7];
    ele[3][8] != ele[5][8];
    ele[3][8] != ele[5][9];
    ele[3][8] != ele[6][8];
    ele[3][8] != ele[7][8];
    ele[3][8] != ele[8][8];
    ele[3][8] != ele[9][8];
    ele[3][9] != ele[10][9];
    ele[3][9] != ele[11][9];
    ele[3][9] != ele[12][9];
    ele[3][9] != ele[13][9];
    ele[3][9] != ele[14][9];
    ele[3][9] != ele[15][9];
    ele[3][9] != ele[16][9];
    ele[3][9] != ele[17][9];
    ele[3][9] != ele[18][9];
    ele[3][9] != ele[19][9];
    ele[3][9] != ele[20][9];
    ele[3][9] != ele[21][9];
    ele[3][9] != ele[22][9];
    ele[3][9] != ele[23][9];
    ele[3][9] != ele[24][9];
    ele[3][9] != ele[25][9];
    ele[3][9] != ele[26][9];
    ele[3][9] != ele[27][9];
    ele[3][9] != ele[28][9];
    ele[3][9] != ele[29][9];
    ele[3][9] != ele[3][10];
    ele[3][9] != ele[3][11];
    ele[3][9] != ele[3][12];
    ele[3][9] != ele[3][13];
    ele[3][9] != ele[3][14];
    ele[3][9] != ele[3][15];
    ele[3][9] != ele[3][16];
    ele[3][9] != ele[3][17];
    ele[3][9] != ele[3][18];
    ele[3][9] != ele[3][19];
    ele[3][9] != ele[3][20];
    ele[3][9] != ele[3][21];
    ele[3][9] != ele[3][22];
    ele[3][9] != ele[3][23];
    ele[3][9] != ele[3][24];
    ele[3][9] != ele[3][25];
    ele[3][9] != ele[3][26];
    ele[3][9] != ele[3][27];
    ele[3][9] != ele[3][28];
    ele[3][9] != ele[3][29];
    ele[3][9] != ele[3][30];
    ele[3][9] != ele[3][31];
    ele[3][9] != ele[3][32];
    ele[3][9] != ele[3][33];
    ele[3][9] != ele[3][34];
    ele[3][9] != ele[3][35];
    ele[3][9] != ele[30][9];
    ele[3][9] != ele[31][9];
    ele[3][9] != ele[32][9];
    ele[3][9] != ele[33][9];
    ele[3][9] != ele[34][9];
    ele[3][9] != ele[35][9];
    ele[3][9] != ele[4][10];
    ele[3][9] != ele[4][11];
    ele[3][9] != ele[4][6];
    ele[3][9] != ele[4][7];
    ele[3][9] != ele[4][8];
    ele[3][9] != ele[4][9];
    ele[3][9] != ele[5][10];
    ele[3][9] != ele[5][11];
    ele[3][9] != ele[5][6];
    ele[3][9] != ele[5][7];
    ele[3][9] != ele[5][8];
    ele[3][9] != ele[5][9];
    ele[3][9] != ele[6][9];
    ele[3][9] != ele[7][9];
    ele[3][9] != ele[8][9];
    ele[3][9] != ele[9][9];
    ele[30][0] != ele[30][1];
    ele[30][0] != ele[30][10];
    ele[30][0] != ele[30][11];
    ele[30][0] != ele[30][12];
    ele[30][0] != ele[30][13];
    ele[30][0] != ele[30][14];
    ele[30][0] != ele[30][15];
    ele[30][0] != ele[30][16];
    ele[30][0] != ele[30][17];
    ele[30][0] != ele[30][18];
    ele[30][0] != ele[30][19];
    ele[30][0] != ele[30][2];
    ele[30][0] != ele[30][20];
    ele[30][0] != ele[30][21];
    ele[30][0] != ele[30][22];
    ele[30][0] != ele[30][23];
    ele[30][0] != ele[30][24];
    ele[30][0] != ele[30][25];
    ele[30][0] != ele[30][26];
    ele[30][0] != ele[30][27];
    ele[30][0] != ele[30][28];
    ele[30][0] != ele[30][29];
    ele[30][0] != ele[30][3];
    ele[30][0] != ele[30][30];
    ele[30][0] != ele[30][31];
    ele[30][0] != ele[30][32];
    ele[30][0] != ele[30][33];
    ele[30][0] != ele[30][34];
    ele[30][0] != ele[30][35];
    ele[30][0] != ele[30][4];
    ele[30][0] != ele[30][5];
    ele[30][0] != ele[30][6];
    ele[30][0] != ele[30][7];
    ele[30][0] != ele[30][8];
    ele[30][0] != ele[30][9];
    ele[30][0] != ele[31][0];
    ele[30][0] != ele[31][1];
    ele[30][0] != ele[31][2];
    ele[30][0] != ele[31][3];
    ele[30][0] != ele[31][4];
    ele[30][0] != ele[31][5];
    ele[30][0] != ele[32][0];
    ele[30][0] != ele[32][1];
    ele[30][0] != ele[32][2];
    ele[30][0] != ele[32][3];
    ele[30][0] != ele[32][4];
    ele[30][0] != ele[32][5];
    ele[30][0] != ele[33][0];
    ele[30][0] != ele[33][1];
    ele[30][0] != ele[33][2];
    ele[30][0] != ele[33][3];
    ele[30][0] != ele[33][4];
    ele[30][0] != ele[33][5];
    ele[30][0] != ele[34][0];
    ele[30][0] != ele[34][1];
    ele[30][0] != ele[34][2];
    ele[30][0] != ele[34][3];
    ele[30][0] != ele[34][4];
    ele[30][0] != ele[34][5];
    ele[30][0] != ele[35][0];
    ele[30][0] != ele[35][1];
    ele[30][0] != ele[35][2];
    ele[30][0] != ele[35][3];
    ele[30][0] != ele[35][4];
    ele[30][0] != ele[35][5];
    ele[30][1] != ele[30][10];
    ele[30][1] != ele[30][11];
    ele[30][1] != ele[30][12];
    ele[30][1] != ele[30][13];
    ele[30][1] != ele[30][14];
    ele[30][1] != ele[30][15];
    ele[30][1] != ele[30][16];
    ele[30][1] != ele[30][17];
    ele[30][1] != ele[30][18];
    ele[30][1] != ele[30][19];
    ele[30][1] != ele[30][2];
    ele[30][1] != ele[30][20];
    ele[30][1] != ele[30][21];
    ele[30][1] != ele[30][22];
    ele[30][1] != ele[30][23];
    ele[30][1] != ele[30][24];
    ele[30][1] != ele[30][25];
    ele[30][1] != ele[30][26];
    ele[30][1] != ele[30][27];
    ele[30][1] != ele[30][28];
    ele[30][1] != ele[30][29];
    ele[30][1] != ele[30][3];
    ele[30][1] != ele[30][30];
    ele[30][1] != ele[30][31];
    ele[30][1] != ele[30][32];
    ele[30][1] != ele[30][33];
    ele[30][1] != ele[30][34];
    ele[30][1] != ele[30][35];
    ele[30][1] != ele[30][4];
    ele[30][1] != ele[30][5];
    ele[30][1] != ele[30][6];
    ele[30][1] != ele[30][7];
    ele[30][1] != ele[30][8];
    ele[30][1] != ele[30][9];
    ele[30][1] != ele[31][0];
    ele[30][1] != ele[31][1];
    ele[30][1] != ele[31][2];
    ele[30][1] != ele[31][3];
    ele[30][1] != ele[31][4];
    ele[30][1] != ele[31][5];
    ele[30][1] != ele[32][0];
    ele[30][1] != ele[32][1];
    ele[30][1] != ele[32][2];
    ele[30][1] != ele[32][3];
    ele[30][1] != ele[32][4];
    ele[30][1] != ele[32][5];
    ele[30][1] != ele[33][0];
    ele[30][1] != ele[33][1];
    ele[30][1] != ele[33][2];
    ele[30][1] != ele[33][3];
    ele[30][1] != ele[33][4];
    ele[30][1] != ele[33][5];
    ele[30][1] != ele[34][0];
    ele[30][1] != ele[34][1];
    ele[30][1] != ele[34][2];
    ele[30][1] != ele[34][3];
    ele[30][1] != ele[34][4];
    ele[30][1] != ele[34][5];
    ele[30][1] != ele[35][0];
    ele[30][1] != ele[35][1];
    ele[30][1] != ele[35][2];
    ele[30][1] != ele[35][3];
    ele[30][1] != ele[35][4];
    ele[30][1] != ele[35][5];
    ele[30][10] != ele[30][11];
    ele[30][10] != ele[30][12];
    ele[30][10] != ele[30][13];
    ele[30][10] != ele[30][14];
    ele[30][10] != ele[30][15];
    ele[30][10] != ele[30][16];
    ele[30][10] != ele[30][17];
    ele[30][10] != ele[30][18];
    ele[30][10] != ele[30][19];
    ele[30][10] != ele[30][20];
    ele[30][10] != ele[30][21];
    ele[30][10] != ele[30][22];
    ele[30][10] != ele[30][23];
    ele[30][10] != ele[30][24];
    ele[30][10] != ele[30][25];
    ele[30][10] != ele[30][26];
    ele[30][10] != ele[30][27];
    ele[30][10] != ele[30][28];
    ele[30][10] != ele[30][29];
    ele[30][10] != ele[30][30];
    ele[30][10] != ele[30][31];
    ele[30][10] != ele[30][32];
    ele[30][10] != ele[30][33];
    ele[30][10] != ele[30][34];
    ele[30][10] != ele[30][35];
    ele[30][10] != ele[31][10];
    ele[30][10] != ele[31][11];
    ele[30][10] != ele[31][6];
    ele[30][10] != ele[31][7];
    ele[30][10] != ele[31][8];
    ele[30][10] != ele[31][9];
    ele[30][10] != ele[32][10];
    ele[30][10] != ele[32][11];
    ele[30][10] != ele[32][6];
    ele[30][10] != ele[32][7];
    ele[30][10] != ele[32][8];
    ele[30][10] != ele[32][9];
    ele[30][10] != ele[33][10];
    ele[30][10] != ele[33][11];
    ele[30][10] != ele[33][6];
    ele[30][10] != ele[33][7];
    ele[30][10] != ele[33][8];
    ele[30][10] != ele[33][9];
    ele[30][10] != ele[34][10];
    ele[30][10] != ele[34][11];
    ele[30][10] != ele[34][6];
    ele[30][10] != ele[34][7];
    ele[30][10] != ele[34][8];
    ele[30][10] != ele[34][9];
    ele[30][10] != ele[35][10];
    ele[30][10] != ele[35][11];
    ele[30][10] != ele[35][6];
    ele[30][10] != ele[35][7];
    ele[30][10] != ele[35][8];
    ele[30][10] != ele[35][9];
    ele[30][11] != ele[30][12];
    ele[30][11] != ele[30][13];
    ele[30][11] != ele[30][14];
    ele[30][11] != ele[30][15];
    ele[30][11] != ele[30][16];
    ele[30][11] != ele[30][17];
    ele[30][11] != ele[30][18];
    ele[30][11] != ele[30][19];
    ele[30][11] != ele[30][20];
    ele[30][11] != ele[30][21];
    ele[30][11] != ele[30][22];
    ele[30][11] != ele[30][23];
    ele[30][11] != ele[30][24];
    ele[30][11] != ele[30][25];
    ele[30][11] != ele[30][26];
    ele[30][11] != ele[30][27];
    ele[30][11] != ele[30][28];
    ele[30][11] != ele[30][29];
    ele[30][11] != ele[30][30];
    ele[30][11] != ele[30][31];
    ele[30][11] != ele[30][32];
    ele[30][11] != ele[30][33];
    ele[30][11] != ele[30][34];
    ele[30][11] != ele[30][35];
    ele[30][11] != ele[31][10];
    ele[30][11] != ele[31][11];
    ele[30][11] != ele[31][6];
    ele[30][11] != ele[31][7];
    ele[30][11] != ele[31][8];
    ele[30][11] != ele[31][9];
    ele[30][11] != ele[32][10];
    ele[30][11] != ele[32][11];
    ele[30][11] != ele[32][6];
    ele[30][11] != ele[32][7];
    ele[30][11] != ele[32][8];
    ele[30][11] != ele[32][9];
    ele[30][11] != ele[33][10];
    ele[30][11] != ele[33][11];
    ele[30][11] != ele[33][6];
    ele[30][11] != ele[33][7];
    ele[30][11] != ele[33][8];
    ele[30][11] != ele[33][9];
    ele[30][11] != ele[34][10];
    ele[30][11] != ele[34][11];
    ele[30][11] != ele[34][6];
    ele[30][11] != ele[34][7];
    ele[30][11] != ele[34][8];
    ele[30][11] != ele[34][9];
    ele[30][11] != ele[35][10];
    ele[30][11] != ele[35][11];
    ele[30][11] != ele[35][6];
    ele[30][11] != ele[35][7];
    ele[30][11] != ele[35][8];
    ele[30][11] != ele[35][9];
    ele[30][12] != ele[30][13];
    ele[30][12] != ele[30][14];
    ele[30][12] != ele[30][15];
    ele[30][12] != ele[30][16];
    ele[30][12] != ele[30][17];
    ele[30][12] != ele[30][18];
    ele[30][12] != ele[30][19];
    ele[30][12] != ele[30][20];
    ele[30][12] != ele[30][21];
    ele[30][12] != ele[30][22];
    ele[30][12] != ele[30][23];
    ele[30][12] != ele[30][24];
    ele[30][12] != ele[30][25];
    ele[30][12] != ele[30][26];
    ele[30][12] != ele[30][27];
    ele[30][12] != ele[30][28];
    ele[30][12] != ele[30][29];
    ele[30][12] != ele[30][30];
    ele[30][12] != ele[30][31];
    ele[30][12] != ele[30][32];
    ele[30][12] != ele[30][33];
    ele[30][12] != ele[30][34];
    ele[30][12] != ele[30][35];
    ele[30][12] != ele[31][12];
    ele[30][12] != ele[31][13];
    ele[30][12] != ele[31][14];
    ele[30][12] != ele[31][15];
    ele[30][12] != ele[31][16];
    ele[30][12] != ele[31][17];
    ele[30][12] != ele[32][12];
    ele[30][12] != ele[32][13];
    ele[30][12] != ele[32][14];
    ele[30][12] != ele[32][15];
    ele[30][12] != ele[32][16];
    ele[30][12] != ele[32][17];
    ele[30][12] != ele[33][12];
    ele[30][12] != ele[33][13];
    ele[30][12] != ele[33][14];
    ele[30][12] != ele[33][15];
    ele[30][12] != ele[33][16];
    ele[30][12] != ele[33][17];
    ele[30][12] != ele[34][12];
    ele[30][12] != ele[34][13];
    ele[30][12] != ele[34][14];
    ele[30][12] != ele[34][15];
    ele[30][12] != ele[34][16];
    ele[30][12] != ele[34][17];
    ele[30][12] != ele[35][12];
    ele[30][12] != ele[35][13];
    ele[30][12] != ele[35][14];
    ele[30][12] != ele[35][15];
    ele[30][12] != ele[35][16];
    ele[30][12] != ele[35][17];
    ele[30][13] != ele[30][14];
    ele[30][13] != ele[30][15];
    ele[30][13] != ele[30][16];
    ele[30][13] != ele[30][17];
    ele[30][13] != ele[30][18];
    ele[30][13] != ele[30][19];
    ele[30][13] != ele[30][20];
    ele[30][13] != ele[30][21];
    ele[30][13] != ele[30][22];
    ele[30][13] != ele[30][23];
    ele[30][13] != ele[30][24];
    ele[30][13] != ele[30][25];
    ele[30][13] != ele[30][26];
    ele[30][13] != ele[30][27];
    ele[30][13] != ele[30][28];
    ele[30][13] != ele[30][29];
    ele[30][13] != ele[30][30];
    ele[30][13] != ele[30][31];
    ele[30][13] != ele[30][32];
    ele[30][13] != ele[30][33];
    ele[30][13] != ele[30][34];
    ele[30][13] != ele[30][35];
    ele[30][13] != ele[31][12];
    ele[30][13] != ele[31][13];
    ele[30][13] != ele[31][14];
    ele[30][13] != ele[31][15];
    ele[30][13] != ele[31][16];
    ele[30][13] != ele[31][17];
    ele[30][13] != ele[32][12];
    ele[30][13] != ele[32][13];
    ele[30][13] != ele[32][14];
    ele[30][13] != ele[32][15];
    ele[30][13] != ele[32][16];
    ele[30][13] != ele[32][17];
    ele[30][13] != ele[33][12];
    ele[30][13] != ele[33][13];
    ele[30][13] != ele[33][14];
    ele[30][13] != ele[33][15];
    ele[30][13] != ele[33][16];
    ele[30][13] != ele[33][17];
    ele[30][13] != ele[34][12];
    ele[30][13] != ele[34][13];
    ele[30][13] != ele[34][14];
    ele[30][13] != ele[34][15];
    ele[30][13] != ele[34][16];
    ele[30][13] != ele[34][17];
    ele[30][13] != ele[35][12];
    ele[30][13] != ele[35][13];
    ele[30][13] != ele[35][14];
    ele[30][13] != ele[35][15];
    ele[30][13] != ele[35][16];
    ele[30][13] != ele[35][17];
    ele[30][14] != ele[30][15];
    ele[30][14] != ele[30][16];
    ele[30][14] != ele[30][17];
    ele[30][14] != ele[30][18];
    ele[30][14] != ele[30][19];
    ele[30][14] != ele[30][20];
    ele[30][14] != ele[30][21];
    ele[30][14] != ele[30][22];
    ele[30][14] != ele[30][23];
    ele[30][14] != ele[30][24];
    ele[30][14] != ele[30][25];
    ele[30][14] != ele[30][26];
    ele[30][14] != ele[30][27];
    ele[30][14] != ele[30][28];
    ele[30][14] != ele[30][29];
    ele[30][14] != ele[30][30];
    ele[30][14] != ele[30][31];
    ele[30][14] != ele[30][32];
    ele[30][14] != ele[30][33];
    ele[30][14] != ele[30][34];
    ele[30][14] != ele[30][35];
    ele[30][14] != ele[31][12];
    ele[30][14] != ele[31][13];
    ele[30][14] != ele[31][14];
    ele[30][14] != ele[31][15];
    ele[30][14] != ele[31][16];
    ele[30][14] != ele[31][17];
    ele[30][14] != ele[32][12];
    ele[30][14] != ele[32][13];
    ele[30][14] != ele[32][14];
    ele[30][14] != ele[32][15];
    ele[30][14] != ele[32][16];
    ele[30][14] != ele[32][17];
    ele[30][14] != ele[33][12];
    ele[30][14] != ele[33][13];
    ele[30][14] != ele[33][14];
    ele[30][14] != ele[33][15];
    ele[30][14] != ele[33][16];
    ele[30][14] != ele[33][17];
    ele[30][14] != ele[34][12];
    ele[30][14] != ele[34][13];
    ele[30][14] != ele[34][14];
    ele[30][14] != ele[34][15];
    ele[30][14] != ele[34][16];
    ele[30][14] != ele[34][17];
    ele[30][14] != ele[35][12];
    ele[30][14] != ele[35][13];
    ele[30][14] != ele[35][14];
    ele[30][14] != ele[35][15];
    ele[30][14] != ele[35][16];
    ele[30][14] != ele[35][17];
    ele[30][15] != ele[30][16];
    ele[30][15] != ele[30][17];
    ele[30][15] != ele[30][18];
    ele[30][15] != ele[30][19];
    ele[30][15] != ele[30][20];
    ele[30][15] != ele[30][21];
    ele[30][15] != ele[30][22];
    ele[30][15] != ele[30][23];
    ele[30][15] != ele[30][24];
    ele[30][15] != ele[30][25];
    ele[30][15] != ele[30][26];
    ele[30][15] != ele[30][27];
    ele[30][15] != ele[30][28];
    ele[30][15] != ele[30][29];
    ele[30][15] != ele[30][30];
    ele[30][15] != ele[30][31];
    ele[30][15] != ele[30][32];
    ele[30][15] != ele[30][33];
    ele[30][15] != ele[30][34];
    ele[30][15] != ele[30][35];
    ele[30][15] != ele[31][12];
    ele[30][15] != ele[31][13];
    ele[30][15] != ele[31][14];
    ele[30][15] != ele[31][15];
    ele[30][15] != ele[31][16];
    ele[30][15] != ele[31][17];
    ele[30][15] != ele[32][12];
    ele[30][15] != ele[32][13];
    ele[30][15] != ele[32][14];
    ele[30][15] != ele[32][15];
    ele[30][15] != ele[32][16];
    ele[30][15] != ele[32][17];
    ele[30][15] != ele[33][12];
    ele[30][15] != ele[33][13];
    ele[30][15] != ele[33][14];
    ele[30][15] != ele[33][15];
    ele[30][15] != ele[33][16];
    ele[30][15] != ele[33][17];
    ele[30][15] != ele[34][12];
    ele[30][15] != ele[34][13];
    ele[30][15] != ele[34][14];
    ele[30][15] != ele[34][15];
    ele[30][15] != ele[34][16];
    ele[30][15] != ele[34][17];
    ele[30][15] != ele[35][12];
    ele[30][15] != ele[35][13];
    ele[30][15] != ele[35][14];
    ele[30][15] != ele[35][15];
    ele[30][15] != ele[35][16];
    ele[30][15] != ele[35][17];
    ele[30][16] != ele[30][17];
    ele[30][16] != ele[30][18];
    ele[30][16] != ele[30][19];
    ele[30][16] != ele[30][20];
    ele[30][16] != ele[30][21];
    ele[30][16] != ele[30][22];
    ele[30][16] != ele[30][23];
    ele[30][16] != ele[30][24];
    ele[30][16] != ele[30][25];
    ele[30][16] != ele[30][26];
    ele[30][16] != ele[30][27];
    ele[30][16] != ele[30][28];
    ele[30][16] != ele[30][29];
    ele[30][16] != ele[30][30];
    ele[30][16] != ele[30][31];
    ele[30][16] != ele[30][32];
    ele[30][16] != ele[30][33];
    ele[30][16] != ele[30][34];
    ele[30][16] != ele[30][35];
    ele[30][16] != ele[31][12];
    ele[30][16] != ele[31][13];
    ele[30][16] != ele[31][14];
    ele[30][16] != ele[31][15];
    ele[30][16] != ele[31][16];
    ele[30][16] != ele[31][17];
    ele[30][16] != ele[32][12];
    ele[30][16] != ele[32][13];
    ele[30][16] != ele[32][14];
    ele[30][16] != ele[32][15];
    ele[30][16] != ele[32][16];
    ele[30][16] != ele[32][17];
    ele[30][16] != ele[33][12];
    ele[30][16] != ele[33][13];
    ele[30][16] != ele[33][14];
    ele[30][16] != ele[33][15];
    ele[30][16] != ele[33][16];
    ele[30][16] != ele[33][17];
    ele[30][16] != ele[34][12];
    ele[30][16] != ele[34][13];
    ele[30][16] != ele[34][14];
    ele[30][16] != ele[34][15];
    ele[30][16] != ele[34][16];
    ele[30][16] != ele[34][17];
    ele[30][16] != ele[35][12];
    ele[30][16] != ele[35][13];
    ele[30][16] != ele[35][14];
    ele[30][16] != ele[35][15];
    ele[30][16] != ele[35][16];
    ele[30][16] != ele[35][17];
    ele[30][17] != ele[30][18];
    ele[30][17] != ele[30][19];
    ele[30][17] != ele[30][20];
    ele[30][17] != ele[30][21];
    ele[30][17] != ele[30][22];
    ele[30][17] != ele[30][23];
    ele[30][17] != ele[30][24];
    ele[30][17] != ele[30][25];
    ele[30][17] != ele[30][26];
    ele[30][17] != ele[30][27];
    ele[30][17] != ele[30][28];
    ele[30][17] != ele[30][29];
    ele[30][17] != ele[30][30];
    ele[30][17] != ele[30][31];
    ele[30][17] != ele[30][32];
    ele[30][17] != ele[30][33];
    ele[30][17] != ele[30][34];
    ele[30][17] != ele[30][35];
    ele[30][17] != ele[31][12];
    ele[30][17] != ele[31][13];
    ele[30][17] != ele[31][14];
    ele[30][17] != ele[31][15];
    ele[30][17] != ele[31][16];
    ele[30][17] != ele[31][17];
    ele[30][17] != ele[32][12];
    ele[30][17] != ele[32][13];
    ele[30][17] != ele[32][14];
    ele[30][17] != ele[32][15];
    ele[30][17] != ele[32][16];
    ele[30][17] != ele[32][17];
    ele[30][17] != ele[33][12];
    ele[30][17] != ele[33][13];
    ele[30][17] != ele[33][14];
    ele[30][17] != ele[33][15];
    ele[30][17] != ele[33][16];
    ele[30][17] != ele[33][17];
    ele[30][17] != ele[34][12];
    ele[30][17] != ele[34][13];
    ele[30][17] != ele[34][14];
    ele[30][17] != ele[34][15];
    ele[30][17] != ele[34][16];
    ele[30][17] != ele[34][17];
    ele[30][17] != ele[35][12];
    ele[30][17] != ele[35][13];
    ele[30][17] != ele[35][14];
    ele[30][17] != ele[35][15];
    ele[30][17] != ele[35][16];
    ele[30][17] != ele[35][17];
    ele[30][18] != ele[30][19];
    ele[30][18] != ele[30][20];
    ele[30][18] != ele[30][21];
    ele[30][18] != ele[30][22];
    ele[30][18] != ele[30][23];
    ele[30][18] != ele[30][24];
    ele[30][18] != ele[30][25];
    ele[30][18] != ele[30][26];
    ele[30][18] != ele[30][27];
    ele[30][18] != ele[30][28];
    ele[30][18] != ele[30][29];
    ele[30][18] != ele[30][30];
    ele[30][18] != ele[30][31];
    ele[30][18] != ele[30][32];
    ele[30][18] != ele[30][33];
    ele[30][18] != ele[30][34];
    ele[30][18] != ele[30][35];
    ele[30][18] != ele[31][18];
    ele[30][18] != ele[31][19];
    ele[30][18] != ele[31][20];
    ele[30][18] != ele[31][21];
    ele[30][18] != ele[31][22];
    ele[30][18] != ele[31][23];
    ele[30][18] != ele[32][18];
    ele[30][18] != ele[32][19];
    ele[30][18] != ele[32][20];
    ele[30][18] != ele[32][21];
    ele[30][18] != ele[32][22];
    ele[30][18] != ele[32][23];
    ele[30][18] != ele[33][18];
    ele[30][18] != ele[33][19];
    ele[30][18] != ele[33][20];
    ele[30][18] != ele[33][21];
    ele[30][18] != ele[33][22];
    ele[30][18] != ele[33][23];
    ele[30][18] != ele[34][18];
    ele[30][18] != ele[34][19];
    ele[30][18] != ele[34][20];
    ele[30][18] != ele[34][21];
    ele[30][18] != ele[34][22];
    ele[30][18] != ele[34][23];
    ele[30][18] != ele[35][18];
    ele[30][18] != ele[35][19];
    ele[30][18] != ele[35][20];
    ele[30][18] != ele[35][21];
    ele[30][18] != ele[35][22];
    ele[30][18] != ele[35][23];
    ele[30][19] != ele[30][20];
    ele[30][19] != ele[30][21];
    ele[30][19] != ele[30][22];
    ele[30][19] != ele[30][23];
    ele[30][19] != ele[30][24];
    ele[30][19] != ele[30][25];
    ele[30][19] != ele[30][26];
    ele[30][19] != ele[30][27];
    ele[30][19] != ele[30][28];
    ele[30][19] != ele[30][29];
    ele[30][19] != ele[30][30];
    ele[30][19] != ele[30][31];
    ele[30][19] != ele[30][32];
    ele[30][19] != ele[30][33];
    ele[30][19] != ele[30][34];
    ele[30][19] != ele[30][35];
    ele[30][19] != ele[31][18];
    ele[30][19] != ele[31][19];
    ele[30][19] != ele[31][20];
    ele[30][19] != ele[31][21];
    ele[30][19] != ele[31][22];
    ele[30][19] != ele[31][23];
    ele[30][19] != ele[32][18];
    ele[30][19] != ele[32][19];
    ele[30][19] != ele[32][20];
    ele[30][19] != ele[32][21];
    ele[30][19] != ele[32][22];
    ele[30][19] != ele[32][23];
    ele[30][19] != ele[33][18];
    ele[30][19] != ele[33][19];
    ele[30][19] != ele[33][20];
    ele[30][19] != ele[33][21];
    ele[30][19] != ele[33][22];
    ele[30][19] != ele[33][23];
    ele[30][19] != ele[34][18];
    ele[30][19] != ele[34][19];
    ele[30][19] != ele[34][20];
    ele[30][19] != ele[34][21];
    ele[30][19] != ele[34][22];
    ele[30][19] != ele[34][23];
    ele[30][19] != ele[35][18];
    ele[30][19] != ele[35][19];
    ele[30][19] != ele[35][20];
    ele[30][19] != ele[35][21];
    ele[30][19] != ele[35][22];
    ele[30][19] != ele[35][23];
    ele[30][2] != ele[30][10];
    ele[30][2] != ele[30][11];
    ele[30][2] != ele[30][12];
    ele[30][2] != ele[30][13];
    ele[30][2] != ele[30][14];
    ele[30][2] != ele[30][15];
    ele[30][2] != ele[30][16];
    ele[30][2] != ele[30][17];
    ele[30][2] != ele[30][18];
    ele[30][2] != ele[30][19];
    ele[30][2] != ele[30][20];
    ele[30][2] != ele[30][21];
    ele[30][2] != ele[30][22];
    ele[30][2] != ele[30][23];
    ele[30][2] != ele[30][24];
    ele[30][2] != ele[30][25];
    ele[30][2] != ele[30][26];
    ele[30][2] != ele[30][27];
    ele[30][2] != ele[30][28];
    ele[30][2] != ele[30][29];
    ele[30][2] != ele[30][3];
    ele[30][2] != ele[30][30];
    ele[30][2] != ele[30][31];
    ele[30][2] != ele[30][32];
    ele[30][2] != ele[30][33];
    ele[30][2] != ele[30][34];
    ele[30][2] != ele[30][35];
    ele[30][2] != ele[30][4];
    ele[30][2] != ele[30][5];
    ele[30][2] != ele[30][6];
    ele[30][2] != ele[30][7];
    ele[30][2] != ele[30][8];
    ele[30][2] != ele[30][9];
    ele[30][2] != ele[31][0];
    ele[30][2] != ele[31][1];
    ele[30][2] != ele[31][2];
    ele[30][2] != ele[31][3];
    ele[30][2] != ele[31][4];
    ele[30][2] != ele[31][5];
    ele[30][2] != ele[32][0];
    ele[30][2] != ele[32][1];
    ele[30][2] != ele[32][2];
    ele[30][2] != ele[32][3];
    ele[30][2] != ele[32][4];
    ele[30][2] != ele[32][5];
    ele[30][2] != ele[33][0];
    ele[30][2] != ele[33][1];
    ele[30][2] != ele[33][2];
    ele[30][2] != ele[33][3];
    ele[30][2] != ele[33][4];
    ele[30][2] != ele[33][5];
    ele[30][2] != ele[34][0];
    ele[30][2] != ele[34][1];
    ele[30][2] != ele[34][2];
    ele[30][2] != ele[34][3];
    ele[30][2] != ele[34][4];
    ele[30][2] != ele[34][5];
    ele[30][2] != ele[35][0];
    ele[30][2] != ele[35][1];
    ele[30][2] != ele[35][2];
    ele[30][2] != ele[35][3];
    ele[30][2] != ele[35][4];
    ele[30][2] != ele[35][5];
    ele[30][20] != ele[30][21];
    ele[30][20] != ele[30][22];
    ele[30][20] != ele[30][23];
    ele[30][20] != ele[30][24];
    ele[30][20] != ele[30][25];
    ele[30][20] != ele[30][26];
    ele[30][20] != ele[30][27];
    ele[30][20] != ele[30][28];
    ele[30][20] != ele[30][29];
    ele[30][20] != ele[30][30];
    ele[30][20] != ele[30][31];
    ele[30][20] != ele[30][32];
    ele[30][20] != ele[30][33];
    ele[30][20] != ele[30][34];
    ele[30][20] != ele[30][35];
    ele[30][20] != ele[31][18];
    ele[30][20] != ele[31][19];
    ele[30][20] != ele[31][20];
    ele[30][20] != ele[31][21];
    ele[30][20] != ele[31][22];
    ele[30][20] != ele[31][23];
    ele[30][20] != ele[32][18];
    ele[30][20] != ele[32][19];
    ele[30][20] != ele[32][20];
    ele[30][20] != ele[32][21];
    ele[30][20] != ele[32][22];
    ele[30][20] != ele[32][23];
    ele[30][20] != ele[33][18];
    ele[30][20] != ele[33][19];
    ele[30][20] != ele[33][20];
    ele[30][20] != ele[33][21];
    ele[30][20] != ele[33][22];
    ele[30][20] != ele[33][23];
    ele[30][20] != ele[34][18];
    ele[30][20] != ele[34][19];
    ele[30][20] != ele[34][20];
    ele[30][20] != ele[34][21];
    ele[30][20] != ele[34][22];
    ele[30][20] != ele[34][23];
    ele[30][20] != ele[35][18];
    ele[30][20] != ele[35][19];
    ele[30][20] != ele[35][20];
    ele[30][20] != ele[35][21];
    ele[30][20] != ele[35][22];
    ele[30][20] != ele[35][23];
    ele[30][21] != ele[30][22];
    ele[30][21] != ele[30][23];
    ele[30][21] != ele[30][24];
    ele[30][21] != ele[30][25];
    ele[30][21] != ele[30][26];
    ele[30][21] != ele[30][27];
    ele[30][21] != ele[30][28];
    ele[30][21] != ele[30][29];
    ele[30][21] != ele[30][30];
    ele[30][21] != ele[30][31];
    ele[30][21] != ele[30][32];
    ele[30][21] != ele[30][33];
    ele[30][21] != ele[30][34];
    ele[30][21] != ele[30][35];
    ele[30][21] != ele[31][18];
    ele[30][21] != ele[31][19];
    ele[30][21] != ele[31][20];
    ele[30][21] != ele[31][21];
    ele[30][21] != ele[31][22];
    ele[30][21] != ele[31][23];
    ele[30][21] != ele[32][18];
    ele[30][21] != ele[32][19];
    ele[30][21] != ele[32][20];
    ele[30][21] != ele[32][21];
    ele[30][21] != ele[32][22];
    ele[30][21] != ele[32][23];
    ele[30][21] != ele[33][18];
    ele[30][21] != ele[33][19];
    ele[30][21] != ele[33][20];
    ele[30][21] != ele[33][21];
    ele[30][21] != ele[33][22];
    ele[30][21] != ele[33][23];
    ele[30][21] != ele[34][18];
    ele[30][21] != ele[34][19];
    ele[30][21] != ele[34][20];
    ele[30][21] != ele[34][21];
    ele[30][21] != ele[34][22];
    ele[30][21] != ele[34][23];
    ele[30][21] != ele[35][18];
    ele[30][21] != ele[35][19];
    ele[30][21] != ele[35][20];
    ele[30][21] != ele[35][21];
    ele[30][21] != ele[35][22];
    ele[30][21] != ele[35][23];
    ele[30][22] != ele[30][23];
    ele[30][22] != ele[30][24];
    ele[30][22] != ele[30][25];
    ele[30][22] != ele[30][26];
    ele[30][22] != ele[30][27];
    ele[30][22] != ele[30][28];
    ele[30][22] != ele[30][29];
    ele[30][22] != ele[30][30];
    ele[30][22] != ele[30][31];
    ele[30][22] != ele[30][32];
    ele[30][22] != ele[30][33];
    ele[30][22] != ele[30][34];
    ele[30][22] != ele[30][35];
    ele[30][22] != ele[31][18];
    ele[30][22] != ele[31][19];
    ele[30][22] != ele[31][20];
    ele[30][22] != ele[31][21];
    ele[30][22] != ele[31][22];
    ele[30][22] != ele[31][23];
    ele[30][22] != ele[32][18];
    ele[30][22] != ele[32][19];
    ele[30][22] != ele[32][20];
    ele[30][22] != ele[32][21];
    ele[30][22] != ele[32][22];
    ele[30][22] != ele[32][23];
    ele[30][22] != ele[33][18];
    ele[30][22] != ele[33][19];
    ele[30][22] != ele[33][20];
    ele[30][22] != ele[33][21];
    ele[30][22] != ele[33][22];
    ele[30][22] != ele[33][23];
    ele[30][22] != ele[34][18];
    ele[30][22] != ele[34][19];
    ele[30][22] != ele[34][20];
    ele[30][22] != ele[34][21];
    ele[30][22] != ele[34][22];
    ele[30][22] != ele[34][23];
    ele[30][22] != ele[35][18];
    ele[30][22] != ele[35][19];
    ele[30][22] != ele[35][20];
    ele[30][22] != ele[35][21];
    ele[30][22] != ele[35][22];
    ele[30][22] != ele[35][23];
    ele[30][23] != ele[30][24];
    ele[30][23] != ele[30][25];
    ele[30][23] != ele[30][26];
    ele[30][23] != ele[30][27];
    ele[30][23] != ele[30][28];
    ele[30][23] != ele[30][29];
    ele[30][23] != ele[30][30];
    ele[30][23] != ele[30][31];
    ele[30][23] != ele[30][32];
    ele[30][23] != ele[30][33];
    ele[30][23] != ele[30][34];
    ele[30][23] != ele[30][35];
    ele[30][23] != ele[31][18];
    ele[30][23] != ele[31][19];
    ele[30][23] != ele[31][20];
    ele[30][23] != ele[31][21];
    ele[30][23] != ele[31][22];
    ele[30][23] != ele[31][23];
    ele[30][23] != ele[32][18];
    ele[30][23] != ele[32][19];
    ele[30][23] != ele[32][20];
    ele[30][23] != ele[32][21];
    ele[30][23] != ele[32][22];
    ele[30][23] != ele[32][23];
    ele[30][23] != ele[33][18];
    ele[30][23] != ele[33][19];
    ele[30][23] != ele[33][20];
    ele[30][23] != ele[33][21];
    ele[30][23] != ele[33][22];
    ele[30][23] != ele[33][23];
    ele[30][23] != ele[34][18];
    ele[30][23] != ele[34][19];
    ele[30][23] != ele[34][20];
    ele[30][23] != ele[34][21];
    ele[30][23] != ele[34][22];
    ele[30][23] != ele[34][23];
    ele[30][23] != ele[35][18];
    ele[30][23] != ele[35][19];
    ele[30][23] != ele[35][20];
    ele[30][23] != ele[35][21];
    ele[30][23] != ele[35][22];
    ele[30][23] != ele[35][23];
    ele[30][24] != ele[30][25];
    ele[30][24] != ele[30][26];
    ele[30][24] != ele[30][27];
    ele[30][24] != ele[30][28];
    ele[30][24] != ele[30][29];
    ele[30][24] != ele[30][30];
    ele[30][24] != ele[30][31];
    ele[30][24] != ele[30][32];
    ele[30][24] != ele[30][33];
    ele[30][24] != ele[30][34];
    ele[30][24] != ele[30][35];
    ele[30][24] != ele[31][24];
    ele[30][24] != ele[31][25];
    ele[30][24] != ele[31][26];
    ele[30][24] != ele[31][27];
    ele[30][24] != ele[31][28];
    ele[30][24] != ele[31][29];
    ele[30][24] != ele[32][24];
    ele[30][24] != ele[32][25];
    ele[30][24] != ele[32][26];
    ele[30][24] != ele[32][27];
    ele[30][24] != ele[32][28];
    ele[30][24] != ele[32][29];
    ele[30][24] != ele[33][24];
    ele[30][24] != ele[33][25];
    ele[30][24] != ele[33][26];
    ele[30][24] != ele[33][27];
    ele[30][24] != ele[33][28];
    ele[30][24] != ele[33][29];
    ele[30][24] != ele[34][24];
    ele[30][24] != ele[34][25];
    ele[30][24] != ele[34][26];
    ele[30][24] != ele[34][27];
    ele[30][24] != ele[34][28];
    ele[30][24] != ele[34][29];
    ele[30][24] != ele[35][24];
    ele[30][24] != ele[35][25];
    ele[30][24] != ele[35][26];
    ele[30][24] != ele[35][27];
    ele[30][24] != ele[35][28];
    ele[30][24] != ele[35][29];
    ele[30][25] != ele[30][26];
    ele[30][25] != ele[30][27];
    ele[30][25] != ele[30][28];
    ele[30][25] != ele[30][29];
    ele[30][25] != ele[30][30];
    ele[30][25] != ele[30][31];
    ele[30][25] != ele[30][32];
    ele[30][25] != ele[30][33];
    ele[30][25] != ele[30][34];
    ele[30][25] != ele[30][35];
    ele[30][25] != ele[31][24];
    ele[30][25] != ele[31][25];
    ele[30][25] != ele[31][26];
    ele[30][25] != ele[31][27];
    ele[30][25] != ele[31][28];
    ele[30][25] != ele[31][29];
    ele[30][25] != ele[32][24];
    ele[30][25] != ele[32][25];
    ele[30][25] != ele[32][26];
    ele[30][25] != ele[32][27];
    ele[30][25] != ele[32][28];
    ele[30][25] != ele[32][29];
    ele[30][25] != ele[33][24];
    ele[30][25] != ele[33][25];
    ele[30][25] != ele[33][26];
    ele[30][25] != ele[33][27];
    ele[30][25] != ele[33][28];
    ele[30][25] != ele[33][29];
    ele[30][25] != ele[34][24];
    ele[30][25] != ele[34][25];
    ele[30][25] != ele[34][26];
    ele[30][25] != ele[34][27];
    ele[30][25] != ele[34][28];
    ele[30][25] != ele[34][29];
    ele[30][25] != ele[35][24];
    ele[30][25] != ele[35][25];
    ele[30][25] != ele[35][26];
    ele[30][25] != ele[35][27];
    ele[30][25] != ele[35][28];
    ele[30][25] != ele[35][29];
    ele[30][26] != ele[30][27];
    ele[30][26] != ele[30][28];
    ele[30][26] != ele[30][29];
    ele[30][26] != ele[30][30];
    ele[30][26] != ele[30][31];
    ele[30][26] != ele[30][32];
    ele[30][26] != ele[30][33];
    ele[30][26] != ele[30][34];
    ele[30][26] != ele[30][35];
    ele[30][26] != ele[31][24];
    ele[30][26] != ele[31][25];
    ele[30][26] != ele[31][26];
    ele[30][26] != ele[31][27];
    ele[30][26] != ele[31][28];
    ele[30][26] != ele[31][29];
    ele[30][26] != ele[32][24];
    ele[30][26] != ele[32][25];
    ele[30][26] != ele[32][26];
    ele[30][26] != ele[32][27];
    ele[30][26] != ele[32][28];
    ele[30][26] != ele[32][29];
    ele[30][26] != ele[33][24];
    ele[30][26] != ele[33][25];
    ele[30][26] != ele[33][26];
    ele[30][26] != ele[33][27];
    ele[30][26] != ele[33][28];
    ele[30][26] != ele[33][29];
    ele[30][26] != ele[34][24];
    ele[30][26] != ele[34][25];
    ele[30][26] != ele[34][26];
    ele[30][26] != ele[34][27];
    ele[30][26] != ele[34][28];
    ele[30][26] != ele[34][29];
    ele[30][26] != ele[35][24];
    ele[30][26] != ele[35][25];
    ele[30][26] != ele[35][26];
    ele[30][26] != ele[35][27];
    ele[30][26] != ele[35][28];
    ele[30][26] != ele[35][29];
    ele[30][27] != ele[30][28];
    ele[30][27] != ele[30][29];
    ele[30][27] != ele[30][30];
    ele[30][27] != ele[30][31];
    ele[30][27] != ele[30][32];
    ele[30][27] != ele[30][33];
    ele[30][27] != ele[30][34];
    ele[30][27] != ele[30][35];
    ele[30][27] != ele[31][24];
    ele[30][27] != ele[31][25];
    ele[30][27] != ele[31][26];
    ele[30][27] != ele[31][27];
    ele[30][27] != ele[31][28];
    ele[30][27] != ele[31][29];
    ele[30][27] != ele[32][24];
    ele[30][27] != ele[32][25];
    ele[30][27] != ele[32][26];
    ele[30][27] != ele[32][27];
    ele[30][27] != ele[32][28];
    ele[30][27] != ele[32][29];
    ele[30][27] != ele[33][24];
    ele[30][27] != ele[33][25];
    ele[30][27] != ele[33][26];
    ele[30][27] != ele[33][27];
    ele[30][27] != ele[33][28];
    ele[30][27] != ele[33][29];
    ele[30][27] != ele[34][24];
    ele[30][27] != ele[34][25];
    ele[30][27] != ele[34][26];
    ele[30][27] != ele[34][27];
    ele[30][27] != ele[34][28];
    ele[30][27] != ele[34][29];
    ele[30][27] != ele[35][24];
    ele[30][27] != ele[35][25];
    ele[30][27] != ele[35][26];
    ele[30][27] != ele[35][27];
    ele[30][27] != ele[35][28];
    ele[30][27] != ele[35][29];
    ele[30][28] != ele[30][29];
    ele[30][28] != ele[30][30];
    ele[30][28] != ele[30][31];
    ele[30][28] != ele[30][32];
    ele[30][28] != ele[30][33];
    ele[30][28] != ele[30][34];
    ele[30][28] != ele[30][35];
    ele[30][28] != ele[31][24];
    ele[30][28] != ele[31][25];
    ele[30][28] != ele[31][26];
    ele[30][28] != ele[31][27];
    ele[30][28] != ele[31][28];
    ele[30][28] != ele[31][29];
    ele[30][28] != ele[32][24];
    ele[30][28] != ele[32][25];
    ele[30][28] != ele[32][26];
    ele[30][28] != ele[32][27];
    ele[30][28] != ele[32][28];
    ele[30][28] != ele[32][29];
    ele[30][28] != ele[33][24];
    ele[30][28] != ele[33][25];
    ele[30][28] != ele[33][26];
    ele[30][28] != ele[33][27];
    ele[30][28] != ele[33][28];
    ele[30][28] != ele[33][29];
    ele[30][28] != ele[34][24];
    ele[30][28] != ele[34][25];
    ele[30][28] != ele[34][26];
    ele[30][28] != ele[34][27];
    ele[30][28] != ele[34][28];
    ele[30][28] != ele[34][29];
    ele[30][28] != ele[35][24];
    ele[30][28] != ele[35][25];
    ele[30][28] != ele[35][26];
    ele[30][28] != ele[35][27];
    ele[30][28] != ele[35][28];
    ele[30][28] != ele[35][29];
    ele[30][29] != ele[30][30];
    ele[30][29] != ele[30][31];
    ele[30][29] != ele[30][32];
    ele[30][29] != ele[30][33];
    ele[30][29] != ele[30][34];
    ele[30][29] != ele[30][35];
    ele[30][29] != ele[31][24];
    ele[30][29] != ele[31][25];
    ele[30][29] != ele[31][26];
    ele[30][29] != ele[31][27];
    ele[30][29] != ele[31][28];
    ele[30][29] != ele[31][29];
    ele[30][29] != ele[32][24];
    ele[30][29] != ele[32][25];
    ele[30][29] != ele[32][26];
    ele[30][29] != ele[32][27];
    ele[30][29] != ele[32][28];
    ele[30][29] != ele[32][29];
    ele[30][29] != ele[33][24];
    ele[30][29] != ele[33][25];
    ele[30][29] != ele[33][26];
    ele[30][29] != ele[33][27];
    ele[30][29] != ele[33][28];
    ele[30][29] != ele[33][29];
    ele[30][29] != ele[34][24];
    ele[30][29] != ele[34][25];
    ele[30][29] != ele[34][26];
    ele[30][29] != ele[34][27];
    ele[30][29] != ele[34][28];
    ele[30][29] != ele[34][29];
    ele[30][29] != ele[35][24];
    ele[30][29] != ele[35][25];
    ele[30][29] != ele[35][26];
    ele[30][29] != ele[35][27];
    ele[30][29] != ele[35][28];
    ele[30][29] != ele[35][29];
    ele[30][3] != ele[30][10];
    ele[30][3] != ele[30][11];
    ele[30][3] != ele[30][12];
    ele[30][3] != ele[30][13];
    ele[30][3] != ele[30][14];
    ele[30][3] != ele[30][15];
    ele[30][3] != ele[30][16];
    ele[30][3] != ele[30][17];
    ele[30][3] != ele[30][18];
    ele[30][3] != ele[30][19];
    ele[30][3] != ele[30][20];
    ele[30][3] != ele[30][21];
    ele[30][3] != ele[30][22];
    ele[30][3] != ele[30][23];
    ele[30][3] != ele[30][24];
    ele[30][3] != ele[30][25];
    ele[30][3] != ele[30][26];
    ele[30][3] != ele[30][27];
    ele[30][3] != ele[30][28];
    ele[30][3] != ele[30][29];
    ele[30][3] != ele[30][30];
    ele[30][3] != ele[30][31];
    ele[30][3] != ele[30][32];
    ele[30][3] != ele[30][33];
    ele[30][3] != ele[30][34];
    ele[30][3] != ele[30][35];
    ele[30][3] != ele[30][4];
    ele[30][3] != ele[30][5];
    ele[30][3] != ele[30][6];
    ele[30][3] != ele[30][7];
    ele[30][3] != ele[30][8];
    ele[30][3] != ele[30][9];
    ele[30][3] != ele[31][0];
    ele[30][3] != ele[31][1];
    ele[30][3] != ele[31][2];
    ele[30][3] != ele[31][3];
    ele[30][3] != ele[31][4];
    ele[30][3] != ele[31][5];
    ele[30][3] != ele[32][0];
    ele[30][3] != ele[32][1];
    ele[30][3] != ele[32][2];
    ele[30][3] != ele[32][3];
    ele[30][3] != ele[32][4];
    ele[30][3] != ele[32][5];
    ele[30][3] != ele[33][0];
    ele[30][3] != ele[33][1];
    ele[30][3] != ele[33][2];
    ele[30][3] != ele[33][3];
    ele[30][3] != ele[33][4];
    ele[30][3] != ele[33][5];
    ele[30][3] != ele[34][0];
    ele[30][3] != ele[34][1];
    ele[30][3] != ele[34][2];
    ele[30][3] != ele[34][3];
    ele[30][3] != ele[34][4];
    ele[30][3] != ele[34][5];
    ele[30][3] != ele[35][0];
    ele[30][3] != ele[35][1];
    ele[30][3] != ele[35][2];
    ele[30][3] != ele[35][3];
    ele[30][3] != ele[35][4];
    ele[30][3] != ele[35][5];
    ele[30][30] != ele[30][31];
    ele[30][30] != ele[30][32];
    ele[30][30] != ele[30][33];
    ele[30][30] != ele[30][34];
    ele[30][30] != ele[30][35];
    ele[30][30] != ele[31][30];
    ele[30][30] != ele[31][31];
    ele[30][30] != ele[31][32];
    ele[30][30] != ele[31][33];
    ele[30][30] != ele[31][34];
    ele[30][30] != ele[31][35];
    ele[30][30] != ele[32][30];
    ele[30][30] != ele[32][31];
    ele[30][30] != ele[32][32];
    ele[30][30] != ele[32][33];
    ele[30][30] != ele[32][34];
    ele[30][30] != ele[32][35];
    ele[30][30] != ele[33][30];
    ele[30][30] != ele[33][31];
    ele[30][30] != ele[33][32];
    ele[30][30] != ele[33][33];
    ele[30][30] != ele[33][34];
    ele[30][30] != ele[33][35];
    ele[30][30] != ele[34][30];
    ele[30][30] != ele[34][31];
    ele[30][30] != ele[34][32];
    ele[30][30] != ele[34][33];
    ele[30][30] != ele[34][34];
    ele[30][30] != ele[34][35];
    ele[30][30] != ele[35][30];
    ele[30][30] != ele[35][31];
    ele[30][30] != ele[35][32];
    ele[30][30] != ele[35][33];
    ele[30][30] != ele[35][34];
    ele[30][30] != ele[35][35];
    ele[30][31] != ele[30][32];
    ele[30][31] != ele[30][33];
    ele[30][31] != ele[30][34];
    ele[30][31] != ele[30][35];
    ele[30][31] != ele[31][30];
    ele[30][31] != ele[31][31];
    ele[30][31] != ele[31][32];
    ele[30][31] != ele[31][33];
    ele[30][31] != ele[31][34];
    ele[30][31] != ele[31][35];
    ele[30][31] != ele[32][30];
    ele[30][31] != ele[32][31];
    ele[30][31] != ele[32][32];
    ele[30][31] != ele[32][33];
    ele[30][31] != ele[32][34];
    ele[30][31] != ele[32][35];
    ele[30][31] != ele[33][30];
    ele[30][31] != ele[33][31];
    ele[30][31] != ele[33][32];
    ele[30][31] != ele[33][33];
    ele[30][31] != ele[33][34];
    ele[30][31] != ele[33][35];
    ele[30][31] != ele[34][30];
    ele[30][31] != ele[34][31];
    ele[30][31] != ele[34][32];
    ele[30][31] != ele[34][33];
    ele[30][31] != ele[34][34];
    ele[30][31] != ele[34][35];
    ele[30][31] != ele[35][30];
    ele[30][31] != ele[35][31];
    ele[30][31] != ele[35][32];
    ele[30][31] != ele[35][33];
    ele[30][31] != ele[35][34];
    ele[30][31] != ele[35][35];
    ele[30][32] != ele[30][33];
    ele[30][32] != ele[30][34];
    ele[30][32] != ele[30][35];
    ele[30][32] != ele[31][30];
    ele[30][32] != ele[31][31];
    ele[30][32] != ele[31][32];
    ele[30][32] != ele[31][33];
    ele[30][32] != ele[31][34];
    ele[30][32] != ele[31][35];
    ele[30][32] != ele[32][30];
    ele[30][32] != ele[32][31];
    ele[30][32] != ele[32][32];
    ele[30][32] != ele[32][33];
    ele[30][32] != ele[32][34];
    ele[30][32] != ele[32][35];
    ele[30][32] != ele[33][30];
    ele[30][32] != ele[33][31];
    ele[30][32] != ele[33][32];
    ele[30][32] != ele[33][33];
    ele[30][32] != ele[33][34];
    ele[30][32] != ele[33][35];
    ele[30][32] != ele[34][30];
    ele[30][32] != ele[34][31];
    ele[30][32] != ele[34][32];
    ele[30][32] != ele[34][33];
    ele[30][32] != ele[34][34];
    ele[30][32] != ele[34][35];
    ele[30][32] != ele[35][30];
    ele[30][32] != ele[35][31];
    ele[30][32] != ele[35][32];
    ele[30][32] != ele[35][33];
    ele[30][32] != ele[35][34];
    ele[30][32] != ele[35][35];
    ele[30][33] != ele[30][34];
    ele[30][33] != ele[30][35];
    ele[30][33] != ele[31][30];
    ele[30][33] != ele[31][31];
    ele[30][33] != ele[31][32];
    ele[30][33] != ele[31][33];
    ele[30][33] != ele[31][34];
    ele[30][33] != ele[31][35];
    ele[30][33] != ele[32][30];
    ele[30][33] != ele[32][31];
    ele[30][33] != ele[32][32];
    ele[30][33] != ele[32][33];
    ele[30][33] != ele[32][34];
    ele[30][33] != ele[32][35];
    ele[30][33] != ele[33][30];
    ele[30][33] != ele[33][31];
    ele[30][33] != ele[33][32];
    ele[30][33] != ele[33][33];
    ele[30][33] != ele[33][34];
    ele[30][33] != ele[33][35];
    ele[30][33] != ele[34][30];
    ele[30][33] != ele[34][31];
    ele[30][33] != ele[34][32];
    ele[30][33] != ele[34][33];
    ele[30][33] != ele[34][34];
    ele[30][33] != ele[34][35];
    ele[30][33] != ele[35][30];
    ele[30][33] != ele[35][31];
    ele[30][33] != ele[35][32];
    ele[30][33] != ele[35][33];
    ele[30][33] != ele[35][34];
    ele[30][33] != ele[35][35];
    ele[30][34] != ele[30][35];
    ele[30][34] != ele[31][30];
    ele[30][34] != ele[31][31];
    ele[30][34] != ele[31][32];
    ele[30][34] != ele[31][33];
    ele[30][34] != ele[31][34];
    ele[30][34] != ele[31][35];
    ele[30][34] != ele[32][30];
    ele[30][34] != ele[32][31];
    ele[30][34] != ele[32][32];
    ele[30][34] != ele[32][33];
    ele[30][34] != ele[32][34];
    ele[30][34] != ele[32][35];
    ele[30][34] != ele[33][30];
    ele[30][34] != ele[33][31];
    ele[30][34] != ele[33][32];
    ele[30][34] != ele[33][33];
    ele[30][34] != ele[33][34];
    ele[30][34] != ele[33][35];
    ele[30][34] != ele[34][30];
    ele[30][34] != ele[34][31];
    ele[30][34] != ele[34][32];
    ele[30][34] != ele[34][33];
    ele[30][34] != ele[34][34];
    ele[30][34] != ele[34][35];
    ele[30][34] != ele[35][30];
    ele[30][34] != ele[35][31];
    ele[30][34] != ele[35][32];
    ele[30][34] != ele[35][33];
    ele[30][34] != ele[35][34];
    ele[30][34] != ele[35][35];
    ele[30][35] != ele[31][30];
    ele[30][35] != ele[31][31];
    ele[30][35] != ele[31][32];
    ele[30][35] != ele[31][33];
    ele[30][35] != ele[31][34];
    ele[30][35] != ele[31][35];
    ele[30][35] != ele[32][30];
    ele[30][35] != ele[32][31];
    ele[30][35] != ele[32][32];
    ele[30][35] != ele[32][33];
    ele[30][35] != ele[32][34];
    ele[30][35] != ele[32][35];
    ele[30][35] != ele[33][30];
    ele[30][35] != ele[33][31];
    ele[30][35] != ele[33][32];
    ele[30][35] != ele[33][33];
    ele[30][35] != ele[33][34];
    ele[30][35] != ele[33][35];
    ele[30][35] != ele[34][30];
    ele[30][35] != ele[34][31];
    ele[30][35] != ele[34][32];
    ele[30][35] != ele[34][33];
    ele[30][35] != ele[34][34];
    ele[30][35] != ele[34][35];
    ele[30][35] != ele[35][30];
    ele[30][35] != ele[35][31];
    ele[30][35] != ele[35][32];
    ele[30][35] != ele[35][33];
    ele[30][35] != ele[35][34];
    ele[30][35] != ele[35][35];
    ele[30][4] != ele[30][10];
    ele[30][4] != ele[30][11];
    ele[30][4] != ele[30][12];
    ele[30][4] != ele[30][13];
    ele[30][4] != ele[30][14];
    ele[30][4] != ele[30][15];
    ele[30][4] != ele[30][16];
    ele[30][4] != ele[30][17];
    ele[30][4] != ele[30][18];
    ele[30][4] != ele[30][19];
    ele[30][4] != ele[30][20];
    ele[30][4] != ele[30][21];
    ele[30][4] != ele[30][22];
    ele[30][4] != ele[30][23];
    ele[30][4] != ele[30][24];
    ele[30][4] != ele[30][25];
    ele[30][4] != ele[30][26];
    ele[30][4] != ele[30][27];
    ele[30][4] != ele[30][28];
    ele[30][4] != ele[30][29];
    ele[30][4] != ele[30][30];
    ele[30][4] != ele[30][31];
    ele[30][4] != ele[30][32];
    ele[30][4] != ele[30][33];
    ele[30][4] != ele[30][34];
    ele[30][4] != ele[30][35];
    ele[30][4] != ele[30][5];
    ele[30][4] != ele[30][6];
    ele[30][4] != ele[30][7];
    ele[30][4] != ele[30][8];
    ele[30][4] != ele[30][9];
    ele[30][4] != ele[31][0];
    ele[30][4] != ele[31][1];
    ele[30][4] != ele[31][2];
    ele[30][4] != ele[31][3];
    ele[30][4] != ele[31][4];
    ele[30][4] != ele[31][5];
    ele[30][4] != ele[32][0];
    ele[30][4] != ele[32][1];
    ele[30][4] != ele[32][2];
    ele[30][4] != ele[32][3];
    ele[30][4] != ele[32][4];
    ele[30][4] != ele[32][5];
    ele[30][4] != ele[33][0];
    ele[30][4] != ele[33][1];
    ele[30][4] != ele[33][2];
    ele[30][4] != ele[33][3];
    ele[30][4] != ele[33][4];
    ele[30][4] != ele[33][5];
    ele[30][4] != ele[34][0];
    ele[30][4] != ele[34][1];
    ele[30][4] != ele[34][2];
    ele[30][4] != ele[34][3];
    ele[30][4] != ele[34][4];
    ele[30][4] != ele[34][5];
    ele[30][4] != ele[35][0];
    ele[30][4] != ele[35][1];
    ele[30][4] != ele[35][2];
    ele[30][4] != ele[35][3];
    ele[30][4] != ele[35][4];
    ele[30][4] != ele[35][5];
    ele[30][5] != ele[30][10];
    ele[30][5] != ele[30][11];
    ele[30][5] != ele[30][12];
    ele[30][5] != ele[30][13];
    ele[30][5] != ele[30][14];
    ele[30][5] != ele[30][15];
    ele[30][5] != ele[30][16];
    ele[30][5] != ele[30][17];
    ele[30][5] != ele[30][18];
    ele[30][5] != ele[30][19];
    ele[30][5] != ele[30][20];
    ele[30][5] != ele[30][21];
    ele[30][5] != ele[30][22];
    ele[30][5] != ele[30][23];
    ele[30][5] != ele[30][24];
    ele[30][5] != ele[30][25];
    ele[30][5] != ele[30][26];
    ele[30][5] != ele[30][27];
    ele[30][5] != ele[30][28];
    ele[30][5] != ele[30][29];
    ele[30][5] != ele[30][30];
    ele[30][5] != ele[30][31];
    ele[30][5] != ele[30][32];
    ele[30][5] != ele[30][33];
    ele[30][5] != ele[30][34];
    ele[30][5] != ele[30][35];
    ele[30][5] != ele[30][6];
    ele[30][5] != ele[30][7];
    ele[30][5] != ele[30][8];
    ele[30][5] != ele[30][9];
    ele[30][5] != ele[31][0];
    ele[30][5] != ele[31][1];
    ele[30][5] != ele[31][2];
    ele[30][5] != ele[31][3];
    ele[30][5] != ele[31][4];
    ele[30][5] != ele[31][5];
    ele[30][5] != ele[32][0];
    ele[30][5] != ele[32][1];
    ele[30][5] != ele[32][2];
    ele[30][5] != ele[32][3];
    ele[30][5] != ele[32][4];
    ele[30][5] != ele[32][5];
    ele[30][5] != ele[33][0];
    ele[30][5] != ele[33][1];
    ele[30][5] != ele[33][2];
    ele[30][5] != ele[33][3];
    ele[30][5] != ele[33][4];
    ele[30][5] != ele[33][5];
    ele[30][5] != ele[34][0];
    ele[30][5] != ele[34][1];
    ele[30][5] != ele[34][2];
    ele[30][5] != ele[34][3];
    ele[30][5] != ele[34][4];
    ele[30][5] != ele[34][5];
    ele[30][5] != ele[35][0];
    ele[30][5] != ele[35][1];
    ele[30][5] != ele[35][2];
    ele[30][5] != ele[35][3];
    ele[30][5] != ele[35][4];
    ele[30][5] != ele[35][5];
    ele[30][6] != ele[30][10];
    ele[30][6] != ele[30][11];
    ele[30][6] != ele[30][12];
    ele[30][6] != ele[30][13];
    ele[30][6] != ele[30][14];
    ele[30][6] != ele[30][15];
    ele[30][6] != ele[30][16];
    ele[30][6] != ele[30][17];
    ele[30][6] != ele[30][18];
    ele[30][6] != ele[30][19];
    ele[30][6] != ele[30][20];
    ele[30][6] != ele[30][21];
    ele[30][6] != ele[30][22];
    ele[30][6] != ele[30][23];
    ele[30][6] != ele[30][24];
    ele[30][6] != ele[30][25];
    ele[30][6] != ele[30][26];
    ele[30][6] != ele[30][27];
    ele[30][6] != ele[30][28];
    ele[30][6] != ele[30][29];
    ele[30][6] != ele[30][30];
    ele[30][6] != ele[30][31];
    ele[30][6] != ele[30][32];
    ele[30][6] != ele[30][33];
    ele[30][6] != ele[30][34];
    ele[30][6] != ele[30][35];
    ele[30][6] != ele[30][7];
    ele[30][6] != ele[30][8];
    ele[30][6] != ele[30][9];
    ele[30][6] != ele[31][10];
    ele[30][6] != ele[31][11];
    ele[30][6] != ele[31][6];
    ele[30][6] != ele[31][7];
    ele[30][6] != ele[31][8];
    ele[30][6] != ele[31][9];
    ele[30][6] != ele[32][10];
    ele[30][6] != ele[32][11];
    ele[30][6] != ele[32][6];
    ele[30][6] != ele[32][7];
    ele[30][6] != ele[32][8];
    ele[30][6] != ele[32][9];
    ele[30][6] != ele[33][10];
    ele[30][6] != ele[33][11];
    ele[30][6] != ele[33][6];
    ele[30][6] != ele[33][7];
    ele[30][6] != ele[33][8];
    ele[30][6] != ele[33][9];
    ele[30][6] != ele[34][10];
    ele[30][6] != ele[34][11];
    ele[30][6] != ele[34][6];
    ele[30][6] != ele[34][7];
    ele[30][6] != ele[34][8];
    ele[30][6] != ele[34][9];
    ele[30][6] != ele[35][10];
    ele[30][6] != ele[35][11];
    ele[30][6] != ele[35][6];
    ele[30][6] != ele[35][7];
    ele[30][6] != ele[35][8];
    ele[30][6] != ele[35][9];
    ele[30][7] != ele[30][10];
    ele[30][7] != ele[30][11];
    ele[30][7] != ele[30][12];
    ele[30][7] != ele[30][13];
    ele[30][7] != ele[30][14];
    ele[30][7] != ele[30][15];
    ele[30][7] != ele[30][16];
    ele[30][7] != ele[30][17];
    ele[30][7] != ele[30][18];
    ele[30][7] != ele[30][19];
    ele[30][7] != ele[30][20];
    ele[30][7] != ele[30][21];
    ele[30][7] != ele[30][22];
    ele[30][7] != ele[30][23];
    ele[30][7] != ele[30][24];
    ele[30][7] != ele[30][25];
    ele[30][7] != ele[30][26];
    ele[30][7] != ele[30][27];
    ele[30][7] != ele[30][28];
    ele[30][7] != ele[30][29];
    ele[30][7] != ele[30][30];
    ele[30][7] != ele[30][31];
    ele[30][7] != ele[30][32];
    ele[30][7] != ele[30][33];
    ele[30][7] != ele[30][34];
    ele[30][7] != ele[30][35];
    ele[30][7] != ele[30][8];
    ele[30][7] != ele[30][9];
    ele[30][7] != ele[31][10];
    ele[30][7] != ele[31][11];
    ele[30][7] != ele[31][6];
    ele[30][7] != ele[31][7];
    ele[30][7] != ele[31][8];
    ele[30][7] != ele[31][9];
    ele[30][7] != ele[32][10];
    ele[30][7] != ele[32][11];
    ele[30][7] != ele[32][6];
    ele[30][7] != ele[32][7];
    ele[30][7] != ele[32][8];
    ele[30][7] != ele[32][9];
    ele[30][7] != ele[33][10];
    ele[30][7] != ele[33][11];
    ele[30][7] != ele[33][6];
    ele[30][7] != ele[33][7];
    ele[30][7] != ele[33][8];
    ele[30][7] != ele[33][9];
    ele[30][7] != ele[34][10];
    ele[30][7] != ele[34][11];
    ele[30][7] != ele[34][6];
    ele[30][7] != ele[34][7];
    ele[30][7] != ele[34][8];
    ele[30][7] != ele[34][9];
    ele[30][7] != ele[35][10];
    ele[30][7] != ele[35][11];
    ele[30][7] != ele[35][6];
    ele[30][7] != ele[35][7];
    ele[30][7] != ele[35][8];
    ele[30][7] != ele[35][9];
    ele[30][8] != ele[30][10];
    ele[30][8] != ele[30][11];
    ele[30][8] != ele[30][12];
    ele[30][8] != ele[30][13];
    ele[30][8] != ele[30][14];
    ele[30][8] != ele[30][15];
    ele[30][8] != ele[30][16];
    ele[30][8] != ele[30][17];
    ele[30][8] != ele[30][18];
    ele[30][8] != ele[30][19];
    ele[30][8] != ele[30][20];
    ele[30][8] != ele[30][21];
    ele[30][8] != ele[30][22];
    ele[30][8] != ele[30][23];
    ele[30][8] != ele[30][24];
    ele[30][8] != ele[30][25];
    ele[30][8] != ele[30][26];
    ele[30][8] != ele[30][27];
    ele[30][8] != ele[30][28];
    ele[30][8] != ele[30][29];
    ele[30][8] != ele[30][30];
    ele[30][8] != ele[30][31];
    ele[30][8] != ele[30][32];
    ele[30][8] != ele[30][33];
    ele[30][8] != ele[30][34];
    ele[30][8] != ele[30][35];
    ele[30][8] != ele[30][9];
    ele[30][8] != ele[31][10];
    ele[30][8] != ele[31][11];
    ele[30][8] != ele[31][6];
    ele[30][8] != ele[31][7];
    ele[30][8] != ele[31][8];
    ele[30][8] != ele[31][9];
    ele[30][8] != ele[32][10];
    ele[30][8] != ele[32][11];
    ele[30][8] != ele[32][6];
    ele[30][8] != ele[32][7];
    ele[30][8] != ele[32][8];
    ele[30][8] != ele[32][9];
    ele[30][8] != ele[33][10];
    ele[30][8] != ele[33][11];
    ele[30][8] != ele[33][6];
    ele[30][8] != ele[33][7];
    ele[30][8] != ele[33][8];
    ele[30][8] != ele[33][9];
    ele[30][8] != ele[34][10];
    ele[30][8] != ele[34][11];
    ele[30][8] != ele[34][6];
    ele[30][8] != ele[34][7];
    ele[30][8] != ele[34][8];
    ele[30][8] != ele[34][9];
    ele[30][8] != ele[35][10];
    ele[30][8] != ele[35][11];
    ele[30][8] != ele[35][6];
    ele[30][8] != ele[35][7];
    ele[30][8] != ele[35][8];
    ele[30][8] != ele[35][9];
    ele[30][9] != ele[30][10];
    ele[30][9] != ele[30][11];
    ele[30][9] != ele[30][12];
    ele[30][9] != ele[30][13];
    ele[30][9] != ele[30][14];
    ele[30][9] != ele[30][15];
    ele[30][9] != ele[30][16];
    ele[30][9] != ele[30][17];
    ele[30][9] != ele[30][18];
    ele[30][9] != ele[30][19];
    ele[30][9] != ele[30][20];
    ele[30][9] != ele[30][21];
    ele[30][9] != ele[30][22];
    ele[30][9] != ele[30][23];
    ele[30][9] != ele[30][24];
    ele[30][9] != ele[30][25];
    ele[30][9] != ele[30][26];
    ele[30][9] != ele[30][27];
    ele[30][9] != ele[30][28];
    ele[30][9] != ele[30][29];
    ele[30][9] != ele[30][30];
    ele[30][9] != ele[30][31];
    ele[30][9] != ele[30][32];
    ele[30][9] != ele[30][33];
    ele[30][9] != ele[30][34];
    ele[30][9] != ele[30][35];
    ele[30][9] != ele[31][10];
    ele[30][9] != ele[31][11];
    ele[30][9] != ele[31][6];
    ele[30][9] != ele[31][7];
    ele[30][9] != ele[31][8];
    ele[30][9] != ele[31][9];
    ele[30][9] != ele[32][10];
    ele[30][9] != ele[32][11];
    ele[30][9] != ele[32][6];
    ele[30][9] != ele[32][7];
    ele[30][9] != ele[32][8];
    ele[30][9] != ele[32][9];
    ele[30][9] != ele[33][10];
    ele[30][9] != ele[33][11];
    ele[30][9] != ele[33][6];
    ele[30][9] != ele[33][7];
    ele[30][9] != ele[33][8];
    ele[30][9] != ele[33][9];
    ele[30][9] != ele[34][10];
    ele[30][9] != ele[34][11];
    ele[30][9] != ele[34][6];
    ele[30][9] != ele[34][7];
    ele[30][9] != ele[34][8];
    ele[30][9] != ele[34][9];
    ele[30][9] != ele[35][10];
    ele[30][9] != ele[35][11];
    ele[30][9] != ele[35][6];
    ele[30][9] != ele[35][7];
    ele[30][9] != ele[35][8];
    ele[30][9] != ele[35][9];
    ele[31][0] != ele[31][1];
    ele[31][0] != ele[31][10];
    ele[31][0] != ele[31][11];
    ele[31][0] != ele[31][12];
    ele[31][0] != ele[31][13];
    ele[31][0] != ele[31][14];
    ele[31][0] != ele[31][15];
    ele[31][0] != ele[31][16];
    ele[31][0] != ele[31][17];
    ele[31][0] != ele[31][18];
    ele[31][0] != ele[31][19];
    ele[31][0] != ele[31][2];
    ele[31][0] != ele[31][20];
    ele[31][0] != ele[31][21];
    ele[31][0] != ele[31][22];
    ele[31][0] != ele[31][23];
    ele[31][0] != ele[31][24];
    ele[31][0] != ele[31][25];
    ele[31][0] != ele[31][26];
    ele[31][0] != ele[31][27];
    ele[31][0] != ele[31][28];
    ele[31][0] != ele[31][29];
    ele[31][0] != ele[31][3];
    ele[31][0] != ele[31][30];
    ele[31][0] != ele[31][31];
    ele[31][0] != ele[31][32];
    ele[31][0] != ele[31][33];
    ele[31][0] != ele[31][34];
    ele[31][0] != ele[31][35];
    ele[31][0] != ele[31][4];
    ele[31][0] != ele[31][5];
    ele[31][0] != ele[31][6];
    ele[31][0] != ele[31][7];
    ele[31][0] != ele[31][8];
    ele[31][0] != ele[31][9];
    ele[31][0] != ele[32][0];
    ele[31][0] != ele[32][1];
    ele[31][0] != ele[32][2];
    ele[31][0] != ele[32][3];
    ele[31][0] != ele[32][4];
    ele[31][0] != ele[32][5];
    ele[31][0] != ele[33][0];
    ele[31][0] != ele[33][1];
    ele[31][0] != ele[33][2];
    ele[31][0] != ele[33][3];
    ele[31][0] != ele[33][4];
    ele[31][0] != ele[33][5];
    ele[31][0] != ele[34][0];
    ele[31][0] != ele[34][1];
    ele[31][0] != ele[34][2];
    ele[31][0] != ele[34][3];
    ele[31][0] != ele[34][4];
    ele[31][0] != ele[34][5];
    ele[31][0] != ele[35][0];
    ele[31][0] != ele[35][1];
    ele[31][0] != ele[35][2];
    ele[31][0] != ele[35][3];
    ele[31][0] != ele[35][4];
    ele[31][0] != ele[35][5];
    ele[31][1] != ele[31][10];
    ele[31][1] != ele[31][11];
    ele[31][1] != ele[31][12];
    ele[31][1] != ele[31][13];
    ele[31][1] != ele[31][14];
    ele[31][1] != ele[31][15];
    ele[31][1] != ele[31][16];
    ele[31][1] != ele[31][17];
    ele[31][1] != ele[31][18];
    ele[31][1] != ele[31][19];
    ele[31][1] != ele[31][2];
    ele[31][1] != ele[31][20];
    ele[31][1] != ele[31][21];
    ele[31][1] != ele[31][22];
    ele[31][1] != ele[31][23];
    ele[31][1] != ele[31][24];
    ele[31][1] != ele[31][25];
    ele[31][1] != ele[31][26];
    ele[31][1] != ele[31][27];
    ele[31][1] != ele[31][28];
    ele[31][1] != ele[31][29];
    ele[31][1] != ele[31][3];
    ele[31][1] != ele[31][30];
    ele[31][1] != ele[31][31];
    ele[31][1] != ele[31][32];
    ele[31][1] != ele[31][33];
    ele[31][1] != ele[31][34];
    ele[31][1] != ele[31][35];
    ele[31][1] != ele[31][4];
    ele[31][1] != ele[31][5];
    ele[31][1] != ele[31][6];
    ele[31][1] != ele[31][7];
    ele[31][1] != ele[31][8];
    ele[31][1] != ele[31][9];
    ele[31][1] != ele[32][0];
    ele[31][1] != ele[32][1];
    ele[31][1] != ele[32][2];
    ele[31][1] != ele[32][3];
    ele[31][1] != ele[32][4];
    ele[31][1] != ele[32][5];
    ele[31][1] != ele[33][0];
    ele[31][1] != ele[33][1];
    ele[31][1] != ele[33][2];
    ele[31][1] != ele[33][3];
    ele[31][1] != ele[33][4];
    ele[31][1] != ele[33][5];
    ele[31][1] != ele[34][0];
    ele[31][1] != ele[34][1];
    ele[31][1] != ele[34][2];
    ele[31][1] != ele[34][3];
    ele[31][1] != ele[34][4];
    ele[31][1] != ele[34][5];
    ele[31][1] != ele[35][0];
    ele[31][1] != ele[35][1];
    ele[31][1] != ele[35][2];
    ele[31][1] != ele[35][3];
    ele[31][1] != ele[35][4];
    ele[31][1] != ele[35][5];
    ele[31][10] != ele[31][11];
    ele[31][10] != ele[31][12];
    ele[31][10] != ele[31][13];
    ele[31][10] != ele[31][14];
    ele[31][10] != ele[31][15];
    ele[31][10] != ele[31][16];
    ele[31][10] != ele[31][17];
    ele[31][10] != ele[31][18];
    ele[31][10] != ele[31][19];
    ele[31][10] != ele[31][20];
    ele[31][10] != ele[31][21];
    ele[31][10] != ele[31][22];
    ele[31][10] != ele[31][23];
    ele[31][10] != ele[31][24];
    ele[31][10] != ele[31][25];
    ele[31][10] != ele[31][26];
    ele[31][10] != ele[31][27];
    ele[31][10] != ele[31][28];
    ele[31][10] != ele[31][29];
    ele[31][10] != ele[31][30];
    ele[31][10] != ele[31][31];
    ele[31][10] != ele[31][32];
    ele[31][10] != ele[31][33];
    ele[31][10] != ele[31][34];
    ele[31][10] != ele[31][35];
    ele[31][10] != ele[32][10];
    ele[31][10] != ele[32][11];
    ele[31][10] != ele[32][6];
    ele[31][10] != ele[32][7];
    ele[31][10] != ele[32][8];
    ele[31][10] != ele[32][9];
    ele[31][10] != ele[33][10];
    ele[31][10] != ele[33][11];
    ele[31][10] != ele[33][6];
    ele[31][10] != ele[33][7];
    ele[31][10] != ele[33][8];
    ele[31][10] != ele[33][9];
    ele[31][10] != ele[34][10];
    ele[31][10] != ele[34][11];
    ele[31][10] != ele[34][6];
    ele[31][10] != ele[34][7];
    ele[31][10] != ele[34][8];
    ele[31][10] != ele[34][9];
    ele[31][10] != ele[35][10];
    ele[31][10] != ele[35][11];
    ele[31][10] != ele[35][6];
    ele[31][10] != ele[35][7];
    ele[31][10] != ele[35][8];
    ele[31][10] != ele[35][9];
    ele[31][11] != ele[31][12];
    ele[31][11] != ele[31][13];
    ele[31][11] != ele[31][14];
    ele[31][11] != ele[31][15];
    ele[31][11] != ele[31][16];
    ele[31][11] != ele[31][17];
    ele[31][11] != ele[31][18];
    ele[31][11] != ele[31][19];
    ele[31][11] != ele[31][20];
    ele[31][11] != ele[31][21];
    ele[31][11] != ele[31][22];
    ele[31][11] != ele[31][23];
    ele[31][11] != ele[31][24];
    ele[31][11] != ele[31][25];
    ele[31][11] != ele[31][26];
    ele[31][11] != ele[31][27];
    ele[31][11] != ele[31][28];
    ele[31][11] != ele[31][29];
    ele[31][11] != ele[31][30];
    ele[31][11] != ele[31][31];
    ele[31][11] != ele[31][32];
    ele[31][11] != ele[31][33];
    ele[31][11] != ele[31][34];
    ele[31][11] != ele[31][35];
    ele[31][11] != ele[32][10];
    ele[31][11] != ele[32][11];
    ele[31][11] != ele[32][6];
    ele[31][11] != ele[32][7];
    ele[31][11] != ele[32][8];
    ele[31][11] != ele[32][9];
    ele[31][11] != ele[33][10];
    ele[31][11] != ele[33][11];
    ele[31][11] != ele[33][6];
    ele[31][11] != ele[33][7];
    ele[31][11] != ele[33][8];
    ele[31][11] != ele[33][9];
    ele[31][11] != ele[34][10];
    ele[31][11] != ele[34][11];
    ele[31][11] != ele[34][6];
    ele[31][11] != ele[34][7];
    ele[31][11] != ele[34][8];
    ele[31][11] != ele[34][9];
    ele[31][11] != ele[35][10];
    ele[31][11] != ele[35][11];
    ele[31][11] != ele[35][6];
    ele[31][11] != ele[35][7];
    ele[31][11] != ele[35][8];
    ele[31][11] != ele[35][9];
    ele[31][12] != ele[31][13];
    ele[31][12] != ele[31][14];
    ele[31][12] != ele[31][15];
    ele[31][12] != ele[31][16];
    ele[31][12] != ele[31][17];
    ele[31][12] != ele[31][18];
    ele[31][12] != ele[31][19];
    ele[31][12] != ele[31][20];
    ele[31][12] != ele[31][21];
    ele[31][12] != ele[31][22];
    ele[31][12] != ele[31][23];
    ele[31][12] != ele[31][24];
    ele[31][12] != ele[31][25];
    ele[31][12] != ele[31][26];
    ele[31][12] != ele[31][27];
    ele[31][12] != ele[31][28];
    ele[31][12] != ele[31][29];
    ele[31][12] != ele[31][30];
    ele[31][12] != ele[31][31];
    ele[31][12] != ele[31][32];
    ele[31][12] != ele[31][33];
    ele[31][12] != ele[31][34];
    ele[31][12] != ele[31][35];
    ele[31][12] != ele[32][12];
    ele[31][12] != ele[32][13];
    ele[31][12] != ele[32][14];
    ele[31][12] != ele[32][15];
    ele[31][12] != ele[32][16];
    ele[31][12] != ele[32][17];
    ele[31][12] != ele[33][12];
    ele[31][12] != ele[33][13];
    ele[31][12] != ele[33][14];
    ele[31][12] != ele[33][15];
    ele[31][12] != ele[33][16];
    ele[31][12] != ele[33][17];
    ele[31][12] != ele[34][12];
    ele[31][12] != ele[34][13];
    ele[31][12] != ele[34][14];
    ele[31][12] != ele[34][15];
    ele[31][12] != ele[34][16];
    ele[31][12] != ele[34][17];
    ele[31][12] != ele[35][12];
    ele[31][12] != ele[35][13];
    ele[31][12] != ele[35][14];
    ele[31][12] != ele[35][15];
    ele[31][12] != ele[35][16];
    ele[31][12] != ele[35][17];
    ele[31][13] != ele[31][14];
    ele[31][13] != ele[31][15];
    ele[31][13] != ele[31][16];
    ele[31][13] != ele[31][17];
    ele[31][13] != ele[31][18];
    ele[31][13] != ele[31][19];
    ele[31][13] != ele[31][20];
    ele[31][13] != ele[31][21];
    ele[31][13] != ele[31][22];
    ele[31][13] != ele[31][23];
    ele[31][13] != ele[31][24];
    ele[31][13] != ele[31][25];
    ele[31][13] != ele[31][26];
    ele[31][13] != ele[31][27];
    ele[31][13] != ele[31][28];
    ele[31][13] != ele[31][29];
    ele[31][13] != ele[31][30];
    ele[31][13] != ele[31][31];
    ele[31][13] != ele[31][32];
    ele[31][13] != ele[31][33];
    ele[31][13] != ele[31][34];
    ele[31][13] != ele[31][35];
    ele[31][13] != ele[32][12];
    ele[31][13] != ele[32][13];
    ele[31][13] != ele[32][14];
    ele[31][13] != ele[32][15];
    ele[31][13] != ele[32][16];
    ele[31][13] != ele[32][17];
    ele[31][13] != ele[33][12];
    ele[31][13] != ele[33][13];
    ele[31][13] != ele[33][14];
    ele[31][13] != ele[33][15];
    ele[31][13] != ele[33][16];
    ele[31][13] != ele[33][17];
    ele[31][13] != ele[34][12];
    ele[31][13] != ele[34][13];
    ele[31][13] != ele[34][14];
    ele[31][13] != ele[34][15];
    ele[31][13] != ele[34][16];
    ele[31][13] != ele[34][17];
    ele[31][13] != ele[35][12];
    ele[31][13] != ele[35][13];
    ele[31][13] != ele[35][14];
    ele[31][13] != ele[35][15];
    ele[31][13] != ele[35][16];
    ele[31][13] != ele[35][17];
    ele[31][14] != ele[31][15];
    ele[31][14] != ele[31][16];
    ele[31][14] != ele[31][17];
    ele[31][14] != ele[31][18];
    ele[31][14] != ele[31][19];
    ele[31][14] != ele[31][20];
    ele[31][14] != ele[31][21];
    ele[31][14] != ele[31][22];
    ele[31][14] != ele[31][23];
    ele[31][14] != ele[31][24];
    ele[31][14] != ele[31][25];
    ele[31][14] != ele[31][26];
    ele[31][14] != ele[31][27];
    ele[31][14] != ele[31][28];
    ele[31][14] != ele[31][29];
    ele[31][14] != ele[31][30];
    ele[31][14] != ele[31][31];
    ele[31][14] != ele[31][32];
    ele[31][14] != ele[31][33];
    ele[31][14] != ele[31][34];
    ele[31][14] != ele[31][35];
    ele[31][14] != ele[32][12];
    ele[31][14] != ele[32][13];
    ele[31][14] != ele[32][14];
    ele[31][14] != ele[32][15];
    ele[31][14] != ele[32][16];
    ele[31][14] != ele[32][17];
    ele[31][14] != ele[33][12];
    ele[31][14] != ele[33][13];
    ele[31][14] != ele[33][14];
    ele[31][14] != ele[33][15];
    ele[31][14] != ele[33][16];
    ele[31][14] != ele[33][17];
    ele[31][14] != ele[34][12];
    ele[31][14] != ele[34][13];
    ele[31][14] != ele[34][14];
    ele[31][14] != ele[34][15];
    ele[31][14] != ele[34][16];
    ele[31][14] != ele[34][17];
    ele[31][14] != ele[35][12];
    ele[31][14] != ele[35][13];
    ele[31][14] != ele[35][14];
    ele[31][14] != ele[35][15];
    ele[31][14] != ele[35][16];
    ele[31][14] != ele[35][17];
    ele[31][15] != ele[31][16];
    ele[31][15] != ele[31][17];
    ele[31][15] != ele[31][18];
    ele[31][15] != ele[31][19];
    ele[31][15] != ele[31][20];
    ele[31][15] != ele[31][21];
    ele[31][15] != ele[31][22];
    ele[31][15] != ele[31][23];
    ele[31][15] != ele[31][24];
    ele[31][15] != ele[31][25];
    ele[31][15] != ele[31][26];
    ele[31][15] != ele[31][27];
    ele[31][15] != ele[31][28];
    ele[31][15] != ele[31][29];
    ele[31][15] != ele[31][30];
    ele[31][15] != ele[31][31];
    ele[31][15] != ele[31][32];
    ele[31][15] != ele[31][33];
    ele[31][15] != ele[31][34];
    ele[31][15] != ele[31][35];
    ele[31][15] != ele[32][12];
    ele[31][15] != ele[32][13];
    ele[31][15] != ele[32][14];
    ele[31][15] != ele[32][15];
    ele[31][15] != ele[32][16];
    ele[31][15] != ele[32][17];
    ele[31][15] != ele[33][12];
    ele[31][15] != ele[33][13];
    ele[31][15] != ele[33][14];
    ele[31][15] != ele[33][15];
    ele[31][15] != ele[33][16];
    ele[31][15] != ele[33][17];
    ele[31][15] != ele[34][12];
    ele[31][15] != ele[34][13];
    ele[31][15] != ele[34][14];
    ele[31][15] != ele[34][15];
    ele[31][15] != ele[34][16];
    ele[31][15] != ele[34][17];
    ele[31][15] != ele[35][12];
    ele[31][15] != ele[35][13];
    ele[31][15] != ele[35][14];
    ele[31][15] != ele[35][15];
    ele[31][15] != ele[35][16];
    ele[31][15] != ele[35][17];
    ele[31][16] != ele[31][17];
    ele[31][16] != ele[31][18];
    ele[31][16] != ele[31][19];
    ele[31][16] != ele[31][20];
    ele[31][16] != ele[31][21];
    ele[31][16] != ele[31][22];
    ele[31][16] != ele[31][23];
    ele[31][16] != ele[31][24];
    ele[31][16] != ele[31][25];
    ele[31][16] != ele[31][26];
    ele[31][16] != ele[31][27];
    ele[31][16] != ele[31][28];
    ele[31][16] != ele[31][29];
    ele[31][16] != ele[31][30];
    ele[31][16] != ele[31][31];
    ele[31][16] != ele[31][32];
    ele[31][16] != ele[31][33];
    ele[31][16] != ele[31][34];
    ele[31][16] != ele[31][35];
    ele[31][16] != ele[32][12];
    ele[31][16] != ele[32][13];
    ele[31][16] != ele[32][14];
    ele[31][16] != ele[32][15];
    ele[31][16] != ele[32][16];
    ele[31][16] != ele[32][17];
    ele[31][16] != ele[33][12];
    ele[31][16] != ele[33][13];
    ele[31][16] != ele[33][14];
    ele[31][16] != ele[33][15];
    ele[31][16] != ele[33][16];
    ele[31][16] != ele[33][17];
    ele[31][16] != ele[34][12];
    ele[31][16] != ele[34][13];
    ele[31][16] != ele[34][14];
    ele[31][16] != ele[34][15];
    ele[31][16] != ele[34][16];
    ele[31][16] != ele[34][17];
    ele[31][16] != ele[35][12];
    ele[31][16] != ele[35][13];
    ele[31][16] != ele[35][14];
    ele[31][16] != ele[35][15];
    ele[31][16] != ele[35][16];
    ele[31][16] != ele[35][17];
    ele[31][17] != ele[31][18];
    ele[31][17] != ele[31][19];
    ele[31][17] != ele[31][20];
    ele[31][17] != ele[31][21];
    ele[31][17] != ele[31][22];
    ele[31][17] != ele[31][23];
    ele[31][17] != ele[31][24];
    ele[31][17] != ele[31][25];
    ele[31][17] != ele[31][26];
    ele[31][17] != ele[31][27];
    ele[31][17] != ele[31][28];
    ele[31][17] != ele[31][29];
    ele[31][17] != ele[31][30];
    ele[31][17] != ele[31][31];
    ele[31][17] != ele[31][32];
    ele[31][17] != ele[31][33];
    ele[31][17] != ele[31][34];
    ele[31][17] != ele[31][35];
    ele[31][17] != ele[32][12];
    ele[31][17] != ele[32][13];
    ele[31][17] != ele[32][14];
    ele[31][17] != ele[32][15];
    ele[31][17] != ele[32][16];
    ele[31][17] != ele[32][17];
    ele[31][17] != ele[33][12];
    ele[31][17] != ele[33][13];
    ele[31][17] != ele[33][14];
    ele[31][17] != ele[33][15];
    ele[31][17] != ele[33][16];
    ele[31][17] != ele[33][17];
    ele[31][17] != ele[34][12];
    ele[31][17] != ele[34][13];
    ele[31][17] != ele[34][14];
    ele[31][17] != ele[34][15];
    ele[31][17] != ele[34][16];
    ele[31][17] != ele[34][17];
    ele[31][17] != ele[35][12];
    ele[31][17] != ele[35][13];
    ele[31][17] != ele[35][14];
    ele[31][17] != ele[35][15];
    ele[31][17] != ele[35][16];
    ele[31][17] != ele[35][17];
    ele[31][18] != ele[31][19];
    ele[31][18] != ele[31][20];
    ele[31][18] != ele[31][21];
    ele[31][18] != ele[31][22];
    ele[31][18] != ele[31][23];
    ele[31][18] != ele[31][24];
    ele[31][18] != ele[31][25];
    ele[31][18] != ele[31][26];
    ele[31][18] != ele[31][27];
    ele[31][18] != ele[31][28];
    ele[31][18] != ele[31][29];
    ele[31][18] != ele[31][30];
    ele[31][18] != ele[31][31];
    ele[31][18] != ele[31][32];
    ele[31][18] != ele[31][33];
    ele[31][18] != ele[31][34];
    ele[31][18] != ele[31][35];
    ele[31][18] != ele[32][18];
    ele[31][18] != ele[32][19];
    ele[31][18] != ele[32][20];
    ele[31][18] != ele[32][21];
    ele[31][18] != ele[32][22];
    ele[31][18] != ele[32][23];
    ele[31][18] != ele[33][18];
    ele[31][18] != ele[33][19];
    ele[31][18] != ele[33][20];
    ele[31][18] != ele[33][21];
    ele[31][18] != ele[33][22];
    ele[31][18] != ele[33][23];
    ele[31][18] != ele[34][18];
    ele[31][18] != ele[34][19];
    ele[31][18] != ele[34][20];
    ele[31][18] != ele[34][21];
    ele[31][18] != ele[34][22];
    ele[31][18] != ele[34][23];
    ele[31][18] != ele[35][18];
    ele[31][18] != ele[35][19];
    ele[31][18] != ele[35][20];
    ele[31][18] != ele[35][21];
    ele[31][18] != ele[35][22];
    ele[31][18] != ele[35][23];
    ele[31][19] != ele[31][20];
    ele[31][19] != ele[31][21];
    ele[31][19] != ele[31][22];
    ele[31][19] != ele[31][23];
    ele[31][19] != ele[31][24];
    ele[31][19] != ele[31][25];
    ele[31][19] != ele[31][26];
    ele[31][19] != ele[31][27];
    ele[31][19] != ele[31][28];
    ele[31][19] != ele[31][29];
    ele[31][19] != ele[31][30];
    ele[31][19] != ele[31][31];
    ele[31][19] != ele[31][32];
    ele[31][19] != ele[31][33];
    ele[31][19] != ele[31][34];
    ele[31][19] != ele[31][35];
    ele[31][19] != ele[32][18];
    ele[31][19] != ele[32][19];
    ele[31][19] != ele[32][20];
    ele[31][19] != ele[32][21];
    ele[31][19] != ele[32][22];
    ele[31][19] != ele[32][23];
    ele[31][19] != ele[33][18];
    ele[31][19] != ele[33][19];
    ele[31][19] != ele[33][20];
    ele[31][19] != ele[33][21];
    ele[31][19] != ele[33][22];
    ele[31][19] != ele[33][23];
    ele[31][19] != ele[34][18];
    ele[31][19] != ele[34][19];
    ele[31][19] != ele[34][20];
    ele[31][19] != ele[34][21];
    ele[31][19] != ele[34][22];
    ele[31][19] != ele[34][23];
    ele[31][19] != ele[35][18];
    ele[31][19] != ele[35][19];
    ele[31][19] != ele[35][20];
    ele[31][19] != ele[35][21];
    ele[31][19] != ele[35][22];
    ele[31][19] != ele[35][23];
    ele[31][2] != ele[31][10];
    ele[31][2] != ele[31][11];
    ele[31][2] != ele[31][12];
    ele[31][2] != ele[31][13];
    ele[31][2] != ele[31][14];
    ele[31][2] != ele[31][15];
    ele[31][2] != ele[31][16];
    ele[31][2] != ele[31][17];
    ele[31][2] != ele[31][18];
    ele[31][2] != ele[31][19];
    ele[31][2] != ele[31][20];
    ele[31][2] != ele[31][21];
    ele[31][2] != ele[31][22];
    ele[31][2] != ele[31][23];
    ele[31][2] != ele[31][24];
    ele[31][2] != ele[31][25];
    ele[31][2] != ele[31][26];
    ele[31][2] != ele[31][27];
    ele[31][2] != ele[31][28];
    ele[31][2] != ele[31][29];
    ele[31][2] != ele[31][3];
    ele[31][2] != ele[31][30];
    ele[31][2] != ele[31][31];
    ele[31][2] != ele[31][32];
    ele[31][2] != ele[31][33];
    ele[31][2] != ele[31][34];
    ele[31][2] != ele[31][35];
    ele[31][2] != ele[31][4];
    ele[31][2] != ele[31][5];
    ele[31][2] != ele[31][6];
    ele[31][2] != ele[31][7];
    ele[31][2] != ele[31][8];
    ele[31][2] != ele[31][9];
    ele[31][2] != ele[32][0];
    ele[31][2] != ele[32][1];
    ele[31][2] != ele[32][2];
    ele[31][2] != ele[32][3];
    ele[31][2] != ele[32][4];
    ele[31][2] != ele[32][5];
    ele[31][2] != ele[33][0];
    ele[31][2] != ele[33][1];
    ele[31][2] != ele[33][2];
    ele[31][2] != ele[33][3];
    ele[31][2] != ele[33][4];
    ele[31][2] != ele[33][5];
    ele[31][2] != ele[34][0];
    ele[31][2] != ele[34][1];
    ele[31][2] != ele[34][2];
    ele[31][2] != ele[34][3];
    ele[31][2] != ele[34][4];
    ele[31][2] != ele[34][5];
    ele[31][2] != ele[35][0];
    ele[31][2] != ele[35][1];
    ele[31][2] != ele[35][2];
    ele[31][2] != ele[35][3];
    ele[31][2] != ele[35][4];
    ele[31][2] != ele[35][5];
    ele[31][20] != ele[31][21];
    ele[31][20] != ele[31][22];
    ele[31][20] != ele[31][23];
    ele[31][20] != ele[31][24];
    ele[31][20] != ele[31][25];
    ele[31][20] != ele[31][26];
    ele[31][20] != ele[31][27];
    ele[31][20] != ele[31][28];
    ele[31][20] != ele[31][29];
    ele[31][20] != ele[31][30];
    ele[31][20] != ele[31][31];
    ele[31][20] != ele[31][32];
    ele[31][20] != ele[31][33];
    ele[31][20] != ele[31][34];
    ele[31][20] != ele[31][35];
    ele[31][20] != ele[32][18];
    ele[31][20] != ele[32][19];
    ele[31][20] != ele[32][20];
    ele[31][20] != ele[32][21];
    ele[31][20] != ele[32][22];
    ele[31][20] != ele[32][23];
    ele[31][20] != ele[33][18];
    ele[31][20] != ele[33][19];
    ele[31][20] != ele[33][20];
    ele[31][20] != ele[33][21];
    ele[31][20] != ele[33][22];
    ele[31][20] != ele[33][23];
    ele[31][20] != ele[34][18];
    ele[31][20] != ele[34][19];
    ele[31][20] != ele[34][20];
    ele[31][20] != ele[34][21];
    ele[31][20] != ele[34][22];
    ele[31][20] != ele[34][23];
    ele[31][20] != ele[35][18];
    ele[31][20] != ele[35][19];
    ele[31][20] != ele[35][20];
    ele[31][20] != ele[35][21];
    ele[31][20] != ele[35][22];
    ele[31][20] != ele[35][23];
    ele[31][21] != ele[31][22];
    ele[31][21] != ele[31][23];
    ele[31][21] != ele[31][24];
    ele[31][21] != ele[31][25];
    ele[31][21] != ele[31][26];
    ele[31][21] != ele[31][27];
    ele[31][21] != ele[31][28];
    ele[31][21] != ele[31][29];
    ele[31][21] != ele[31][30];
    ele[31][21] != ele[31][31];
    ele[31][21] != ele[31][32];
    ele[31][21] != ele[31][33];
    ele[31][21] != ele[31][34];
    ele[31][21] != ele[31][35];
    ele[31][21] != ele[32][18];
    ele[31][21] != ele[32][19];
    ele[31][21] != ele[32][20];
    ele[31][21] != ele[32][21];
    ele[31][21] != ele[32][22];
    ele[31][21] != ele[32][23];
    ele[31][21] != ele[33][18];
    ele[31][21] != ele[33][19];
    ele[31][21] != ele[33][20];
    ele[31][21] != ele[33][21];
    ele[31][21] != ele[33][22];
    ele[31][21] != ele[33][23];
    ele[31][21] != ele[34][18];
    ele[31][21] != ele[34][19];
    ele[31][21] != ele[34][20];
    ele[31][21] != ele[34][21];
    ele[31][21] != ele[34][22];
    ele[31][21] != ele[34][23];
    ele[31][21] != ele[35][18];
    ele[31][21] != ele[35][19];
    ele[31][21] != ele[35][20];
    ele[31][21] != ele[35][21];
    ele[31][21] != ele[35][22];
    ele[31][21] != ele[35][23];
    ele[31][22] != ele[31][23];
    ele[31][22] != ele[31][24];
    ele[31][22] != ele[31][25];
    ele[31][22] != ele[31][26];
    ele[31][22] != ele[31][27];
    ele[31][22] != ele[31][28];
    ele[31][22] != ele[31][29];
    ele[31][22] != ele[31][30];
    ele[31][22] != ele[31][31];
    ele[31][22] != ele[31][32];
    ele[31][22] != ele[31][33];
    ele[31][22] != ele[31][34];
    ele[31][22] != ele[31][35];
    ele[31][22] != ele[32][18];
    ele[31][22] != ele[32][19];
    ele[31][22] != ele[32][20];
    ele[31][22] != ele[32][21];
    ele[31][22] != ele[32][22];
    ele[31][22] != ele[32][23];
    ele[31][22] != ele[33][18];
    ele[31][22] != ele[33][19];
    ele[31][22] != ele[33][20];
    ele[31][22] != ele[33][21];
    ele[31][22] != ele[33][22];
    ele[31][22] != ele[33][23];
    ele[31][22] != ele[34][18];
    ele[31][22] != ele[34][19];
    ele[31][22] != ele[34][20];
    ele[31][22] != ele[34][21];
    ele[31][22] != ele[34][22];
    ele[31][22] != ele[34][23];
    ele[31][22] != ele[35][18];
    ele[31][22] != ele[35][19];
    ele[31][22] != ele[35][20];
    ele[31][22] != ele[35][21];
    ele[31][22] != ele[35][22];
    ele[31][22] != ele[35][23];
    ele[31][23] != ele[31][24];
    ele[31][23] != ele[31][25];
    ele[31][23] != ele[31][26];
    ele[31][23] != ele[31][27];
    ele[31][23] != ele[31][28];
    ele[31][23] != ele[31][29];
    ele[31][23] != ele[31][30];
    ele[31][23] != ele[31][31];
    ele[31][23] != ele[31][32];
    ele[31][23] != ele[31][33];
    ele[31][23] != ele[31][34];
    ele[31][23] != ele[31][35];
    ele[31][23] != ele[32][18];
    ele[31][23] != ele[32][19];
    ele[31][23] != ele[32][20];
    ele[31][23] != ele[32][21];
    ele[31][23] != ele[32][22];
    ele[31][23] != ele[32][23];
    ele[31][23] != ele[33][18];
    ele[31][23] != ele[33][19];
    ele[31][23] != ele[33][20];
    ele[31][23] != ele[33][21];
    ele[31][23] != ele[33][22];
    ele[31][23] != ele[33][23];
    ele[31][23] != ele[34][18];
    ele[31][23] != ele[34][19];
    ele[31][23] != ele[34][20];
    ele[31][23] != ele[34][21];
    ele[31][23] != ele[34][22];
    ele[31][23] != ele[34][23];
    ele[31][23] != ele[35][18];
    ele[31][23] != ele[35][19];
    ele[31][23] != ele[35][20];
    ele[31][23] != ele[35][21];
    ele[31][23] != ele[35][22];
    ele[31][23] != ele[35][23];
    ele[31][24] != ele[31][25];
    ele[31][24] != ele[31][26];
    ele[31][24] != ele[31][27];
    ele[31][24] != ele[31][28];
    ele[31][24] != ele[31][29];
    ele[31][24] != ele[31][30];
    ele[31][24] != ele[31][31];
    ele[31][24] != ele[31][32];
    ele[31][24] != ele[31][33];
    ele[31][24] != ele[31][34];
    ele[31][24] != ele[31][35];
    ele[31][24] != ele[32][24];
    ele[31][24] != ele[32][25];
    ele[31][24] != ele[32][26];
    ele[31][24] != ele[32][27];
    ele[31][24] != ele[32][28];
    ele[31][24] != ele[32][29];
    ele[31][24] != ele[33][24];
    ele[31][24] != ele[33][25];
    ele[31][24] != ele[33][26];
    ele[31][24] != ele[33][27];
    ele[31][24] != ele[33][28];
    ele[31][24] != ele[33][29];
    ele[31][24] != ele[34][24];
    ele[31][24] != ele[34][25];
    ele[31][24] != ele[34][26];
    ele[31][24] != ele[34][27];
    ele[31][24] != ele[34][28];
    ele[31][24] != ele[34][29];
    ele[31][24] != ele[35][24];
    ele[31][24] != ele[35][25];
    ele[31][24] != ele[35][26];
    ele[31][24] != ele[35][27];
    ele[31][24] != ele[35][28];
    ele[31][24] != ele[35][29];
    ele[31][25] != ele[31][26];
    ele[31][25] != ele[31][27];
    ele[31][25] != ele[31][28];
    ele[31][25] != ele[31][29];
    ele[31][25] != ele[31][30];
    ele[31][25] != ele[31][31];
    ele[31][25] != ele[31][32];
    ele[31][25] != ele[31][33];
    ele[31][25] != ele[31][34];
    ele[31][25] != ele[31][35];
    ele[31][25] != ele[32][24];
    ele[31][25] != ele[32][25];
    ele[31][25] != ele[32][26];
    ele[31][25] != ele[32][27];
    ele[31][25] != ele[32][28];
    ele[31][25] != ele[32][29];
    ele[31][25] != ele[33][24];
    ele[31][25] != ele[33][25];
    ele[31][25] != ele[33][26];
    ele[31][25] != ele[33][27];
    ele[31][25] != ele[33][28];
    ele[31][25] != ele[33][29];
    ele[31][25] != ele[34][24];
    ele[31][25] != ele[34][25];
    ele[31][25] != ele[34][26];
    ele[31][25] != ele[34][27];
    ele[31][25] != ele[34][28];
    ele[31][25] != ele[34][29];
    ele[31][25] != ele[35][24];
    ele[31][25] != ele[35][25];
    ele[31][25] != ele[35][26];
    ele[31][25] != ele[35][27];
    ele[31][25] != ele[35][28];
    ele[31][25] != ele[35][29];
    ele[31][26] != ele[31][27];
    ele[31][26] != ele[31][28];
    ele[31][26] != ele[31][29];
    ele[31][26] != ele[31][30];
    ele[31][26] != ele[31][31];
    ele[31][26] != ele[31][32];
    ele[31][26] != ele[31][33];
    ele[31][26] != ele[31][34];
    ele[31][26] != ele[31][35];
    ele[31][26] != ele[32][24];
    ele[31][26] != ele[32][25];
    ele[31][26] != ele[32][26];
    ele[31][26] != ele[32][27];
    ele[31][26] != ele[32][28];
    ele[31][26] != ele[32][29];
    ele[31][26] != ele[33][24];
    ele[31][26] != ele[33][25];
    ele[31][26] != ele[33][26];
    ele[31][26] != ele[33][27];
    ele[31][26] != ele[33][28];
    ele[31][26] != ele[33][29];
    ele[31][26] != ele[34][24];
    ele[31][26] != ele[34][25];
    ele[31][26] != ele[34][26];
    ele[31][26] != ele[34][27];
    ele[31][26] != ele[34][28];
    ele[31][26] != ele[34][29];
    ele[31][26] != ele[35][24];
    ele[31][26] != ele[35][25];
    ele[31][26] != ele[35][26];
    ele[31][26] != ele[35][27];
    ele[31][26] != ele[35][28];
    ele[31][26] != ele[35][29];
    ele[31][27] != ele[31][28];
    ele[31][27] != ele[31][29];
    ele[31][27] != ele[31][30];
    ele[31][27] != ele[31][31];
    ele[31][27] != ele[31][32];
    ele[31][27] != ele[31][33];
    ele[31][27] != ele[31][34];
    ele[31][27] != ele[31][35];
    ele[31][27] != ele[32][24];
    ele[31][27] != ele[32][25];
    ele[31][27] != ele[32][26];
    ele[31][27] != ele[32][27];
    ele[31][27] != ele[32][28];
    ele[31][27] != ele[32][29];
    ele[31][27] != ele[33][24];
    ele[31][27] != ele[33][25];
    ele[31][27] != ele[33][26];
    ele[31][27] != ele[33][27];
    ele[31][27] != ele[33][28];
    ele[31][27] != ele[33][29];
    ele[31][27] != ele[34][24];
    ele[31][27] != ele[34][25];
    ele[31][27] != ele[34][26];
    ele[31][27] != ele[34][27];
    ele[31][27] != ele[34][28];
    ele[31][27] != ele[34][29];
    ele[31][27] != ele[35][24];
    ele[31][27] != ele[35][25];
    ele[31][27] != ele[35][26];
    ele[31][27] != ele[35][27];
    ele[31][27] != ele[35][28];
    ele[31][27] != ele[35][29];
    ele[31][28] != ele[31][29];
    ele[31][28] != ele[31][30];
    ele[31][28] != ele[31][31];
    ele[31][28] != ele[31][32];
    ele[31][28] != ele[31][33];
    ele[31][28] != ele[31][34];
    ele[31][28] != ele[31][35];
    ele[31][28] != ele[32][24];
    ele[31][28] != ele[32][25];
    ele[31][28] != ele[32][26];
    ele[31][28] != ele[32][27];
    ele[31][28] != ele[32][28];
    ele[31][28] != ele[32][29];
    ele[31][28] != ele[33][24];
    ele[31][28] != ele[33][25];
    ele[31][28] != ele[33][26];
    ele[31][28] != ele[33][27];
    ele[31][28] != ele[33][28];
    ele[31][28] != ele[33][29];
    ele[31][28] != ele[34][24];
    ele[31][28] != ele[34][25];
    ele[31][28] != ele[34][26];
    ele[31][28] != ele[34][27];
    ele[31][28] != ele[34][28];
    ele[31][28] != ele[34][29];
    ele[31][28] != ele[35][24];
    ele[31][28] != ele[35][25];
    ele[31][28] != ele[35][26];
    ele[31][28] != ele[35][27];
    ele[31][28] != ele[35][28];
    ele[31][28] != ele[35][29];
    ele[31][29] != ele[31][30];
    ele[31][29] != ele[31][31];
    ele[31][29] != ele[31][32];
    ele[31][29] != ele[31][33];
    ele[31][29] != ele[31][34];
    ele[31][29] != ele[31][35];
    ele[31][29] != ele[32][24];
    ele[31][29] != ele[32][25];
    ele[31][29] != ele[32][26];
    ele[31][29] != ele[32][27];
    ele[31][29] != ele[32][28];
    ele[31][29] != ele[32][29];
    ele[31][29] != ele[33][24];
    ele[31][29] != ele[33][25];
    ele[31][29] != ele[33][26];
    ele[31][29] != ele[33][27];
    ele[31][29] != ele[33][28];
    ele[31][29] != ele[33][29];
    ele[31][29] != ele[34][24];
    ele[31][29] != ele[34][25];
    ele[31][29] != ele[34][26];
    ele[31][29] != ele[34][27];
    ele[31][29] != ele[34][28];
    ele[31][29] != ele[34][29];
    ele[31][29] != ele[35][24];
    ele[31][29] != ele[35][25];
    ele[31][29] != ele[35][26];
    ele[31][29] != ele[35][27];
    ele[31][29] != ele[35][28];
    ele[31][29] != ele[35][29];
    ele[31][3] != ele[31][10];
    ele[31][3] != ele[31][11];
    ele[31][3] != ele[31][12];
    ele[31][3] != ele[31][13];
    ele[31][3] != ele[31][14];
    ele[31][3] != ele[31][15];
    ele[31][3] != ele[31][16];
    ele[31][3] != ele[31][17];
    ele[31][3] != ele[31][18];
    ele[31][3] != ele[31][19];
    ele[31][3] != ele[31][20];
    ele[31][3] != ele[31][21];
    ele[31][3] != ele[31][22];
    ele[31][3] != ele[31][23];
    ele[31][3] != ele[31][24];
    ele[31][3] != ele[31][25];
    ele[31][3] != ele[31][26];
    ele[31][3] != ele[31][27];
    ele[31][3] != ele[31][28];
    ele[31][3] != ele[31][29];
    ele[31][3] != ele[31][30];
    ele[31][3] != ele[31][31];
    ele[31][3] != ele[31][32];
    ele[31][3] != ele[31][33];
    ele[31][3] != ele[31][34];
    ele[31][3] != ele[31][35];
    ele[31][3] != ele[31][4];
    ele[31][3] != ele[31][5];
    ele[31][3] != ele[31][6];
    ele[31][3] != ele[31][7];
    ele[31][3] != ele[31][8];
    ele[31][3] != ele[31][9];
    ele[31][3] != ele[32][0];
    ele[31][3] != ele[32][1];
    ele[31][3] != ele[32][2];
    ele[31][3] != ele[32][3];
    ele[31][3] != ele[32][4];
    ele[31][3] != ele[32][5];
    ele[31][3] != ele[33][0];
    ele[31][3] != ele[33][1];
    ele[31][3] != ele[33][2];
    ele[31][3] != ele[33][3];
    ele[31][3] != ele[33][4];
    ele[31][3] != ele[33][5];
    ele[31][3] != ele[34][0];
    ele[31][3] != ele[34][1];
    ele[31][3] != ele[34][2];
    ele[31][3] != ele[34][3];
    ele[31][3] != ele[34][4];
    ele[31][3] != ele[34][5];
    ele[31][3] != ele[35][0];
    ele[31][3] != ele[35][1];
    ele[31][3] != ele[35][2];
    ele[31][3] != ele[35][3];
    ele[31][3] != ele[35][4];
    ele[31][3] != ele[35][5];
    ele[31][30] != ele[31][31];
    ele[31][30] != ele[31][32];
    ele[31][30] != ele[31][33];
    ele[31][30] != ele[31][34];
    ele[31][30] != ele[31][35];
    ele[31][30] != ele[32][30];
    ele[31][30] != ele[32][31];
    ele[31][30] != ele[32][32];
    ele[31][30] != ele[32][33];
    ele[31][30] != ele[32][34];
    ele[31][30] != ele[32][35];
    ele[31][30] != ele[33][30];
    ele[31][30] != ele[33][31];
    ele[31][30] != ele[33][32];
    ele[31][30] != ele[33][33];
    ele[31][30] != ele[33][34];
    ele[31][30] != ele[33][35];
    ele[31][30] != ele[34][30];
    ele[31][30] != ele[34][31];
    ele[31][30] != ele[34][32];
    ele[31][30] != ele[34][33];
    ele[31][30] != ele[34][34];
    ele[31][30] != ele[34][35];
    ele[31][30] != ele[35][30];
    ele[31][30] != ele[35][31];
    ele[31][30] != ele[35][32];
    ele[31][30] != ele[35][33];
    ele[31][30] != ele[35][34];
    ele[31][30] != ele[35][35];
    ele[31][31] != ele[31][32];
    ele[31][31] != ele[31][33];
    ele[31][31] != ele[31][34];
    ele[31][31] != ele[31][35];
    ele[31][31] != ele[32][30];
    ele[31][31] != ele[32][31];
    ele[31][31] != ele[32][32];
    ele[31][31] != ele[32][33];
    ele[31][31] != ele[32][34];
    ele[31][31] != ele[32][35];
    ele[31][31] != ele[33][30];
    ele[31][31] != ele[33][31];
    ele[31][31] != ele[33][32];
    ele[31][31] != ele[33][33];
    ele[31][31] != ele[33][34];
    ele[31][31] != ele[33][35];
    ele[31][31] != ele[34][30];
    ele[31][31] != ele[34][31];
    ele[31][31] != ele[34][32];
    ele[31][31] != ele[34][33];
    ele[31][31] != ele[34][34];
    ele[31][31] != ele[34][35];
    ele[31][31] != ele[35][30];
    ele[31][31] != ele[35][31];
    ele[31][31] != ele[35][32];
    ele[31][31] != ele[35][33];
    ele[31][31] != ele[35][34];
    ele[31][31] != ele[35][35];
    ele[31][32] != ele[31][33];
    ele[31][32] != ele[31][34];
    ele[31][32] != ele[31][35];
    ele[31][32] != ele[32][30];
    ele[31][32] != ele[32][31];
    ele[31][32] != ele[32][32];
    ele[31][32] != ele[32][33];
    ele[31][32] != ele[32][34];
    ele[31][32] != ele[32][35];
    ele[31][32] != ele[33][30];
    ele[31][32] != ele[33][31];
    ele[31][32] != ele[33][32];
    ele[31][32] != ele[33][33];
    ele[31][32] != ele[33][34];
    ele[31][32] != ele[33][35];
    ele[31][32] != ele[34][30];
    ele[31][32] != ele[34][31];
    ele[31][32] != ele[34][32];
    ele[31][32] != ele[34][33];
    ele[31][32] != ele[34][34];
    ele[31][32] != ele[34][35];
    ele[31][32] != ele[35][30];
    ele[31][32] != ele[35][31];
    ele[31][32] != ele[35][32];
    ele[31][32] != ele[35][33];
    ele[31][32] != ele[35][34];
    ele[31][32] != ele[35][35];
    ele[31][33] != ele[31][34];
    ele[31][33] != ele[31][35];
    ele[31][33] != ele[32][30];
    ele[31][33] != ele[32][31];
    ele[31][33] != ele[32][32];
    ele[31][33] != ele[32][33];
    ele[31][33] != ele[32][34];
    ele[31][33] != ele[32][35];
    ele[31][33] != ele[33][30];
    ele[31][33] != ele[33][31];
    ele[31][33] != ele[33][32];
    ele[31][33] != ele[33][33];
    ele[31][33] != ele[33][34];
    ele[31][33] != ele[33][35];
    ele[31][33] != ele[34][30];
    ele[31][33] != ele[34][31];
    ele[31][33] != ele[34][32];
    ele[31][33] != ele[34][33];
    ele[31][33] != ele[34][34];
    ele[31][33] != ele[34][35];
    ele[31][33] != ele[35][30];
    ele[31][33] != ele[35][31];
    ele[31][33] != ele[35][32];
    ele[31][33] != ele[35][33];
    ele[31][33] != ele[35][34];
    ele[31][33] != ele[35][35];
    ele[31][34] != ele[31][35];
    ele[31][34] != ele[32][30];
    ele[31][34] != ele[32][31];
    ele[31][34] != ele[32][32];
    ele[31][34] != ele[32][33];
    ele[31][34] != ele[32][34];
    ele[31][34] != ele[32][35];
    ele[31][34] != ele[33][30];
    ele[31][34] != ele[33][31];
    ele[31][34] != ele[33][32];
    ele[31][34] != ele[33][33];
    ele[31][34] != ele[33][34];
    ele[31][34] != ele[33][35];
    ele[31][34] != ele[34][30];
    ele[31][34] != ele[34][31];
    ele[31][34] != ele[34][32];
    ele[31][34] != ele[34][33];
    ele[31][34] != ele[34][34];
    ele[31][34] != ele[34][35];
    ele[31][34] != ele[35][30];
    ele[31][34] != ele[35][31];
    ele[31][34] != ele[35][32];
    ele[31][34] != ele[35][33];
    ele[31][34] != ele[35][34];
    ele[31][34] != ele[35][35];
    ele[31][35] != ele[32][30];
    ele[31][35] != ele[32][31];
    ele[31][35] != ele[32][32];
    ele[31][35] != ele[32][33];
    ele[31][35] != ele[32][34];
    ele[31][35] != ele[32][35];
    ele[31][35] != ele[33][30];
    ele[31][35] != ele[33][31];
    ele[31][35] != ele[33][32];
    ele[31][35] != ele[33][33];
    ele[31][35] != ele[33][34];
    ele[31][35] != ele[33][35];
    ele[31][35] != ele[34][30];
    ele[31][35] != ele[34][31];
    ele[31][35] != ele[34][32];
    ele[31][35] != ele[34][33];
    ele[31][35] != ele[34][34];
    ele[31][35] != ele[34][35];
    ele[31][35] != ele[35][30];
    ele[31][35] != ele[35][31];
    ele[31][35] != ele[35][32];
    ele[31][35] != ele[35][33];
    ele[31][35] != ele[35][34];
    ele[31][35] != ele[35][35];
    ele[31][4] != ele[31][10];
    ele[31][4] != ele[31][11];
    ele[31][4] != ele[31][12];
    ele[31][4] != ele[31][13];
    ele[31][4] != ele[31][14];
    ele[31][4] != ele[31][15];
    ele[31][4] != ele[31][16];
    ele[31][4] != ele[31][17];
    ele[31][4] != ele[31][18];
    ele[31][4] != ele[31][19];
    ele[31][4] != ele[31][20];
    ele[31][4] != ele[31][21];
    ele[31][4] != ele[31][22];
    ele[31][4] != ele[31][23];
    ele[31][4] != ele[31][24];
    ele[31][4] != ele[31][25];
    ele[31][4] != ele[31][26];
    ele[31][4] != ele[31][27];
    ele[31][4] != ele[31][28];
    ele[31][4] != ele[31][29];
    ele[31][4] != ele[31][30];
    ele[31][4] != ele[31][31];
    ele[31][4] != ele[31][32];
    ele[31][4] != ele[31][33];
    ele[31][4] != ele[31][34];
    ele[31][4] != ele[31][35];
    ele[31][4] != ele[31][5];
    ele[31][4] != ele[31][6];
    ele[31][4] != ele[31][7];
    ele[31][4] != ele[31][8];
    ele[31][4] != ele[31][9];
    ele[31][4] != ele[32][0];
    ele[31][4] != ele[32][1];
    ele[31][4] != ele[32][2];
    ele[31][4] != ele[32][3];
    ele[31][4] != ele[32][4];
    ele[31][4] != ele[32][5];
    ele[31][4] != ele[33][0];
    ele[31][4] != ele[33][1];
    ele[31][4] != ele[33][2];
    ele[31][4] != ele[33][3];
    ele[31][4] != ele[33][4];
    ele[31][4] != ele[33][5];
    ele[31][4] != ele[34][0];
    ele[31][4] != ele[34][1];
    ele[31][4] != ele[34][2];
    ele[31][4] != ele[34][3];
    ele[31][4] != ele[34][4];
    ele[31][4] != ele[34][5];
    ele[31][4] != ele[35][0];
    ele[31][4] != ele[35][1];
    ele[31][4] != ele[35][2];
    ele[31][4] != ele[35][3];
    ele[31][4] != ele[35][4];
    ele[31][4] != ele[35][5];
    ele[31][5] != ele[31][10];
    ele[31][5] != ele[31][11];
    ele[31][5] != ele[31][12];
    ele[31][5] != ele[31][13];
    ele[31][5] != ele[31][14];
    ele[31][5] != ele[31][15];
    ele[31][5] != ele[31][16];
    ele[31][5] != ele[31][17];
    ele[31][5] != ele[31][18];
    ele[31][5] != ele[31][19];
    ele[31][5] != ele[31][20];
    ele[31][5] != ele[31][21];
    ele[31][5] != ele[31][22];
    ele[31][5] != ele[31][23];
    ele[31][5] != ele[31][24];
    ele[31][5] != ele[31][25];
    ele[31][5] != ele[31][26];
    ele[31][5] != ele[31][27];
    ele[31][5] != ele[31][28];
    ele[31][5] != ele[31][29];
    ele[31][5] != ele[31][30];
    ele[31][5] != ele[31][31];
    ele[31][5] != ele[31][32];
    ele[31][5] != ele[31][33];
    ele[31][5] != ele[31][34];
    ele[31][5] != ele[31][35];
    ele[31][5] != ele[31][6];
    ele[31][5] != ele[31][7];
    ele[31][5] != ele[31][8];
    ele[31][5] != ele[31][9];
    ele[31][5] != ele[32][0];
    ele[31][5] != ele[32][1];
    ele[31][5] != ele[32][2];
    ele[31][5] != ele[32][3];
    ele[31][5] != ele[32][4];
    ele[31][5] != ele[32][5];
    ele[31][5] != ele[33][0];
    ele[31][5] != ele[33][1];
    ele[31][5] != ele[33][2];
    ele[31][5] != ele[33][3];
    ele[31][5] != ele[33][4];
    ele[31][5] != ele[33][5];
    ele[31][5] != ele[34][0];
    ele[31][5] != ele[34][1];
    ele[31][5] != ele[34][2];
    ele[31][5] != ele[34][3];
    ele[31][5] != ele[34][4];
    ele[31][5] != ele[34][5];
    ele[31][5] != ele[35][0];
    ele[31][5] != ele[35][1];
    ele[31][5] != ele[35][2];
    ele[31][5] != ele[35][3];
    ele[31][5] != ele[35][4];
    ele[31][5] != ele[35][5];
    ele[31][6] != ele[31][10];
    ele[31][6] != ele[31][11];
    ele[31][6] != ele[31][12];
    ele[31][6] != ele[31][13];
    ele[31][6] != ele[31][14];
    ele[31][6] != ele[31][15];
    ele[31][6] != ele[31][16];
    ele[31][6] != ele[31][17];
    ele[31][6] != ele[31][18];
    ele[31][6] != ele[31][19];
    ele[31][6] != ele[31][20];
    ele[31][6] != ele[31][21];
    ele[31][6] != ele[31][22];
    ele[31][6] != ele[31][23];
    ele[31][6] != ele[31][24];
    ele[31][6] != ele[31][25];
    ele[31][6] != ele[31][26];
    ele[31][6] != ele[31][27];
    ele[31][6] != ele[31][28];
    ele[31][6] != ele[31][29];
    ele[31][6] != ele[31][30];
    ele[31][6] != ele[31][31];
    ele[31][6] != ele[31][32];
    ele[31][6] != ele[31][33];
    ele[31][6] != ele[31][34];
    ele[31][6] != ele[31][35];
    ele[31][6] != ele[31][7];
    ele[31][6] != ele[31][8];
    ele[31][6] != ele[31][9];
    ele[31][6] != ele[32][10];
    ele[31][6] != ele[32][11];
    ele[31][6] != ele[32][6];
    ele[31][6] != ele[32][7];
    ele[31][6] != ele[32][8];
    ele[31][6] != ele[32][9];
    ele[31][6] != ele[33][10];
    ele[31][6] != ele[33][11];
    ele[31][6] != ele[33][6];
    ele[31][6] != ele[33][7];
    ele[31][6] != ele[33][8];
    ele[31][6] != ele[33][9];
    ele[31][6] != ele[34][10];
    ele[31][6] != ele[34][11];
    ele[31][6] != ele[34][6];
    ele[31][6] != ele[34][7];
    ele[31][6] != ele[34][8];
    ele[31][6] != ele[34][9];
    ele[31][6] != ele[35][10];
    ele[31][6] != ele[35][11];
    ele[31][6] != ele[35][6];
    ele[31][6] != ele[35][7];
    ele[31][6] != ele[35][8];
    ele[31][6] != ele[35][9];
    ele[31][7] != ele[31][10];
    ele[31][7] != ele[31][11];
    ele[31][7] != ele[31][12];
    ele[31][7] != ele[31][13];
    ele[31][7] != ele[31][14];
    ele[31][7] != ele[31][15];
    ele[31][7] != ele[31][16];
    ele[31][7] != ele[31][17];
    ele[31][7] != ele[31][18];
    ele[31][7] != ele[31][19];
    ele[31][7] != ele[31][20];
    ele[31][7] != ele[31][21];
    ele[31][7] != ele[31][22];
    ele[31][7] != ele[31][23];
    ele[31][7] != ele[31][24];
    ele[31][7] != ele[31][25];
    ele[31][7] != ele[31][26];
    ele[31][7] != ele[31][27];
    ele[31][7] != ele[31][28];
    ele[31][7] != ele[31][29];
    ele[31][7] != ele[31][30];
    ele[31][7] != ele[31][31];
    ele[31][7] != ele[31][32];
    ele[31][7] != ele[31][33];
    ele[31][7] != ele[31][34];
    ele[31][7] != ele[31][35];
    ele[31][7] != ele[31][8];
    ele[31][7] != ele[31][9];
    ele[31][7] != ele[32][10];
    ele[31][7] != ele[32][11];
    ele[31][7] != ele[32][6];
    ele[31][7] != ele[32][7];
    ele[31][7] != ele[32][8];
    ele[31][7] != ele[32][9];
    ele[31][7] != ele[33][10];
    ele[31][7] != ele[33][11];
    ele[31][7] != ele[33][6];
    ele[31][7] != ele[33][7];
    ele[31][7] != ele[33][8];
    ele[31][7] != ele[33][9];
    ele[31][7] != ele[34][10];
    ele[31][7] != ele[34][11];
    ele[31][7] != ele[34][6];
    ele[31][7] != ele[34][7];
    ele[31][7] != ele[34][8];
    ele[31][7] != ele[34][9];
    ele[31][7] != ele[35][10];
    ele[31][7] != ele[35][11];
    ele[31][7] != ele[35][6];
    ele[31][7] != ele[35][7];
    ele[31][7] != ele[35][8];
    ele[31][7] != ele[35][9];
    ele[31][8] != ele[31][10];
    ele[31][8] != ele[31][11];
    ele[31][8] != ele[31][12];
    ele[31][8] != ele[31][13];
    ele[31][8] != ele[31][14];
    ele[31][8] != ele[31][15];
    ele[31][8] != ele[31][16];
    ele[31][8] != ele[31][17];
    ele[31][8] != ele[31][18];
    ele[31][8] != ele[31][19];
    ele[31][8] != ele[31][20];
    ele[31][8] != ele[31][21];
    ele[31][8] != ele[31][22];
    ele[31][8] != ele[31][23];
    ele[31][8] != ele[31][24];
    ele[31][8] != ele[31][25];
    ele[31][8] != ele[31][26];
    ele[31][8] != ele[31][27];
    ele[31][8] != ele[31][28];
    ele[31][8] != ele[31][29];
    ele[31][8] != ele[31][30];
    ele[31][8] != ele[31][31];
    ele[31][8] != ele[31][32];
    ele[31][8] != ele[31][33];
    ele[31][8] != ele[31][34];
    ele[31][8] != ele[31][35];
    ele[31][8] != ele[31][9];
    ele[31][8] != ele[32][10];
    ele[31][8] != ele[32][11];
    ele[31][8] != ele[32][6];
    ele[31][8] != ele[32][7];
    ele[31][8] != ele[32][8];
    ele[31][8] != ele[32][9];
    ele[31][8] != ele[33][10];
    ele[31][8] != ele[33][11];
    ele[31][8] != ele[33][6];
    ele[31][8] != ele[33][7];
    ele[31][8] != ele[33][8];
    ele[31][8] != ele[33][9];
    ele[31][8] != ele[34][10];
    ele[31][8] != ele[34][11];
    ele[31][8] != ele[34][6];
    ele[31][8] != ele[34][7];
    ele[31][8] != ele[34][8];
    ele[31][8] != ele[34][9];
    ele[31][8] != ele[35][10];
    ele[31][8] != ele[35][11];
    ele[31][8] != ele[35][6];
    ele[31][8] != ele[35][7];
    ele[31][8] != ele[35][8];
    ele[31][8] != ele[35][9];
    ele[31][9] != ele[31][10];
    ele[31][9] != ele[31][11];
    ele[31][9] != ele[31][12];
    ele[31][9] != ele[31][13];
    ele[31][9] != ele[31][14];
    ele[31][9] != ele[31][15];
    ele[31][9] != ele[31][16];
    ele[31][9] != ele[31][17];
    ele[31][9] != ele[31][18];
    ele[31][9] != ele[31][19];
    ele[31][9] != ele[31][20];
    ele[31][9] != ele[31][21];
    ele[31][9] != ele[31][22];
    ele[31][9] != ele[31][23];
    ele[31][9] != ele[31][24];
    ele[31][9] != ele[31][25];
    ele[31][9] != ele[31][26];
    ele[31][9] != ele[31][27];
    ele[31][9] != ele[31][28];
    ele[31][9] != ele[31][29];
    ele[31][9] != ele[31][30];
    ele[31][9] != ele[31][31];
    ele[31][9] != ele[31][32];
    ele[31][9] != ele[31][33];
    ele[31][9] != ele[31][34];
    ele[31][9] != ele[31][35];
    ele[31][9] != ele[32][10];
    ele[31][9] != ele[32][11];
    ele[31][9] != ele[32][6];
    ele[31][9] != ele[32][7];
    ele[31][9] != ele[32][8];
    ele[31][9] != ele[32][9];
    ele[31][9] != ele[33][10];
    ele[31][9] != ele[33][11];
    ele[31][9] != ele[33][6];
    ele[31][9] != ele[33][7];
    ele[31][9] != ele[33][8];
    ele[31][9] != ele[33][9];
    ele[31][9] != ele[34][10];
    ele[31][9] != ele[34][11];
    ele[31][9] != ele[34][6];
    ele[31][9] != ele[34][7];
    ele[31][9] != ele[34][8];
    ele[31][9] != ele[34][9];
    ele[31][9] != ele[35][10];
    ele[31][9] != ele[35][11];
    ele[31][9] != ele[35][6];
    ele[31][9] != ele[35][7];
    ele[31][9] != ele[35][8];
    ele[31][9] != ele[35][9];
    ele[32][0] != ele[32][1];
    ele[32][0] != ele[32][10];
    ele[32][0] != ele[32][11];
    ele[32][0] != ele[32][12];
    ele[32][0] != ele[32][13];
    ele[32][0] != ele[32][14];
    ele[32][0] != ele[32][15];
    ele[32][0] != ele[32][16];
    ele[32][0] != ele[32][17];
    ele[32][0] != ele[32][18];
    ele[32][0] != ele[32][19];
    ele[32][0] != ele[32][2];
    ele[32][0] != ele[32][20];
    ele[32][0] != ele[32][21];
    ele[32][0] != ele[32][22];
    ele[32][0] != ele[32][23];
    ele[32][0] != ele[32][24];
    ele[32][0] != ele[32][25];
    ele[32][0] != ele[32][26];
    ele[32][0] != ele[32][27];
    ele[32][0] != ele[32][28];
    ele[32][0] != ele[32][29];
    ele[32][0] != ele[32][3];
    ele[32][0] != ele[32][30];
    ele[32][0] != ele[32][31];
    ele[32][0] != ele[32][32];
    ele[32][0] != ele[32][33];
    ele[32][0] != ele[32][34];
    ele[32][0] != ele[32][35];
    ele[32][0] != ele[32][4];
    ele[32][0] != ele[32][5];
    ele[32][0] != ele[32][6];
    ele[32][0] != ele[32][7];
    ele[32][0] != ele[32][8];
    ele[32][0] != ele[32][9];
    ele[32][0] != ele[33][0];
    ele[32][0] != ele[33][1];
    ele[32][0] != ele[33][2];
    ele[32][0] != ele[33][3];
    ele[32][0] != ele[33][4];
    ele[32][0] != ele[33][5];
    ele[32][0] != ele[34][0];
    ele[32][0] != ele[34][1];
    ele[32][0] != ele[34][2];
    ele[32][0] != ele[34][3];
    ele[32][0] != ele[34][4];
    ele[32][0] != ele[34][5];
    ele[32][0] != ele[35][0];
    ele[32][0] != ele[35][1];
    ele[32][0] != ele[35][2];
    ele[32][0] != ele[35][3];
    ele[32][0] != ele[35][4];
    ele[32][0] != ele[35][5];
    ele[32][1] != ele[32][10];
    ele[32][1] != ele[32][11];
    ele[32][1] != ele[32][12];
    ele[32][1] != ele[32][13];
    ele[32][1] != ele[32][14];
    ele[32][1] != ele[32][15];
    ele[32][1] != ele[32][16];
    ele[32][1] != ele[32][17];
    ele[32][1] != ele[32][18];
    ele[32][1] != ele[32][19];
    ele[32][1] != ele[32][2];
    ele[32][1] != ele[32][20];
    ele[32][1] != ele[32][21];
    ele[32][1] != ele[32][22];
    ele[32][1] != ele[32][23];
    ele[32][1] != ele[32][24];
    ele[32][1] != ele[32][25];
    ele[32][1] != ele[32][26];
    ele[32][1] != ele[32][27];
    ele[32][1] != ele[32][28];
    ele[32][1] != ele[32][29];
    ele[32][1] != ele[32][3];
    ele[32][1] != ele[32][30];
    ele[32][1] != ele[32][31];
    ele[32][1] != ele[32][32];
    ele[32][1] != ele[32][33];
    ele[32][1] != ele[32][34];
    ele[32][1] != ele[32][35];
    ele[32][1] != ele[32][4];
    ele[32][1] != ele[32][5];
    ele[32][1] != ele[32][6];
    ele[32][1] != ele[32][7];
    ele[32][1] != ele[32][8];
    ele[32][1] != ele[32][9];
    ele[32][1] != ele[33][0];
    ele[32][1] != ele[33][1];
    ele[32][1] != ele[33][2];
    ele[32][1] != ele[33][3];
    ele[32][1] != ele[33][4];
    ele[32][1] != ele[33][5];
    ele[32][1] != ele[34][0];
    ele[32][1] != ele[34][1];
    ele[32][1] != ele[34][2];
    ele[32][1] != ele[34][3];
    ele[32][1] != ele[34][4];
    ele[32][1] != ele[34][5];
    ele[32][1] != ele[35][0];
    ele[32][1] != ele[35][1];
    ele[32][1] != ele[35][2];
    ele[32][1] != ele[35][3];
    ele[32][1] != ele[35][4];
    ele[32][1] != ele[35][5];
    ele[32][10] != ele[32][11];
    ele[32][10] != ele[32][12];
    ele[32][10] != ele[32][13];
    ele[32][10] != ele[32][14];
    ele[32][10] != ele[32][15];
    ele[32][10] != ele[32][16];
    ele[32][10] != ele[32][17];
    ele[32][10] != ele[32][18];
    ele[32][10] != ele[32][19];
    ele[32][10] != ele[32][20];
    ele[32][10] != ele[32][21];
    ele[32][10] != ele[32][22];
    ele[32][10] != ele[32][23];
    ele[32][10] != ele[32][24];
    ele[32][10] != ele[32][25];
    ele[32][10] != ele[32][26];
    ele[32][10] != ele[32][27];
    ele[32][10] != ele[32][28];
    ele[32][10] != ele[32][29];
    ele[32][10] != ele[32][30];
    ele[32][10] != ele[32][31];
    ele[32][10] != ele[32][32];
    ele[32][10] != ele[32][33];
    ele[32][10] != ele[32][34];
    ele[32][10] != ele[32][35];
    ele[32][10] != ele[33][10];
    ele[32][10] != ele[33][11];
    ele[32][10] != ele[33][6];
    ele[32][10] != ele[33][7];
    ele[32][10] != ele[33][8];
    ele[32][10] != ele[33][9];
    ele[32][10] != ele[34][10];
    ele[32][10] != ele[34][11];
    ele[32][10] != ele[34][6];
    ele[32][10] != ele[34][7];
    ele[32][10] != ele[34][8];
    ele[32][10] != ele[34][9];
    ele[32][10] != ele[35][10];
    ele[32][10] != ele[35][11];
    ele[32][10] != ele[35][6];
    ele[32][10] != ele[35][7];
    ele[32][10] != ele[35][8];
    ele[32][10] != ele[35][9];
    ele[32][11] != ele[32][12];
    ele[32][11] != ele[32][13];
    ele[32][11] != ele[32][14];
    ele[32][11] != ele[32][15];
    ele[32][11] != ele[32][16];
    ele[32][11] != ele[32][17];
    ele[32][11] != ele[32][18];
    ele[32][11] != ele[32][19];
    ele[32][11] != ele[32][20];
    ele[32][11] != ele[32][21];
    ele[32][11] != ele[32][22];
    ele[32][11] != ele[32][23];
    ele[32][11] != ele[32][24];
    ele[32][11] != ele[32][25];
    ele[32][11] != ele[32][26];
    ele[32][11] != ele[32][27];
    ele[32][11] != ele[32][28];
    ele[32][11] != ele[32][29];
    ele[32][11] != ele[32][30];
    ele[32][11] != ele[32][31];
    ele[32][11] != ele[32][32];
    ele[32][11] != ele[32][33];
    ele[32][11] != ele[32][34];
    ele[32][11] != ele[32][35];
    ele[32][11] != ele[33][10];
    ele[32][11] != ele[33][11];
    ele[32][11] != ele[33][6];
    ele[32][11] != ele[33][7];
    ele[32][11] != ele[33][8];
    ele[32][11] != ele[33][9];
    ele[32][11] != ele[34][10];
    ele[32][11] != ele[34][11];
    ele[32][11] != ele[34][6];
    ele[32][11] != ele[34][7];
    ele[32][11] != ele[34][8];
    ele[32][11] != ele[34][9];
    ele[32][11] != ele[35][10];
    ele[32][11] != ele[35][11];
    ele[32][11] != ele[35][6];
    ele[32][11] != ele[35][7];
    ele[32][11] != ele[35][8];
    ele[32][11] != ele[35][9];
    ele[32][12] != ele[32][13];
    ele[32][12] != ele[32][14];
    ele[32][12] != ele[32][15];
    ele[32][12] != ele[32][16];
    ele[32][12] != ele[32][17];
    ele[32][12] != ele[32][18];
    ele[32][12] != ele[32][19];
    ele[32][12] != ele[32][20];
    ele[32][12] != ele[32][21];
    ele[32][12] != ele[32][22];
    ele[32][12] != ele[32][23];
    ele[32][12] != ele[32][24];
    ele[32][12] != ele[32][25];
    ele[32][12] != ele[32][26];
    ele[32][12] != ele[32][27];
    ele[32][12] != ele[32][28];
    ele[32][12] != ele[32][29];
    ele[32][12] != ele[32][30];
    ele[32][12] != ele[32][31];
    ele[32][12] != ele[32][32];
    ele[32][12] != ele[32][33];
    ele[32][12] != ele[32][34];
    ele[32][12] != ele[32][35];
    ele[32][12] != ele[33][12];
    ele[32][12] != ele[33][13];
    ele[32][12] != ele[33][14];
    ele[32][12] != ele[33][15];
    ele[32][12] != ele[33][16];
    ele[32][12] != ele[33][17];
    ele[32][12] != ele[34][12];
    ele[32][12] != ele[34][13];
    ele[32][12] != ele[34][14];
    ele[32][12] != ele[34][15];
    ele[32][12] != ele[34][16];
    ele[32][12] != ele[34][17];
    ele[32][12] != ele[35][12];
    ele[32][12] != ele[35][13];
    ele[32][12] != ele[35][14];
    ele[32][12] != ele[35][15];
    ele[32][12] != ele[35][16];
    ele[32][12] != ele[35][17];
    ele[32][13] != ele[32][14];
    ele[32][13] != ele[32][15];
    ele[32][13] != ele[32][16];
    ele[32][13] != ele[32][17];
    ele[32][13] != ele[32][18];
    ele[32][13] != ele[32][19];
    ele[32][13] != ele[32][20];
    ele[32][13] != ele[32][21];
    ele[32][13] != ele[32][22];
    ele[32][13] != ele[32][23];
    ele[32][13] != ele[32][24];
    ele[32][13] != ele[32][25];
    ele[32][13] != ele[32][26];
    ele[32][13] != ele[32][27];
    ele[32][13] != ele[32][28];
    ele[32][13] != ele[32][29];
    ele[32][13] != ele[32][30];
    ele[32][13] != ele[32][31];
    ele[32][13] != ele[32][32];
    ele[32][13] != ele[32][33];
    ele[32][13] != ele[32][34];
    ele[32][13] != ele[32][35];
    ele[32][13] != ele[33][12];
    ele[32][13] != ele[33][13];
    ele[32][13] != ele[33][14];
    ele[32][13] != ele[33][15];
    ele[32][13] != ele[33][16];
    ele[32][13] != ele[33][17];
    ele[32][13] != ele[34][12];
    ele[32][13] != ele[34][13];
    ele[32][13] != ele[34][14];
    ele[32][13] != ele[34][15];
    ele[32][13] != ele[34][16];
    ele[32][13] != ele[34][17];
    ele[32][13] != ele[35][12];
    ele[32][13] != ele[35][13];
    ele[32][13] != ele[35][14];
    ele[32][13] != ele[35][15];
    ele[32][13] != ele[35][16];
    ele[32][13] != ele[35][17];
    ele[32][14] != ele[32][15];
    ele[32][14] != ele[32][16];
    ele[32][14] != ele[32][17];
    ele[32][14] != ele[32][18];
    ele[32][14] != ele[32][19];
    ele[32][14] != ele[32][20];
    ele[32][14] != ele[32][21];
    ele[32][14] != ele[32][22];
    ele[32][14] != ele[32][23];
    ele[32][14] != ele[32][24];
    ele[32][14] != ele[32][25];
    ele[32][14] != ele[32][26];
    ele[32][14] != ele[32][27];
    ele[32][14] != ele[32][28];
    ele[32][14] != ele[32][29];
    ele[32][14] != ele[32][30];
    ele[32][14] != ele[32][31];
    ele[32][14] != ele[32][32];
    ele[32][14] != ele[32][33];
    ele[32][14] != ele[32][34];
    ele[32][14] != ele[32][35];
    ele[32][14] != ele[33][12];
    ele[32][14] != ele[33][13];
    ele[32][14] != ele[33][14];
    ele[32][14] != ele[33][15];
    ele[32][14] != ele[33][16];
    ele[32][14] != ele[33][17];
    ele[32][14] != ele[34][12];
    ele[32][14] != ele[34][13];
    ele[32][14] != ele[34][14];
    ele[32][14] != ele[34][15];
    ele[32][14] != ele[34][16];
    ele[32][14] != ele[34][17];
    ele[32][14] != ele[35][12];
    ele[32][14] != ele[35][13];
    ele[32][14] != ele[35][14];
    ele[32][14] != ele[35][15];
    ele[32][14] != ele[35][16];
    ele[32][14] != ele[35][17];
    ele[32][15] != ele[32][16];
    ele[32][15] != ele[32][17];
    ele[32][15] != ele[32][18];
    ele[32][15] != ele[32][19];
    ele[32][15] != ele[32][20];
    ele[32][15] != ele[32][21];
    ele[32][15] != ele[32][22];
    ele[32][15] != ele[32][23];
    ele[32][15] != ele[32][24];
    ele[32][15] != ele[32][25];
    ele[32][15] != ele[32][26];
    ele[32][15] != ele[32][27];
    ele[32][15] != ele[32][28];
    ele[32][15] != ele[32][29];
    ele[32][15] != ele[32][30];
    ele[32][15] != ele[32][31];
    ele[32][15] != ele[32][32];
    ele[32][15] != ele[32][33];
    ele[32][15] != ele[32][34];
    ele[32][15] != ele[32][35];
    ele[32][15] != ele[33][12];
    ele[32][15] != ele[33][13];
    ele[32][15] != ele[33][14];
    ele[32][15] != ele[33][15];
    ele[32][15] != ele[33][16];
    ele[32][15] != ele[33][17];
    ele[32][15] != ele[34][12];
    ele[32][15] != ele[34][13];
    ele[32][15] != ele[34][14];
    ele[32][15] != ele[34][15];
    ele[32][15] != ele[34][16];
    ele[32][15] != ele[34][17];
    ele[32][15] != ele[35][12];
    ele[32][15] != ele[35][13];
    ele[32][15] != ele[35][14];
    ele[32][15] != ele[35][15];
    ele[32][15] != ele[35][16];
    ele[32][15] != ele[35][17];
    ele[32][16] != ele[32][17];
    ele[32][16] != ele[32][18];
    ele[32][16] != ele[32][19];
    ele[32][16] != ele[32][20];
    ele[32][16] != ele[32][21];
    ele[32][16] != ele[32][22];
    ele[32][16] != ele[32][23];
    ele[32][16] != ele[32][24];
    ele[32][16] != ele[32][25];
    ele[32][16] != ele[32][26];
    ele[32][16] != ele[32][27];
    ele[32][16] != ele[32][28];
    ele[32][16] != ele[32][29];
    ele[32][16] != ele[32][30];
    ele[32][16] != ele[32][31];
    ele[32][16] != ele[32][32];
    ele[32][16] != ele[32][33];
    ele[32][16] != ele[32][34];
    ele[32][16] != ele[32][35];
    ele[32][16] != ele[33][12];
    ele[32][16] != ele[33][13];
    ele[32][16] != ele[33][14];
    ele[32][16] != ele[33][15];
    ele[32][16] != ele[33][16];
    ele[32][16] != ele[33][17];
    ele[32][16] != ele[34][12];
    ele[32][16] != ele[34][13];
    ele[32][16] != ele[34][14];
    ele[32][16] != ele[34][15];
    ele[32][16] != ele[34][16];
    ele[32][16] != ele[34][17];
    ele[32][16] != ele[35][12];
    ele[32][16] != ele[35][13];
    ele[32][16] != ele[35][14];
    ele[32][16] != ele[35][15];
    ele[32][16] != ele[35][16];
    ele[32][16] != ele[35][17];
    ele[32][17] != ele[32][18];
    ele[32][17] != ele[32][19];
    ele[32][17] != ele[32][20];
    ele[32][17] != ele[32][21];
    ele[32][17] != ele[32][22];
    ele[32][17] != ele[32][23];
    ele[32][17] != ele[32][24];
    ele[32][17] != ele[32][25];
    ele[32][17] != ele[32][26];
    ele[32][17] != ele[32][27];
    ele[32][17] != ele[32][28];
    ele[32][17] != ele[32][29];
    ele[32][17] != ele[32][30];
    ele[32][17] != ele[32][31];
    ele[32][17] != ele[32][32];
    ele[32][17] != ele[32][33];
    ele[32][17] != ele[32][34];
    ele[32][17] != ele[32][35];
    ele[32][17] != ele[33][12];
    ele[32][17] != ele[33][13];
    ele[32][17] != ele[33][14];
    ele[32][17] != ele[33][15];
    ele[32][17] != ele[33][16];
    ele[32][17] != ele[33][17];
    ele[32][17] != ele[34][12];
    ele[32][17] != ele[34][13];
    ele[32][17] != ele[34][14];
    ele[32][17] != ele[34][15];
    ele[32][17] != ele[34][16];
    ele[32][17] != ele[34][17];
    ele[32][17] != ele[35][12];
    ele[32][17] != ele[35][13];
    ele[32][17] != ele[35][14];
    ele[32][17] != ele[35][15];
    ele[32][17] != ele[35][16];
    ele[32][17] != ele[35][17];
    ele[32][18] != ele[32][19];
    ele[32][18] != ele[32][20];
    ele[32][18] != ele[32][21];
    ele[32][18] != ele[32][22];
    ele[32][18] != ele[32][23];
    ele[32][18] != ele[32][24];
    ele[32][18] != ele[32][25];
    ele[32][18] != ele[32][26];
    ele[32][18] != ele[32][27];
    ele[32][18] != ele[32][28];
    ele[32][18] != ele[32][29];
    ele[32][18] != ele[32][30];
    ele[32][18] != ele[32][31];
    ele[32][18] != ele[32][32];
    ele[32][18] != ele[32][33];
    ele[32][18] != ele[32][34];
    ele[32][18] != ele[32][35];
    ele[32][18] != ele[33][18];
    ele[32][18] != ele[33][19];
    ele[32][18] != ele[33][20];
    ele[32][18] != ele[33][21];
    ele[32][18] != ele[33][22];
    ele[32][18] != ele[33][23];
    ele[32][18] != ele[34][18];
    ele[32][18] != ele[34][19];
    ele[32][18] != ele[34][20];
    ele[32][18] != ele[34][21];
    ele[32][18] != ele[34][22];
    ele[32][18] != ele[34][23];
    ele[32][18] != ele[35][18];
    ele[32][18] != ele[35][19];
    ele[32][18] != ele[35][20];
    ele[32][18] != ele[35][21];
    ele[32][18] != ele[35][22];
    ele[32][18] != ele[35][23];
    ele[32][19] != ele[32][20];
    ele[32][19] != ele[32][21];
    ele[32][19] != ele[32][22];
    ele[32][19] != ele[32][23];
    ele[32][19] != ele[32][24];
    ele[32][19] != ele[32][25];
    ele[32][19] != ele[32][26];
    ele[32][19] != ele[32][27];
    ele[32][19] != ele[32][28];
    ele[32][19] != ele[32][29];
    ele[32][19] != ele[32][30];
    ele[32][19] != ele[32][31];
    ele[32][19] != ele[32][32];
    ele[32][19] != ele[32][33];
    ele[32][19] != ele[32][34];
    ele[32][19] != ele[32][35];
    ele[32][19] != ele[33][18];
    ele[32][19] != ele[33][19];
    ele[32][19] != ele[33][20];
    ele[32][19] != ele[33][21];
    ele[32][19] != ele[33][22];
    ele[32][19] != ele[33][23];
    ele[32][19] != ele[34][18];
    ele[32][19] != ele[34][19];
    ele[32][19] != ele[34][20];
    ele[32][19] != ele[34][21];
    ele[32][19] != ele[34][22];
    ele[32][19] != ele[34][23];
    ele[32][19] != ele[35][18];
    ele[32][19] != ele[35][19];
    ele[32][19] != ele[35][20];
    ele[32][19] != ele[35][21];
    ele[32][19] != ele[35][22];
    ele[32][19] != ele[35][23];
    ele[32][2] != ele[32][10];
    ele[32][2] != ele[32][11];
    ele[32][2] != ele[32][12];
    ele[32][2] != ele[32][13];
    ele[32][2] != ele[32][14];
    ele[32][2] != ele[32][15];
    ele[32][2] != ele[32][16];
    ele[32][2] != ele[32][17];
    ele[32][2] != ele[32][18];
    ele[32][2] != ele[32][19];
    ele[32][2] != ele[32][20];
    ele[32][2] != ele[32][21];
    ele[32][2] != ele[32][22];
    ele[32][2] != ele[32][23];
    ele[32][2] != ele[32][24];
    ele[32][2] != ele[32][25];
    ele[32][2] != ele[32][26];
    ele[32][2] != ele[32][27];
    ele[32][2] != ele[32][28];
    ele[32][2] != ele[32][29];
    ele[32][2] != ele[32][3];
    ele[32][2] != ele[32][30];
    ele[32][2] != ele[32][31];
    ele[32][2] != ele[32][32];
    ele[32][2] != ele[32][33];
    ele[32][2] != ele[32][34];
    ele[32][2] != ele[32][35];
    ele[32][2] != ele[32][4];
    ele[32][2] != ele[32][5];
    ele[32][2] != ele[32][6];
    ele[32][2] != ele[32][7];
    ele[32][2] != ele[32][8];
    ele[32][2] != ele[32][9];
    ele[32][2] != ele[33][0];
    ele[32][2] != ele[33][1];
    ele[32][2] != ele[33][2];
    ele[32][2] != ele[33][3];
    ele[32][2] != ele[33][4];
    ele[32][2] != ele[33][5];
    ele[32][2] != ele[34][0];
    ele[32][2] != ele[34][1];
    ele[32][2] != ele[34][2];
    ele[32][2] != ele[34][3];
    ele[32][2] != ele[34][4];
    ele[32][2] != ele[34][5];
    ele[32][2] != ele[35][0];
    ele[32][2] != ele[35][1];
    ele[32][2] != ele[35][2];
    ele[32][2] != ele[35][3];
    ele[32][2] != ele[35][4];
    ele[32][2] != ele[35][5];
    ele[32][20] != ele[32][21];
    ele[32][20] != ele[32][22];
    ele[32][20] != ele[32][23];
    ele[32][20] != ele[32][24];
    ele[32][20] != ele[32][25];
    ele[32][20] != ele[32][26];
    ele[32][20] != ele[32][27];
    ele[32][20] != ele[32][28];
    ele[32][20] != ele[32][29];
    ele[32][20] != ele[32][30];
    ele[32][20] != ele[32][31];
    ele[32][20] != ele[32][32];
    ele[32][20] != ele[32][33];
    ele[32][20] != ele[32][34];
    ele[32][20] != ele[32][35];
    ele[32][20] != ele[33][18];
    ele[32][20] != ele[33][19];
    ele[32][20] != ele[33][20];
    ele[32][20] != ele[33][21];
    ele[32][20] != ele[33][22];
    ele[32][20] != ele[33][23];
    ele[32][20] != ele[34][18];
    ele[32][20] != ele[34][19];
    ele[32][20] != ele[34][20];
    ele[32][20] != ele[34][21];
    ele[32][20] != ele[34][22];
    ele[32][20] != ele[34][23];
    ele[32][20] != ele[35][18];
    ele[32][20] != ele[35][19];
    ele[32][20] != ele[35][20];
    ele[32][20] != ele[35][21];
    ele[32][20] != ele[35][22];
    ele[32][20] != ele[35][23];
    ele[32][21] != ele[32][22];
    ele[32][21] != ele[32][23];
    ele[32][21] != ele[32][24];
    ele[32][21] != ele[32][25];
    ele[32][21] != ele[32][26];
    ele[32][21] != ele[32][27];
    ele[32][21] != ele[32][28];
    ele[32][21] != ele[32][29];
    ele[32][21] != ele[32][30];
    ele[32][21] != ele[32][31];
    ele[32][21] != ele[32][32];
    ele[32][21] != ele[32][33];
    ele[32][21] != ele[32][34];
    ele[32][21] != ele[32][35];
    ele[32][21] != ele[33][18];
    ele[32][21] != ele[33][19];
    ele[32][21] != ele[33][20];
    ele[32][21] != ele[33][21];
    ele[32][21] != ele[33][22];
    ele[32][21] != ele[33][23];
    ele[32][21] != ele[34][18];
    ele[32][21] != ele[34][19];
    ele[32][21] != ele[34][20];
    ele[32][21] != ele[34][21];
    ele[32][21] != ele[34][22];
    ele[32][21] != ele[34][23];
    ele[32][21] != ele[35][18];
    ele[32][21] != ele[35][19];
    ele[32][21] != ele[35][20];
    ele[32][21] != ele[35][21];
    ele[32][21] != ele[35][22];
    ele[32][21] != ele[35][23];
    ele[32][22] != ele[32][23];
    ele[32][22] != ele[32][24];
    ele[32][22] != ele[32][25];
    ele[32][22] != ele[32][26];
    ele[32][22] != ele[32][27];
    ele[32][22] != ele[32][28];
    ele[32][22] != ele[32][29];
    ele[32][22] != ele[32][30];
    ele[32][22] != ele[32][31];
    ele[32][22] != ele[32][32];
    ele[32][22] != ele[32][33];
    ele[32][22] != ele[32][34];
    ele[32][22] != ele[32][35];
    ele[32][22] != ele[33][18];
    ele[32][22] != ele[33][19];
    ele[32][22] != ele[33][20];
    ele[32][22] != ele[33][21];
    ele[32][22] != ele[33][22];
    ele[32][22] != ele[33][23];
    ele[32][22] != ele[34][18];
    ele[32][22] != ele[34][19];
    ele[32][22] != ele[34][20];
    ele[32][22] != ele[34][21];
    ele[32][22] != ele[34][22];
    ele[32][22] != ele[34][23];
    ele[32][22] != ele[35][18];
    ele[32][22] != ele[35][19];
    ele[32][22] != ele[35][20];
    ele[32][22] != ele[35][21];
    ele[32][22] != ele[35][22];
    ele[32][22] != ele[35][23];
    ele[32][23] != ele[32][24];
    ele[32][23] != ele[32][25];
    ele[32][23] != ele[32][26];
    ele[32][23] != ele[32][27];
    ele[32][23] != ele[32][28];
    ele[32][23] != ele[32][29];
    ele[32][23] != ele[32][30];
    ele[32][23] != ele[32][31];
    ele[32][23] != ele[32][32];
    ele[32][23] != ele[32][33];
    ele[32][23] != ele[32][34];
    ele[32][23] != ele[32][35];
    ele[32][23] != ele[33][18];
    ele[32][23] != ele[33][19];
    ele[32][23] != ele[33][20];
    ele[32][23] != ele[33][21];
    ele[32][23] != ele[33][22];
    ele[32][23] != ele[33][23];
    ele[32][23] != ele[34][18];
    ele[32][23] != ele[34][19];
    ele[32][23] != ele[34][20];
    ele[32][23] != ele[34][21];
    ele[32][23] != ele[34][22];
    ele[32][23] != ele[34][23];
    ele[32][23] != ele[35][18];
    ele[32][23] != ele[35][19];
    ele[32][23] != ele[35][20];
    ele[32][23] != ele[35][21];
    ele[32][23] != ele[35][22];
    ele[32][23] != ele[35][23];
    ele[32][24] != ele[32][25];
    ele[32][24] != ele[32][26];
    ele[32][24] != ele[32][27];
    ele[32][24] != ele[32][28];
    ele[32][24] != ele[32][29];
    ele[32][24] != ele[32][30];
    ele[32][24] != ele[32][31];
    ele[32][24] != ele[32][32];
    ele[32][24] != ele[32][33];
    ele[32][24] != ele[32][34];
    ele[32][24] != ele[32][35];
    ele[32][24] != ele[33][24];
    ele[32][24] != ele[33][25];
    ele[32][24] != ele[33][26];
    ele[32][24] != ele[33][27];
    ele[32][24] != ele[33][28];
    ele[32][24] != ele[33][29];
    ele[32][24] != ele[34][24];
    ele[32][24] != ele[34][25];
    ele[32][24] != ele[34][26];
    ele[32][24] != ele[34][27];
    ele[32][24] != ele[34][28];
    ele[32][24] != ele[34][29];
    ele[32][24] != ele[35][24];
    ele[32][24] != ele[35][25];
    ele[32][24] != ele[35][26];
    ele[32][24] != ele[35][27];
    ele[32][24] != ele[35][28];
    ele[32][24] != ele[35][29];
    ele[32][25] != ele[32][26];
    ele[32][25] != ele[32][27];
    ele[32][25] != ele[32][28];
    ele[32][25] != ele[32][29];
    ele[32][25] != ele[32][30];
    ele[32][25] != ele[32][31];
    ele[32][25] != ele[32][32];
    ele[32][25] != ele[32][33];
    ele[32][25] != ele[32][34];
    ele[32][25] != ele[32][35];
    ele[32][25] != ele[33][24];
    ele[32][25] != ele[33][25];
    ele[32][25] != ele[33][26];
    ele[32][25] != ele[33][27];
    ele[32][25] != ele[33][28];
    ele[32][25] != ele[33][29];
    ele[32][25] != ele[34][24];
    ele[32][25] != ele[34][25];
    ele[32][25] != ele[34][26];
    ele[32][25] != ele[34][27];
    ele[32][25] != ele[34][28];
    ele[32][25] != ele[34][29];
    ele[32][25] != ele[35][24];
    ele[32][25] != ele[35][25];
    ele[32][25] != ele[35][26];
    ele[32][25] != ele[35][27];
    ele[32][25] != ele[35][28];
    ele[32][25] != ele[35][29];
    ele[32][26] != ele[32][27];
    ele[32][26] != ele[32][28];
    ele[32][26] != ele[32][29];
    ele[32][26] != ele[32][30];
    ele[32][26] != ele[32][31];
    ele[32][26] != ele[32][32];
    ele[32][26] != ele[32][33];
    ele[32][26] != ele[32][34];
    ele[32][26] != ele[32][35];
    ele[32][26] != ele[33][24];
    ele[32][26] != ele[33][25];
    ele[32][26] != ele[33][26];
    ele[32][26] != ele[33][27];
    ele[32][26] != ele[33][28];
    ele[32][26] != ele[33][29];
    ele[32][26] != ele[34][24];
    ele[32][26] != ele[34][25];
    ele[32][26] != ele[34][26];
    ele[32][26] != ele[34][27];
    ele[32][26] != ele[34][28];
    ele[32][26] != ele[34][29];
    ele[32][26] != ele[35][24];
    ele[32][26] != ele[35][25];
    ele[32][26] != ele[35][26];
    ele[32][26] != ele[35][27];
    ele[32][26] != ele[35][28];
    ele[32][26] != ele[35][29];
    ele[32][27] != ele[32][28];
    ele[32][27] != ele[32][29];
    ele[32][27] != ele[32][30];
    ele[32][27] != ele[32][31];
    ele[32][27] != ele[32][32];
    ele[32][27] != ele[32][33];
    ele[32][27] != ele[32][34];
    ele[32][27] != ele[32][35];
    ele[32][27] != ele[33][24];
    ele[32][27] != ele[33][25];
    ele[32][27] != ele[33][26];
    ele[32][27] != ele[33][27];
    ele[32][27] != ele[33][28];
    ele[32][27] != ele[33][29];
    ele[32][27] != ele[34][24];
    ele[32][27] != ele[34][25];
    ele[32][27] != ele[34][26];
    ele[32][27] != ele[34][27];
    ele[32][27] != ele[34][28];
    ele[32][27] != ele[34][29];
    ele[32][27] != ele[35][24];
    ele[32][27] != ele[35][25];
    ele[32][27] != ele[35][26];
    ele[32][27] != ele[35][27];
    ele[32][27] != ele[35][28];
    ele[32][27] != ele[35][29];
    ele[32][28] != ele[32][29];
    ele[32][28] != ele[32][30];
    ele[32][28] != ele[32][31];
    ele[32][28] != ele[32][32];
    ele[32][28] != ele[32][33];
    ele[32][28] != ele[32][34];
    ele[32][28] != ele[32][35];
    ele[32][28] != ele[33][24];
    ele[32][28] != ele[33][25];
    ele[32][28] != ele[33][26];
    ele[32][28] != ele[33][27];
    ele[32][28] != ele[33][28];
    ele[32][28] != ele[33][29];
    ele[32][28] != ele[34][24];
    ele[32][28] != ele[34][25];
    ele[32][28] != ele[34][26];
    ele[32][28] != ele[34][27];
    ele[32][28] != ele[34][28];
    ele[32][28] != ele[34][29];
    ele[32][28] != ele[35][24];
    ele[32][28] != ele[35][25];
    ele[32][28] != ele[35][26];
    ele[32][28] != ele[35][27];
    ele[32][28] != ele[35][28];
    ele[32][28] != ele[35][29];
    ele[32][29] != ele[32][30];
    ele[32][29] != ele[32][31];
    ele[32][29] != ele[32][32];
    ele[32][29] != ele[32][33];
    ele[32][29] != ele[32][34];
    ele[32][29] != ele[32][35];
    ele[32][29] != ele[33][24];
    ele[32][29] != ele[33][25];
    ele[32][29] != ele[33][26];
    ele[32][29] != ele[33][27];
    ele[32][29] != ele[33][28];
    ele[32][29] != ele[33][29];
    ele[32][29] != ele[34][24];
    ele[32][29] != ele[34][25];
    ele[32][29] != ele[34][26];
    ele[32][29] != ele[34][27];
    ele[32][29] != ele[34][28];
    ele[32][29] != ele[34][29];
    ele[32][29] != ele[35][24];
    ele[32][29] != ele[35][25];
    ele[32][29] != ele[35][26];
    ele[32][29] != ele[35][27];
    ele[32][29] != ele[35][28];
    ele[32][29] != ele[35][29];
    ele[32][3] != ele[32][10];
    ele[32][3] != ele[32][11];
    ele[32][3] != ele[32][12];
    ele[32][3] != ele[32][13];
    ele[32][3] != ele[32][14];
    ele[32][3] != ele[32][15];
    ele[32][3] != ele[32][16];
    ele[32][3] != ele[32][17];
    ele[32][3] != ele[32][18];
    ele[32][3] != ele[32][19];
    ele[32][3] != ele[32][20];
    ele[32][3] != ele[32][21];
    ele[32][3] != ele[32][22];
    ele[32][3] != ele[32][23];
    ele[32][3] != ele[32][24];
    ele[32][3] != ele[32][25];
    ele[32][3] != ele[32][26];
    ele[32][3] != ele[32][27];
    ele[32][3] != ele[32][28];
    ele[32][3] != ele[32][29];
    ele[32][3] != ele[32][30];
    ele[32][3] != ele[32][31];
    ele[32][3] != ele[32][32];
    ele[32][3] != ele[32][33];
    ele[32][3] != ele[32][34];
    ele[32][3] != ele[32][35];
    ele[32][3] != ele[32][4];
    ele[32][3] != ele[32][5];
    ele[32][3] != ele[32][6];
    ele[32][3] != ele[32][7];
    ele[32][3] != ele[32][8];
    ele[32][3] != ele[32][9];
    ele[32][3] != ele[33][0];
    ele[32][3] != ele[33][1];
    ele[32][3] != ele[33][2];
    ele[32][3] != ele[33][3];
    ele[32][3] != ele[33][4];
    ele[32][3] != ele[33][5];
    ele[32][3] != ele[34][0];
    ele[32][3] != ele[34][1];
    ele[32][3] != ele[34][2];
    ele[32][3] != ele[34][3];
    ele[32][3] != ele[34][4];
    ele[32][3] != ele[34][5];
    ele[32][3] != ele[35][0];
    ele[32][3] != ele[35][1];
    ele[32][3] != ele[35][2];
    ele[32][3] != ele[35][3];
    ele[32][3] != ele[35][4];
    ele[32][3] != ele[35][5];
    ele[32][30] != ele[32][31];
    ele[32][30] != ele[32][32];
    ele[32][30] != ele[32][33];
    ele[32][30] != ele[32][34];
    ele[32][30] != ele[32][35];
    ele[32][30] != ele[33][30];
    ele[32][30] != ele[33][31];
    ele[32][30] != ele[33][32];
    ele[32][30] != ele[33][33];
    ele[32][30] != ele[33][34];
    ele[32][30] != ele[33][35];
    ele[32][30] != ele[34][30];
    ele[32][30] != ele[34][31];
    ele[32][30] != ele[34][32];
    ele[32][30] != ele[34][33];
    ele[32][30] != ele[34][34];
    ele[32][30] != ele[34][35];
    ele[32][30] != ele[35][30];
    ele[32][30] != ele[35][31];
    ele[32][30] != ele[35][32];
    ele[32][30] != ele[35][33];
    ele[32][30] != ele[35][34];
    ele[32][30] != ele[35][35];
    ele[32][31] != ele[32][32];
    ele[32][31] != ele[32][33];
    ele[32][31] != ele[32][34];
    ele[32][31] != ele[32][35];
    ele[32][31] != ele[33][30];
    ele[32][31] != ele[33][31];
    ele[32][31] != ele[33][32];
    ele[32][31] != ele[33][33];
    ele[32][31] != ele[33][34];
    ele[32][31] != ele[33][35];
    ele[32][31] != ele[34][30];
    ele[32][31] != ele[34][31];
    ele[32][31] != ele[34][32];
    ele[32][31] != ele[34][33];
    ele[32][31] != ele[34][34];
    ele[32][31] != ele[34][35];
    ele[32][31] != ele[35][30];
    ele[32][31] != ele[35][31];
    ele[32][31] != ele[35][32];
    ele[32][31] != ele[35][33];
    ele[32][31] != ele[35][34];
    ele[32][31] != ele[35][35];
    ele[32][32] != ele[32][33];
    ele[32][32] != ele[32][34];
    ele[32][32] != ele[32][35];
    ele[32][32] != ele[33][30];
    ele[32][32] != ele[33][31];
    ele[32][32] != ele[33][32];
    ele[32][32] != ele[33][33];
    ele[32][32] != ele[33][34];
    ele[32][32] != ele[33][35];
    ele[32][32] != ele[34][30];
    ele[32][32] != ele[34][31];
    ele[32][32] != ele[34][32];
    ele[32][32] != ele[34][33];
    ele[32][32] != ele[34][34];
    ele[32][32] != ele[34][35];
    ele[32][32] != ele[35][30];
    ele[32][32] != ele[35][31];
    ele[32][32] != ele[35][32];
    ele[32][32] != ele[35][33];
    ele[32][32] != ele[35][34];
    ele[32][32] != ele[35][35];
    ele[32][33] != ele[32][34];
    ele[32][33] != ele[32][35];
    ele[32][33] != ele[33][30];
    ele[32][33] != ele[33][31];
    ele[32][33] != ele[33][32];
    ele[32][33] != ele[33][33];
    ele[32][33] != ele[33][34];
    ele[32][33] != ele[33][35];
    ele[32][33] != ele[34][30];
    ele[32][33] != ele[34][31];
    ele[32][33] != ele[34][32];
    ele[32][33] != ele[34][33];
    ele[32][33] != ele[34][34];
    ele[32][33] != ele[34][35];
    ele[32][33] != ele[35][30];
    ele[32][33] != ele[35][31];
    ele[32][33] != ele[35][32];
    ele[32][33] != ele[35][33];
    ele[32][33] != ele[35][34];
    ele[32][33] != ele[35][35];
    ele[32][34] != ele[32][35];
    ele[32][34] != ele[33][30];
    ele[32][34] != ele[33][31];
    ele[32][34] != ele[33][32];
    ele[32][34] != ele[33][33];
    ele[32][34] != ele[33][34];
    ele[32][34] != ele[33][35];
    ele[32][34] != ele[34][30];
    ele[32][34] != ele[34][31];
    ele[32][34] != ele[34][32];
    ele[32][34] != ele[34][33];
    ele[32][34] != ele[34][34];
    ele[32][34] != ele[34][35];
    ele[32][34] != ele[35][30];
    ele[32][34] != ele[35][31];
    ele[32][34] != ele[35][32];
    ele[32][34] != ele[35][33];
    ele[32][34] != ele[35][34];
    ele[32][34] != ele[35][35];
    ele[32][35] != ele[33][30];
    ele[32][35] != ele[33][31];
    ele[32][35] != ele[33][32];
    ele[32][35] != ele[33][33];
    ele[32][35] != ele[33][34];
    ele[32][35] != ele[33][35];
    ele[32][35] != ele[34][30];
    ele[32][35] != ele[34][31];
    ele[32][35] != ele[34][32];
    ele[32][35] != ele[34][33];
    ele[32][35] != ele[34][34];
    ele[32][35] != ele[34][35];
    ele[32][35] != ele[35][30];
    ele[32][35] != ele[35][31];
    ele[32][35] != ele[35][32];
    ele[32][35] != ele[35][33];
    ele[32][35] != ele[35][34];
    ele[32][35] != ele[35][35];
    ele[32][4] != ele[32][10];
    ele[32][4] != ele[32][11];
    ele[32][4] != ele[32][12];
    ele[32][4] != ele[32][13];
    ele[32][4] != ele[32][14];
    ele[32][4] != ele[32][15];
    ele[32][4] != ele[32][16];
    ele[32][4] != ele[32][17];
    ele[32][4] != ele[32][18];
    ele[32][4] != ele[32][19];
    ele[32][4] != ele[32][20];
    ele[32][4] != ele[32][21];
    ele[32][4] != ele[32][22];
    ele[32][4] != ele[32][23];
    ele[32][4] != ele[32][24];
    ele[32][4] != ele[32][25];
    ele[32][4] != ele[32][26];
    ele[32][4] != ele[32][27];
    ele[32][4] != ele[32][28];
    ele[32][4] != ele[32][29];
    ele[32][4] != ele[32][30];
    ele[32][4] != ele[32][31];
    ele[32][4] != ele[32][32];
    ele[32][4] != ele[32][33];
    ele[32][4] != ele[32][34];
    ele[32][4] != ele[32][35];
    ele[32][4] != ele[32][5];
    ele[32][4] != ele[32][6];
    ele[32][4] != ele[32][7];
    ele[32][4] != ele[32][8];
    ele[32][4] != ele[32][9];
    ele[32][4] != ele[33][0];
    ele[32][4] != ele[33][1];
    ele[32][4] != ele[33][2];
    ele[32][4] != ele[33][3];
    ele[32][4] != ele[33][4];
    ele[32][4] != ele[33][5];
    ele[32][4] != ele[34][0];
    ele[32][4] != ele[34][1];
    ele[32][4] != ele[34][2];
    ele[32][4] != ele[34][3];
    ele[32][4] != ele[34][4];
    ele[32][4] != ele[34][5];
    ele[32][4] != ele[35][0];
    ele[32][4] != ele[35][1];
    ele[32][4] != ele[35][2];
    ele[32][4] != ele[35][3];
    ele[32][4] != ele[35][4];
    ele[32][4] != ele[35][5];
    ele[32][5] != ele[32][10];
    ele[32][5] != ele[32][11];
    ele[32][5] != ele[32][12];
    ele[32][5] != ele[32][13];
    ele[32][5] != ele[32][14];
    ele[32][5] != ele[32][15];
    ele[32][5] != ele[32][16];
    ele[32][5] != ele[32][17];
    ele[32][5] != ele[32][18];
    ele[32][5] != ele[32][19];
    ele[32][5] != ele[32][20];
    ele[32][5] != ele[32][21];
    ele[32][5] != ele[32][22];
    ele[32][5] != ele[32][23];
    ele[32][5] != ele[32][24];
    ele[32][5] != ele[32][25];
    ele[32][5] != ele[32][26];
    ele[32][5] != ele[32][27];
    ele[32][5] != ele[32][28];
    ele[32][5] != ele[32][29];
    ele[32][5] != ele[32][30];
    ele[32][5] != ele[32][31];
    ele[32][5] != ele[32][32];
    ele[32][5] != ele[32][33];
    ele[32][5] != ele[32][34];
    ele[32][5] != ele[32][35];
    ele[32][5] != ele[32][6];
    ele[32][5] != ele[32][7];
    ele[32][5] != ele[32][8];
    ele[32][5] != ele[32][9];
    ele[32][5] != ele[33][0];
    ele[32][5] != ele[33][1];
    ele[32][5] != ele[33][2];
    ele[32][5] != ele[33][3];
    ele[32][5] != ele[33][4];
    ele[32][5] != ele[33][5];
    ele[32][5] != ele[34][0];
    ele[32][5] != ele[34][1];
    ele[32][5] != ele[34][2];
    ele[32][5] != ele[34][3];
    ele[32][5] != ele[34][4];
    ele[32][5] != ele[34][5];
    ele[32][5] != ele[35][0];
    ele[32][5] != ele[35][1];
    ele[32][5] != ele[35][2];
    ele[32][5] != ele[35][3];
    ele[32][5] != ele[35][4];
    ele[32][5] != ele[35][5];
    ele[32][6] != ele[32][10];
    ele[32][6] != ele[32][11];
    ele[32][6] != ele[32][12];
    ele[32][6] != ele[32][13];
    ele[32][6] != ele[32][14];
    ele[32][6] != ele[32][15];
    ele[32][6] != ele[32][16];
    ele[32][6] != ele[32][17];
    ele[32][6] != ele[32][18];
    ele[32][6] != ele[32][19];
    ele[32][6] != ele[32][20];
    ele[32][6] != ele[32][21];
    ele[32][6] != ele[32][22];
    ele[32][6] != ele[32][23];
    ele[32][6] != ele[32][24];
    ele[32][6] != ele[32][25];
    ele[32][6] != ele[32][26];
    ele[32][6] != ele[32][27];
    ele[32][6] != ele[32][28];
    ele[32][6] != ele[32][29];
    ele[32][6] != ele[32][30];
    ele[32][6] != ele[32][31];
    ele[32][6] != ele[32][32];
    ele[32][6] != ele[32][33];
    ele[32][6] != ele[32][34];
    ele[32][6] != ele[32][35];
    ele[32][6] != ele[32][7];
    ele[32][6] != ele[32][8];
    ele[32][6] != ele[32][9];
    ele[32][6] != ele[33][10];
    ele[32][6] != ele[33][11];
    ele[32][6] != ele[33][6];
    ele[32][6] != ele[33][7];
    ele[32][6] != ele[33][8];
    ele[32][6] != ele[33][9];
    ele[32][6] != ele[34][10];
    ele[32][6] != ele[34][11];
    ele[32][6] != ele[34][6];
    ele[32][6] != ele[34][7];
    ele[32][6] != ele[34][8];
    ele[32][6] != ele[34][9];
    ele[32][6] != ele[35][10];
    ele[32][6] != ele[35][11];
    ele[32][6] != ele[35][6];
    ele[32][6] != ele[35][7];
    ele[32][6] != ele[35][8];
    ele[32][6] != ele[35][9];
    ele[32][7] != ele[32][10];
    ele[32][7] != ele[32][11];
    ele[32][7] != ele[32][12];
    ele[32][7] != ele[32][13];
    ele[32][7] != ele[32][14];
    ele[32][7] != ele[32][15];
    ele[32][7] != ele[32][16];
    ele[32][7] != ele[32][17];
    ele[32][7] != ele[32][18];
    ele[32][7] != ele[32][19];
    ele[32][7] != ele[32][20];
    ele[32][7] != ele[32][21];
    ele[32][7] != ele[32][22];
    ele[32][7] != ele[32][23];
    ele[32][7] != ele[32][24];
    ele[32][7] != ele[32][25];
    ele[32][7] != ele[32][26];
    ele[32][7] != ele[32][27];
    ele[32][7] != ele[32][28];
    ele[32][7] != ele[32][29];
    ele[32][7] != ele[32][30];
    ele[32][7] != ele[32][31];
    ele[32][7] != ele[32][32];
    ele[32][7] != ele[32][33];
    ele[32][7] != ele[32][34];
    ele[32][7] != ele[32][35];
    ele[32][7] != ele[32][8];
    ele[32][7] != ele[32][9];
    ele[32][7] != ele[33][10];
    ele[32][7] != ele[33][11];
    ele[32][7] != ele[33][6];
    ele[32][7] != ele[33][7];
    ele[32][7] != ele[33][8];
    ele[32][7] != ele[33][9];
    ele[32][7] != ele[34][10];
    ele[32][7] != ele[34][11];
    ele[32][7] != ele[34][6];
    ele[32][7] != ele[34][7];
    ele[32][7] != ele[34][8];
    ele[32][7] != ele[34][9];
    ele[32][7] != ele[35][10];
    ele[32][7] != ele[35][11];
    ele[32][7] != ele[35][6];
    ele[32][7] != ele[35][7];
    ele[32][7] != ele[35][8];
    ele[32][7] != ele[35][9];
    ele[32][8] != ele[32][10];
    ele[32][8] != ele[32][11];
    ele[32][8] != ele[32][12];
    ele[32][8] != ele[32][13];
    ele[32][8] != ele[32][14];
    ele[32][8] != ele[32][15];
    ele[32][8] != ele[32][16];
    ele[32][8] != ele[32][17];
    ele[32][8] != ele[32][18];
    ele[32][8] != ele[32][19];
    ele[32][8] != ele[32][20];
    ele[32][8] != ele[32][21];
    ele[32][8] != ele[32][22];
    ele[32][8] != ele[32][23];
    ele[32][8] != ele[32][24];
    ele[32][8] != ele[32][25];
    ele[32][8] != ele[32][26];
    ele[32][8] != ele[32][27];
    ele[32][8] != ele[32][28];
    ele[32][8] != ele[32][29];
    ele[32][8] != ele[32][30];
    ele[32][8] != ele[32][31];
    ele[32][8] != ele[32][32];
    ele[32][8] != ele[32][33];
    ele[32][8] != ele[32][34];
    ele[32][8] != ele[32][35];
    ele[32][8] != ele[32][9];
    ele[32][8] != ele[33][10];
    ele[32][8] != ele[33][11];
    ele[32][8] != ele[33][6];
    ele[32][8] != ele[33][7];
    ele[32][8] != ele[33][8];
    ele[32][8] != ele[33][9];
    ele[32][8] != ele[34][10];
    ele[32][8] != ele[34][11];
    ele[32][8] != ele[34][6];
    ele[32][8] != ele[34][7];
    ele[32][8] != ele[34][8];
    ele[32][8] != ele[34][9];
    ele[32][8] != ele[35][10];
    ele[32][8] != ele[35][11];
    ele[32][8] != ele[35][6];
    ele[32][8] != ele[35][7];
    ele[32][8] != ele[35][8];
    ele[32][8] != ele[35][9];
    ele[32][9] != ele[32][10];
    ele[32][9] != ele[32][11];
    ele[32][9] != ele[32][12];
    ele[32][9] != ele[32][13];
    ele[32][9] != ele[32][14];
    ele[32][9] != ele[32][15];
    ele[32][9] != ele[32][16];
    ele[32][9] != ele[32][17];
    ele[32][9] != ele[32][18];
    ele[32][9] != ele[32][19];
    ele[32][9] != ele[32][20];
    ele[32][9] != ele[32][21];
    ele[32][9] != ele[32][22];
    ele[32][9] != ele[32][23];
    ele[32][9] != ele[32][24];
    ele[32][9] != ele[32][25];
    ele[32][9] != ele[32][26];
    ele[32][9] != ele[32][27];
    ele[32][9] != ele[32][28];
    ele[32][9] != ele[32][29];
    ele[32][9] != ele[32][30];
    ele[32][9] != ele[32][31];
    ele[32][9] != ele[32][32];
    ele[32][9] != ele[32][33];
    ele[32][9] != ele[32][34];
    ele[32][9] != ele[32][35];
    ele[32][9] != ele[33][10];
    ele[32][9] != ele[33][11];
    ele[32][9] != ele[33][6];
    ele[32][9] != ele[33][7];
    ele[32][9] != ele[33][8];
    ele[32][9] != ele[33][9];
    ele[32][9] != ele[34][10];
    ele[32][9] != ele[34][11];
    ele[32][9] != ele[34][6];
    ele[32][9] != ele[34][7];
    ele[32][9] != ele[34][8];
    ele[32][9] != ele[34][9];
    ele[32][9] != ele[35][10];
    ele[32][9] != ele[35][11];
    ele[32][9] != ele[35][6];
    ele[32][9] != ele[35][7];
    ele[32][9] != ele[35][8];
    ele[32][9] != ele[35][9];
    ele[33][0] != ele[33][1];
    ele[33][0] != ele[33][10];
    ele[33][0] != ele[33][11];
    ele[33][0] != ele[33][12];
    ele[33][0] != ele[33][13];
    ele[33][0] != ele[33][14];
    ele[33][0] != ele[33][15];
    ele[33][0] != ele[33][16];
    ele[33][0] != ele[33][17];
    ele[33][0] != ele[33][18];
    ele[33][0] != ele[33][19];
    ele[33][0] != ele[33][2];
    ele[33][0] != ele[33][20];
    ele[33][0] != ele[33][21];
    ele[33][0] != ele[33][22];
    ele[33][0] != ele[33][23];
    ele[33][0] != ele[33][24];
    ele[33][0] != ele[33][25];
    ele[33][0] != ele[33][26];
    ele[33][0] != ele[33][27];
    ele[33][0] != ele[33][28];
    ele[33][0] != ele[33][29];
    ele[33][0] != ele[33][3];
    ele[33][0] != ele[33][30];
    ele[33][0] != ele[33][31];
    ele[33][0] != ele[33][32];
    ele[33][0] != ele[33][33];
    ele[33][0] != ele[33][34];
    ele[33][0] != ele[33][35];
    ele[33][0] != ele[33][4];
    ele[33][0] != ele[33][5];
    ele[33][0] != ele[33][6];
    ele[33][0] != ele[33][7];
    ele[33][0] != ele[33][8];
    ele[33][0] != ele[33][9];
    ele[33][0] != ele[34][0];
    ele[33][0] != ele[34][1];
    ele[33][0] != ele[34][2];
    ele[33][0] != ele[34][3];
    ele[33][0] != ele[34][4];
    ele[33][0] != ele[34][5];
    ele[33][0] != ele[35][0];
    ele[33][0] != ele[35][1];
    ele[33][0] != ele[35][2];
    ele[33][0] != ele[35][3];
    ele[33][0] != ele[35][4];
    ele[33][0] != ele[35][5];
    ele[33][1] != ele[33][10];
    ele[33][1] != ele[33][11];
    ele[33][1] != ele[33][12];
    ele[33][1] != ele[33][13];
    ele[33][1] != ele[33][14];
    ele[33][1] != ele[33][15];
    ele[33][1] != ele[33][16];
    ele[33][1] != ele[33][17];
    ele[33][1] != ele[33][18];
    ele[33][1] != ele[33][19];
    ele[33][1] != ele[33][2];
    ele[33][1] != ele[33][20];
    ele[33][1] != ele[33][21];
    ele[33][1] != ele[33][22];
    ele[33][1] != ele[33][23];
    ele[33][1] != ele[33][24];
    ele[33][1] != ele[33][25];
    ele[33][1] != ele[33][26];
    ele[33][1] != ele[33][27];
    ele[33][1] != ele[33][28];
    ele[33][1] != ele[33][29];
    ele[33][1] != ele[33][3];
    ele[33][1] != ele[33][30];
    ele[33][1] != ele[33][31];
    ele[33][1] != ele[33][32];
    ele[33][1] != ele[33][33];
    ele[33][1] != ele[33][34];
    ele[33][1] != ele[33][35];
    ele[33][1] != ele[33][4];
    ele[33][1] != ele[33][5];
    ele[33][1] != ele[33][6];
    ele[33][1] != ele[33][7];
    ele[33][1] != ele[33][8];
    ele[33][1] != ele[33][9];
    ele[33][1] != ele[34][0];
    ele[33][1] != ele[34][1];
    ele[33][1] != ele[34][2];
    ele[33][1] != ele[34][3];
    ele[33][1] != ele[34][4];
    ele[33][1] != ele[34][5];
    ele[33][1] != ele[35][0];
    ele[33][1] != ele[35][1];
    ele[33][1] != ele[35][2];
    ele[33][1] != ele[35][3];
    ele[33][1] != ele[35][4];
    ele[33][1] != ele[35][5];
    ele[33][10] != ele[33][11];
    ele[33][10] != ele[33][12];
    ele[33][10] != ele[33][13];
    ele[33][10] != ele[33][14];
    ele[33][10] != ele[33][15];
    ele[33][10] != ele[33][16];
    ele[33][10] != ele[33][17];
    ele[33][10] != ele[33][18];
    ele[33][10] != ele[33][19];
    ele[33][10] != ele[33][20];
    ele[33][10] != ele[33][21];
    ele[33][10] != ele[33][22];
    ele[33][10] != ele[33][23];
    ele[33][10] != ele[33][24];
    ele[33][10] != ele[33][25];
    ele[33][10] != ele[33][26];
    ele[33][10] != ele[33][27];
    ele[33][10] != ele[33][28];
    ele[33][10] != ele[33][29];
    ele[33][10] != ele[33][30];
    ele[33][10] != ele[33][31];
    ele[33][10] != ele[33][32];
    ele[33][10] != ele[33][33];
    ele[33][10] != ele[33][34];
    ele[33][10] != ele[33][35];
    ele[33][10] != ele[34][10];
    ele[33][10] != ele[34][11];
    ele[33][10] != ele[34][6];
    ele[33][10] != ele[34][7];
    ele[33][10] != ele[34][8];
    ele[33][10] != ele[34][9];
    ele[33][10] != ele[35][10];
    ele[33][10] != ele[35][11];
    ele[33][10] != ele[35][6];
    ele[33][10] != ele[35][7];
    ele[33][10] != ele[35][8];
    ele[33][10] != ele[35][9];
    ele[33][11] != ele[33][12];
    ele[33][11] != ele[33][13];
    ele[33][11] != ele[33][14];
    ele[33][11] != ele[33][15];
    ele[33][11] != ele[33][16];
    ele[33][11] != ele[33][17];
    ele[33][11] != ele[33][18];
    ele[33][11] != ele[33][19];
    ele[33][11] != ele[33][20];
    ele[33][11] != ele[33][21];
    ele[33][11] != ele[33][22];
    ele[33][11] != ele[33][23];
    ele[33][11] != ele[33][24];
    ele[33][11] != ele[33][25];
    ele[33][11] != ele[33][26];
    ele[33][11] != ele[33][27];
    ele[33][11] != ele[33][28];
    ele[33][11] != ele[33][29];
    ele[33][11] != ele[33][30];
    ele[33][11] != ele[33][31];
    ele[33][11] != ele[33][32];
    ele[33][11] != ele[33][33];
    ele[33][11] != ele[33][34];
    ele[33][11] != ele[33][35];
    ele[33][11] != ele[34][10];
    ele[33][11] != ele[34][11];
    ele[33][11] != ele[34][6];
    ele[33][11] != ele[34][7];
    ele[33][11] != ele[34][8];
    ele[33][11] != ele[34][9];
    ele[33][11] != ele[35][10];
    ele[33][11] != ele[35][11];
    ele[33][11] != ele[35][6];
    ele[33][11] != ele[35][7];
    ele[33][11] != ele[35][8];
    ele[33][11] != ele[35][9];
    ele[33][12] != ele[33][13];
    ele[33][12] != ele[33][14];
    ele[33][12] != ele[33][15];
    ele[33][12] != ele[33][16];
    ele[33][12] != ele[33][17];
    ele[33][12] != ele[33][18];
    ele[33][12] != ele[33][19];
    ele[33][12] != ele[33][20];
    ele[33][12] != ele[33][21];
    ele[33][12] != ele[33][22];
    ele[33][12] != ele[33][23];
    ele[33][12] != ele[33][24];
    ele[33][12] != ele[33][25];
    ele[33][12] != ele[33][26];
    ele[33][12] != ele[33][27];
    ele[33][12] != ele[33][28];
    ele[33][12] != ele[33][29];
    ele[33][12] != ele[33][30];
    ele[33][12] != ele[33][31];
    ele[33][12] != ele[33][32];
    ele[33][12] != ele[33][33];
    ele[33][12] != ele[33][34];
    ele[33][12] != ele[33][35];
    ele[33][12] != ele[34][12];
    ele[33][12] != ele[34][13];
    ele[33][12] != ele[34][14];
    ele[33][12] != ele[34][15];
    ele[33][12] != ele[34][16];
    ele[33][12] != ele[34][17];
    ele[33][12] != ele[35][12];
    ele[33][12] != ele[35][13];
    ele[33][12] != ele[35][14];
    ele[33][12] != ele[35][15];
    ele[33][12] != ele[35][16];
    ele[33][12] != ele[35][17];
    ele[33][13] != ele[33][14];
    ele[33][13] != ele[33][15];
    ele[33][13] != ele[33][16];
    ele[33][13] != ele[33][17];
    ele[33][13] != ele[33][18];
    ele[33][13] != ele[33][19];
    ele[33][13] != ele[33][20];
    ele[33][13] != ele[33][21];
    ele[33][13] != ele[33][22];
    ele[33][13] != ele[33][23];
    ele[33][13] != ele[33][24];
    ele[33][13] != ele[33][25];
    ele[33][13] != ele[33][26];
    ele[33][13] != ele[33][27];
    ele[33][13] != ele[33][28];
    ele[33][13] != ele[33][29];
    ele[33][13] != ele[33][30];
    ele[33][13] != ele[33][31];
    ele[33][13] != ele[33][32];
    ele[33][13] != ele[33][33];
    ele[33][13] != ele[33][34];
    ele[33][13] != ele[33][35];
    ele[33][13] != ele[34][12];
    ele[33][13] != ele[34][13];
    ele[33][13] != ele[34][14];
    ele[33][13] != ele[34][15];
    ele[33][13] != ele[34][16];
    ele[33][13] != ele[34][17];
    ele[33][13] != ele[35][12];
    ele[33][13] != ele[35][13];
    ele[33][13] != ele[35][14];
    ele[33][13] != ele[35][15];
    ele[33][13] != ele[35][16];
    ele[33][13] != ele[35][17];
    ele[33][14] != ele[33][15];
    ele[33][14] != ele[33][16];
    ele[33][14] != ele[33][17];
    ele[33][14] != ele[33][18];
    ele[33][14] != ele[33][19];
    ele[33][14] != ele[33][20];
    ele[33][14] != ele[33][21];
    ele[33][14] != ele[33][22];
    ele[33][14] != ele[33][23];
    ele[33][14] != ele[33][24];
    ele[33][14] != ele[33][25];
    ele[33][14] != ele[33][26];
    ele[33][14] != ele[33][27];
    ele[33][14] != ele[33][28];
    ele[33][14] != ele[33][29];
    ele[33][14] != ele[33][30];
    ele[33][14] != ele[33][31];
    ele[33][14] != ele[33][32];
    ele[33][14] != ele[33][33];
    ele[33][14] != ele[33][34];
    ele[33][14] != ele[33][35];
    ele[33][14] != ele[34][12];
    ele[33][14] != ele[34][13];
    ele[33][14] != ele[34][14];
    ele[33][14] != ele[34][15];
    ele[33][14] != ele[34][16];
    ele[33][14] != ele[34][17];
    ele[33][14] != ele[35][12];
    ele[33][14] != ele[35][13];
    ele[33][14] != ele[35][14];
    ele[33][14] != ele[35][15];
    ele[33][14] != ele[35][16];
    ele[33][14] != ele[35][17];
    ele[33][15] != ele[33][16];
    ele[33][15] != ele[33][17];
    ele[33][15] != ele[33][18];
    ele[33][15] != ele[33][19];
    ele[33][15] != ele[33][20];
    ele[33][15] != ele[33][21];
    ele[33][15] != ele[33][22];
    ele[33][15] != ele[33][23];
    ele[33][15] != ele[33][24];
    ele[33][15] != ele[33][25];
    ele[33][15] != ele[33][26];
    ele[33][15] != ele[33][27];
    ele[33][15] != ele[33][28];
    ele[33][15] != ele[33][29];
    ele[33][15] != ele[33][30];
    ele[33][15] != ele[33][31];
    ele[33][15] != ele[33][32];
    ele[33][15] != ele[33][33];
    ele[33][15] != ele[33][34];
    ele[33][15] != ele[33][35];
    ele[33][15] != ele[34][12];
    ele[33][15] != ele[34][13];
    ele[33][15] != ele[34][14];
    ele[33][15] != ele[34][15];
    ele[33][15] != ele[34][16];
    ele[33][15] != ele[34][17];
    ele[33][15] != ele[35][12];
    ele[33][15] != ele[35][13];
    ele[33][15] != ele[35][14];
    ele[33][15] != ele[35][15];
    ele[33][15] != ele[35][16];
    ele[33][15] != ele[35][17];
    ele[33][16] != ele[33][17];
    ele[33][16] != ele[33][18];
    ele[33][16] != ele[33][19];
    ele[33][16] != ele[33][20];
    ele[33][16] != ele[33][21];
    ele[33][16] != ele[33][22];
    ele[33][16] != ele[33][23];
    ele[33][16] != ele[33][24];
    ele[33][16] != ele[33][25];
    ele[33][16] != ele[33][26];
    ele[33][16] != ele[33][27];
    ele[33][16] != ele[33][28];
    ele[33][16] != ele[33][29];
    ele[33][16] != ele[33][30];
    ele[33][16] != ele[33][31];
    ele[33][16] != ele[33][32];
    ele[33][16] != ele[33][33];
    ele[33][16] != ele[33][34];
    ele[33][16] != ele[33][35];
    ele[33][16] != ele[34][12];
    ele[33][16] != ele[34][13];
    ele[33][16] != ele[34][14];
    ele[33][16] != ele[34][15];
    ele[33][16] != ele[34][16];
    ele[33][16] != ele[34][17];
    ele[33][16] != ele[35][12];
    ele[33][16] != ele[35][13];
    ele[33][16] != ele[35][14];
    ele[33][16] != ele[35][15];
    ele[33][16] != ele[35][16];
    ele[33][16] != ele[35][17];
    ele[33][17] != ele[33][18];
    ele[33][17] != ele[33][19];
    ele[33][17] != ele[33][20];
    ele[33][17] != ele[33][21];
    ele[33][17] != ele[33][22];
    ele[33][17] != ele[33][23];
    ele[33][17] != ele[33][24];
    ele[33][17] != ele[33][25];
    ele[33][17] != ele[33][26];
    ele[33][17] != ele[33][27];
    ele[33][17] != ele[33][28];
    ele[33][17] != ele[33][29];
    ele[33][17] != ele[33][30];
    ele[33][17] != ele[33][31];
    ele[33][17] != ele[33][32];
    ele[33][17] != ele[33][33];
    ele[33][17] != ele[33][34];
    ele[33][17] != ele[33][35];
    ele[33][17] != ele[34][12];
    ele[33][17] != ele[34][13];
    ele[33][17] != ele[34][14];
    ele[33][17] != ele[34][15];
    ele[33][17] != ele[34][16];
    ele[33][17] != ele[34][17];
    ele[33][17] != ele[35][12];
    ele[33][17] != ele[35][13];
    ele[33][17] != ele[35][14];
    ele[33][17] != ele[35][15];
    ele[33][17] != ele[35][16];
    ele[33][17] != ele[35][17];
    ele[33][18] != ele[33][19];
    ele[33][18] != ele[33][20];
    ele[33][18] != ele[33][21];
    ele[33][18] != ele[33][22];
    ele[33][18] != ele[33][23];
    ele[33][18] != ele[33][24];
    ele[33][18] != ele[33][25];
    ele[33][18] != ele[33][26];
    ele[33][18] != ele[33][27];
    ele[33][18] != ele[33][28];
    ele[33][18] != ele[33][29];
    ele[33][18] != ele[33][30];
    ele[33][18] != ele[33][31];
    ele[33][18] != ele[33][32];
    ele[33][18] != ele[33][33];
    ele[33][18] != ele[33][34];
    ele[33][18] != ele[33][35];
    ele[33][18] != ele[34][18];
    ele[33][18] != ele[34][19];
    ele[33][18] != ele[34][20];
    ele[33][18] != ele[34][21];
    ele[33][18] != ele[34][22];
    ele[33][18] != ele[34][23];
    ele[33][18] != ele[35][18];
    ele[33][18] != ele[35][19];
    ele[33][18] != ele[35][20];
    ele[33][18] != ele[35][21];
    ele[33][18] != ele[35][22];
    ele[33][18] != ele[35][23];
    ele[33][19] != ele[33][20];
    ele[33][19] != ele[33][21];
    ele[33][19] != ele[33][22];
    ele[33][19] != ele[33][23];
    ele[33][19] != ele[33][24];
    ele[33][19] != ele[33][25];
    ele[33][19] != ele[33][26];
    ele[33][19] != ele[33][27];
    ele[33][19] != ele[33][28];
    ele[33][19] != ele[33][29];
    ele[33][19] != ele[33][30];
    ele[33][19] != ele[33][31];
    ele[33][19] != ele[33][32];
    ele[33][19] != ele[33][33];
    ele[33][19] != ele[33][34];
    ele[33][19] != ele[33][35];
    ele[33][19] != ele[34][18];
    ele[33][19] != ele[34][19];
    ele[33][19] != ele[34][20];
    ele[33][19] != ele[34][21];
    ele[33][19] != ele[34][22];
    ele[33][19] != ele[34][23];
    ele[33][19] != ele[35][18];
    ele[33][19] != ele[35][19];
    ele[33][19] != ele[35][20];
    ele[33][19] != ele[35][21];
    ele[33][19] != ele[35][22];
    ele[33][19] != ele[35][23];
    ele[33][2] != ele[33][10];
    ele[33][2] != ele[33][11];
    ele[33][2] != ele[33][12];
    ele[33][2] != ele[33][13];
    ele[33][2] != ele[33][14];
    ele[33][2] != ele[33][15];
    ele[33][2] != ele[33][16];
    ele[33][2] != ele[33][17];
    ele[33][2] != ele[33][18];
    ele[33][2] != ele[33][19];
    ele[33][2] != ele[33][20];
    ele[33][2] != ele[33][21];
    ele[33][2] != ele[33][22];
    ele[33][2] != ele[33][23];
    ele[33][2] != ele[33][24];
    ele[33][2] != ele[33][25];
    ele[33][2] != ele[33][26];
    ele[33][2] != ele[33][27];
    ele[33][2] != ele[33][28];
    ele[33][2] != ele[33][29];
    ele[33][2] != ele[33][3];
    ele[33][2] != ele[33][30];
    ele[33][2] != ele[33][31];
    ele[33][2] != ele[33][32];
    ele[33][2] != ele[33][33];
    ele[33][2] != ele[33][34];
    ele[33][2] != ele[33][35];
    ele[33][2] != ele[33][4];
    ele[33][2] != ele[33][5];
    ele[33][2] != ele[33][6];
    ele[33][2] != ele[33][7];
    ele[33][2] != ele[33][8];
    ele[33][2] != ele[33][9];
    ele[33][2] != ele[34][0];
    ele[33][2] != ele[34][1];
    ele[33][2] != ele[34][2];
    ele[33][2] != ele[34][3];
    ele[33][2] != ele[34][4];
    ele[33][2] != ele[34][5];
    ele[33][2] != ele[35][0];
    ele[33][2] != ele[35][1];
    ele[33][2] != ele[35][2];
    ele[33][2] != ele[35][3];
    ele[33][2] != ele[35][4];
    ele[33][2] != ele[35][5];
    ele[33][20] != ele[33][21];
    ele[33][20] != ele[33][22];
    ele[33][20] != ele[33][23];
    ele[33][20] != ele[33][24];
    ele[33][20] != ele[33][25];
    ele[33][20] != ele[33][26];
    ele[33][20] != ele[33][27];
    ele[33][20] != ele[33][28];
    ele[33][20] != ele[33][29];
    ele[33][20] != ele[33][30];
    ele[33][20] != ele[33][31];
    ele[33][20] != ele[33][32];
    ele[33][20] != ele[33][33];
    ele[33][20] != ele[33][34];
    ele[33][20] != ele[33][35];
    ele[33][20] != ele[34][18];
    ele[33][20] != ele[34][19];
    ele[33][20] != ele[34][20];
    ele[33][20] != ele[34][21];
    ele[33][20] != ele[34][22];
    ele[33][20] != ele[34][23];
    ele[33][20] != ele[35][18];
    ele[33][20] != ele[35][19];
    ele[33][20] != ele[35][20];
    ele[33][20] != ele[35][21];
    ele[33][20] != ele[35][22];
    ele[33][20] != ele[35][23];
    ele[33][21] != ele[33][22];
    ele[33][21] != ele[33][23];
    ele[33][21] != ele[33][24];
    ele[33][21] != ele[33][25];
    ele[33][21] != ele[33][26];
    ele[33][21] != ele[33][27];
    ele[33][21] != ele[33][28];
    ele[33][21] != ele[33][29];
    ele[33][21] != ele[33][30];
    ele[33][21] != ele[33][31];
    ele[33][21] != ele[33][32];
    ele[33][21] != ele[33][33];
    ele[33][21] != ele[33][34];
    ele[33][21] != ele[33][35];
    ele[33][21] != ele[34][18];
    ele[33][21] != ele[34][19];
    ele[33][21] != ele[34][20];
    ele[33][21] != ele[34][21];
    ele[33][21] != ele[34][22];
    ele[33][21] != ele[34][23];
    ele[33][21] != ele[35][18];
    ele[33][21] != ele[35][19];
    ele[33][21] != ele[35][20];
    ele[33][21] != ele[35][21];
    ele[33][21] != ele[35][22];
    ele[33][21] != ele[35][23];
    ele[33][22] != ele[33][23];
    ele[33][22] != ele[33][24];
    ele[33][22] != ele[33][25];
    ele[33][22] != ele[33][26];
    ele[33][22] != ele[33][27];
    ele[33][22] != ele[33][28];
    ele[33][22] != ele[33][29];
    ele[33][22] != ele[33][30];
    ele[33][22] != ele[33][31];
    ele[33][22] != ele[33][32];
    ele[33][22] != ele[33][33];
    ele[33][22] != ele[33][34];
    ele[33][22] != ele[33][35];
    ele[33][22] != ele[34][18];
    ele[33][22] != ele[34][19];
    ele[33][22] != ele[34][20];
    ele[33][22] != ele[34][21];
    ele[33][22] != ele[34][22];
    ele[33][22] != ele[34][23];
    ele[33][22] != ele[35][18];
    ele[33][22] != ele[35][19];
    ele[33][22] != ele[35][20];
    ele[33][22] != ele[35][21];
    ele[33][22] != ele[35][22];
    ele[33][22] != ele[35][23];
    ele[33][23] != ele[33][24];
    ele[33][23] != ele[33][25];
    ele[33][23] != ele[33][26];
    ele[33][23] != ele[33][27];
    ele[33][23] != ele[33][28];
    ele[33][23] != ele[33][29];
    ele[33][23] != ele[33][30];
    ele[33][23] != ele[33][31];
    ele[33][23] != ele[33][32];
    ele[33][23] != ele[33][33];
    ele[33][23] != ele[33][34];
    ele[33][23] != ele[33][35];
    ele[33][23] != ele[34][18];
    ele[33][23] != ele[34][19];
    ele[33][23] != ele[34][20];
    ele[33][23] != ele[34][21];
    ele[33][23] != ele[34][22];
    ele[33][23] != ele[34][23];
    ele[33][23] != ele[35][18];
    ele[33][23] != ele[35][19];
    ele[33][23] != ele[35][20];
    ele[33][23] != ele[35][21];
    ele[33][23] != ele[35][22];
    ele[33][23] != ele[35][23];
    ele[33][24] != ele[33][25];
    ele[33][24] != ele[33][26];
    ele[33][24] != ele[33][27];
    ele[33][24] != ele[33][28];
    ele[33][24] != ele[33][29];
    ele[33][24] != ele[33][30];
    ele[33][24] != ele[33][31];
    ele[33][24] != ele[33][32];
    ele[33][24] != ele[33][33];
    ele[33][24] != ele[33][34];
    ele[33][24] != ele[33][35];
    ele[33][24] != ele[34][24];
    ele[33][24] != ele[34][25];
    ele[33][24] != ele[34][26];
    ele[33][24] != ele[34][27];
    ele[33][24] != ele[34][28];
    ele[33][24] != ele[34][29];
    ele[33][24] != ele[35][24];
    ele[33][24] != ele[35][25];
    ele[33][24] != ele[35][26];
    ele[33][24] != ele[35][27];
    ele[33][24] != ele[35][28];
    ele[33][24] != ele[35][29];
    ele[33][25] != ele[33][26];
    ele[33][25] != ele[33][27];
    ele[33][25] != ele[33][28];
    ele[33][25] != ele[33][29];
    ele[33][25] != ele[33][30];
    ele[33][25] != ele[33][31];
    ele[33][25] != ele[33][32];
    ele[33][25] != ele[33][33];
    ele[33][25] != ele[33][34];
    ele[33][25] != ele[33][35];
    ele[33][25] != ele[34][24];
    ele[33][25] != ele[34][25];
    ele[33][25] != ele[34][26];
    ele[33][25] != ele[34][27];
    ele[33][25] != ele[34][28];
    ele[33][25] != ele[34][29];
    ele[33][25] != ele[35][24];
    ele[33][25] != ele[35][25];
    ele[33][25] != ele[35][26];
    ele[33][25] != ele[35][27];
    ele[33][25] != ele[35][28];
    ele[33][25] != ele[35][29];
    ele[33][26] != ele[33][27];
    ele[33][26] != ele[33][28];
    ele[33][26] != ele[33][29];
    ele[33][26] != ele[33][30];
    ele[33][26] != ele[33][31];
    ele[33][26] != ele[33][32];
    ele[33][26] != ele[33][33];
    ele[33][26] != ele[33][34];
    ele[33][26] != ele[33][35];
    ele[33][26] != ele[34][24];
    ele[33][26] != ele[34][25];
    ele[33][26] != ele[34][26];
    ele[33][26] != ele[34][27];
    ele[33][26] != ele[34][28];
    ele[33][26] != ele[34][29];
    ele[33][26] != ele[35][24];
    ele[33][26] != ele[35][25];
    ele[33][26] != ele[35][26];
    ele[33][26] != ele[35][27];
    ele[33][26] != ele[35][28];
    ele[33][26] != ele[35][29];
    ele[33][27] != ele[33][28];
    ele[33][27] != ele[33][29];
    ele[33][27] != ele[33][30];
    ele[33][27] != ele[33][31];
    ele[33][27] != ele[33][32];
    ele[33][27] != ele[33][33];
    ele[33][27] != ele[33][34];
    ele[33][27] != ele[33][35];
    ele[33][27] != ele[34][24];
    ele[33][27] != ele[34][25];
    ele[33][27] != ele[34][26];
    ele[33][27] != ele[34][27];
    ele[33][27] != ele[34][28];
    ele[33][27] != ele[34][29];
    ele[33][27] != ele[35][24];
    ele[33][27] != ele[35][25];
    ele[33][27] != ele[35][26];
    ele[33][27] != ele[35][27];
    ele[33][27] != ele[35][28];
    ele[33][27] != ele[35][29];
    ele[33][28] != ele[33][29];
    ele[33][28] != ele[33][30];
    ele[33][28] != ele[33][31];
    ele[33][28] != ele[33][32];
    ele[33][28] != ele[33][33];
    ele[33][28] != ele[33][34];
    ele[33][28] != ele[33][35];
    ele[33][28] != ele[34][24];
    ele[33][28] != ele[34][25];
    ele[33][28] != ele[34][26];
    ele[33][28] != ele[34][27];
    ele[33][28] != ele[34][28];
    ele[33][28] != ele[34][29];
    ele[33][28] != ele[35][24];
    ele[33][28] != ele[35][25];
    ele[33][28] != ele[35][26];
    ele[33][28] != ele[35][27];
    ele[33][28] != ele[35][28];
    ele[33][28] != ele[35][29];
    ele[33][29] != ele[33][30];
    ele[33][29] != ele[33][31];
    ele[33][29] != ele[33][32];
    ele[33][29] != ele[33][33];
    ele[33][29] != ele[33][34];
    ele[33][29] != ele[33][35];
    ele[33][29] != ele[34][24];
    ele[33][29] != ele[34][25];
    ele[33][29] != ele[34][26];
    ele[33][29] != ele[34][27];
    ele[33][29] != ele[34][28];
    ele[33][29] != ele[34][29];
    ele[33][29] != ele[35][24];
    ele[33][29] != ele[35][25];
    ele[33][29] != ele[35][26];
    ele[33][29] != ele[35][27];
    ele[33][29] != ele[35][28];
    ele[33][29] != ele[35][29];
    ele[33][3] != ele[33][10];
    ele[33][3] != ele[33][11];
    ele[33][3] != ele[33][12];
    ele[33][3] != ele[33][13];
    ele[33][3] != ele[33][14];
    ele[33][3] != ele[33][15];
    ele[33][3] != ele[33][16];
    ele[33][3] != ele[33][17];
    ele[33][3] != ele[33][18];
    ele[33][3] != ele[33][19];
    ele[33][3] != ele[33][20];
    ele[33][3] != ele[33][21];
    ele[33][3] != ele[33][22];
    ele[33][3] != ele[33][23];
    ele[33][3] != ele[33][24];
    ele[33][3] != ele[33][25];
    ele[33][3] != ele[33][26];
    ele[33][3] != ele[33][27];
    ele[33][3] != ele[33][28];
    ele[33][3] != ele[33][29];
    ele[33][3] != ele[33][30];
    ele[33][3] != ele[33][31];
    ele[33][3] != ele[33][32];
    ele[33][3] != ele[33][33];
    ele[33][3] != ele[33][34];
    ele[33][3] != ele[33][35];
    ele[33][3] != ele[33][4];
    ele[33][3] != ele[33][5];
    ele[33][3] != ele[33][6];
    ele[33][3] != ele[33][7];
    ele[33][3] != ele[33][8];
    ele[33][3] != ele[33][9];
    ele[33][3] != ele[34][0];
    ele[33][3] != ele[34][1];
    ele[33][3] != ele[34][2];
    ele[33][3] != ele[34][3];
    ele[33][3] != ele[34][4];
    ele[33][3] != ele[34][5];
    ele[33][3] != ele[35][0];
    ele[33][3] != ele[35][1];
    ele[33][3] != ele[35][2];
    ele[33][3] != ele[35][3];
    ele[33][3] != ele[35][4];
    ele[33][3] != ele[35][5];
    ele[33][30] != ele[33][31];
    ele[33][30] != ele[33][32];
    ele[33][30] != ele[33][33];
    ele[33][30] != ele[33][34];
    ele[33][30] != ele[33][35];
    ele[33][30] != ele[34][30];
    ele[33][30] != ele[34][31];
    ele[33][30] != ele[34][32];
    ele[33][30] != ele[34][33];
    ele[33][30] != ele[34][34];
    ele[33][30] != ele[34][35];
    ele[33][30] != ele[35][30];
    ele[33][30] != ele[35][31];
    ele[33][30] != ele[35][32];
    ele[33][30] != ele[35][33];
    ele[33][30] != ele[35][34];
    ele[33][30] != ele[35][35];
    ele[33][31] != ele[33][32];
    ele[33][31] != ele[33][33];
    ele[33][31] != ele[33][34];
    ele[33][31] != ele[33][35];
    ele[33][31] != ele[34][30];
    ele[33][31] != ele[34][31];
    ele[33][31] != ele[34][32];
    ele[33][31] != ele[34][33];
    ele[33][31] != ele[34][34];
    ele[33][31] != ele[34][35];
    ele[33][31] != ele[35][30];
    ele[33][31] != ele[35][31];
    ele[33][31] != ele[35][32];
    ele[33][31] != ele[35][33];
    ele[33][31] != ele[35][34];
    ele[33][31] != ele[35][35];
    ele[33][32] != ele[33][33];
    ele[33][32] != ele[33][34];
    ele[33][32] != ele[33][35];
    ele[33][32] != ele[34][30];
    ele[33][32] != ele[34][31];
    ele[33][32] != ele[34][32];
    ele[33][32] != ele[34][33];
    ele[33][32] != ele[34][34];
    ele[33][32] != ele[34][35];
    ele[33][32] != ele[35][30];
    ele[33][32] != ele[35][31];
    ele[33][32] != ele[35][32];
    ele[33][32] != ele[35][33];
    ele[33][32] != ele[35][34];
    ele[33][32] != ele[35][35];
    ele[33][33] != ele[33][34];
    ele[33][33] != ele[33][35];
    ele[33][33] != ele[34][30];
    ele[33][33] != ele[34][31];
    ele[33][33] != ele[34][32];
    ele[33][33] != ele[34][33];
    ele[33][33] != ele[34][34];
    ele[33][33] != ele[34][35];
    ele[33][33] != ele[35][30];
    ele[33][33] != ele[35][31];
    ele[33][33] != ele[35][32];
    ele[33][33] != ele[35][33];
    ele[33][33] != ele[35][34];
    ele[33][33] != ele[35][35];
    ele[33][34] != ele[33][35];
    ele[33][34] != ele[34][30];
    ele[33][34] != ele[34][31];
    ele[33][34] != ele[34][32];
    ele[33][34] != ele[34][33];
    ele[33][34] != ele[34][34];
    ele[33][34] != ele[34][35];
    ele[33][34] != ele[35][30];
    ele[33][34] != ele[35][31];
    ele[33][34] != ele[35][32];
    ele[33][34] != ele[35][33];
    ele[33][34] != ele[35][34];
    ele[33][34] != ele[35][35];
    ele[33][35] != ele[34][30];
    ele[33][35] != ele[34][31];
    ele[33][35] != ele[34][32];
    ele[33][35] != ele[34][33];
    ele[33][35] != ele[34][34];
    ele[33][35] != ele[34][35];
    ele[33][35] != ele[35][30];
    ele[33][35] != ele[35][31];
    ele[33][35] != ele[35][32];
    ele[33][35] != ele[35][33];
    ele[33][35] != ele[35][34];
    ele[33][35] != ele[35][35];
    ele[33][4] != ele[33][10];
    ele[33][4] != ele[33][11];
    ele[33][4] != ele[33][12];
    ele[33][4] != ele[33][13];
    ele[33][4] != ele[33][14];
    ele[33][4] != ele[33][15];
    ele[33][4] != ele[33][16];
    ele[33][4] != ele[33][17];
    ele[33][4] != ele[33][18];
    ele[33][4] != ele[33][19];
    ele[33][4] != ele[33][20];
    ele[33][4] != ele[33][21];
    ele[33][4] != ele[33][22];
    ele[33][4] != ele[33][23];
    ele[33][4] != ele[33][24];
    ele[33][4] != ele[33][25];
    ele[33][4] != ele[33][26];
    ele[33][4] != ele[33][27];
    ele[33][4] != ele[33][28];
    ele[33][4] != ele[33][29];
    ele[33][4] != ele[33][30];
    ele[33][4] != ele[33][31];
    ele[33][4] != ele[33][32];
    ele[33][4] != ele[33][33];
    ele[33][4] != ele[33][34];
    ele[33][4] != ele[33][35];
    ele[33][4] != ele[33][5];
    ele[33][4] != ele[33][6];
    ele[33][4] != ele[33][7];
    ele[33][4] != ele[33][8];
    ele[33][4] != ele[33][9];
    ele[33][4] != ele[34][0];
    ele[33][4] != ele[34][1];
    ele[33][4] != ele[34][2];
    ele[33][4] != ele[34][3];
    ele[33][4] != ele[34][4];
    ele[33][4] != ele[34][5];
    ele[33][4] != ele[35][0];
    ele[33][4] != ele[35][1];
    ele[33][4] != ele[35][2];
    ele[33][4] != ele[35][3];
    ele[33][4] != ele[35][4];
    ele[33][4] != ele[35][5];
    ele[33][5] != ele[33][10];
    ele[33][5] != ele[33][11];
    ele[33][5] != ele[33][12];
    ele[33][5] != ele[33][13];
    ele[33][5] != ele[33][14];
    ele[33][5] != ele[33][15];
    ele[33][5] != ele[33][16];
    ele[33][5] != ele[33][17];
    ele[33][5] != ele[33][18];
    ele[33][5] != ele[33][19];
    ele[33][5] != ele[33][20];
    ele[33][5] != ele[33][21];
    ele[33][5] != ele[33][22];
    ele[33][5] != ele[33][23];
    ele[33][5] != ele[33][24];
    ele[33][5] != ele[33][25];
    ele[33][5] != ele[33][26];
    ele[33][5] != ele[33][27];
    ele[33][5] != ele[33][28];
    ele[33][5] != ele[33][29];
    ele[33][5] != ele[33][30];
    ele[33][5] != ele[33][31];
    ele[33][5] != ele[33][32];
    ele[33][5] != ele[33][33];
    ele[33][5] != ele[33][34];
    ele[33][5] != ele[33][35];
    ele[33][5] != ele[33][6];
    ele[33][5] != ele[33][7];
    ele[33][5] != ele[33][8];
    ele[33][5] != ele[33][9];
    ele[33][5] != ele[34][0];
    ele[33][5] != ele[34][1];
    ele[33][5] != ele[34][2];
    ele[33][5] != ele[34][3];
    ele[33][5] != ele[34][4];
    ele[33][5] != ele[34][5];
    ele[33][5] != ele[35][0];
    ele[33][5] != ele[35][1];
    ele[33][5] != ele[35][2];
    ele[33][5] != ele[35][3];
    ele[33][5] != ele[35][4];
    ele[33][5] != ele[35][5];
    ele[33][6] != ele[33][10];
    ele[33][6] != ele[33][11];
    ele[33][6] != ele[33][12];
    ele[33][6] != ele[33][13];
    ele[33][6] != ele[33][14];
    ele[33][6] != ele[33][15];
    ele[33][6] != ele[33][16];
    ele[33][6] != ele[33][17];
    ele[33][6] != ele[33][18];
    ele[33][6] != ele[33][19];
    ele[33][6] != ele[33][20];
    ele[33][6] != ele[33][21];
    ele[33][6] != ele[33][22];
    ele[33][6] != ele[33][23];
    ele[33][6] != ele[33][24];
    ele[33][6] != ele[33][25];
    ele[33][6] != ele[33][26];
    ele[33][6] != ele[33][27];
    ele[33][6] != ele[33][28];
    ele[33][6] != ele[33][29];
    ele[33][6] != ele[33][30];
    ele[33][6] != ele[33][31];
    ele[33][6] != ele[33][32];
    ele[33][6] != ele[33][33];
    ele[33][6] != ele[33][34];
    ele[33][6] != ele[33][35];
    ele[33][6] != ele[33][7];
    ele[33][6] != ele[33][8];
    ele[33][6] != ele[33][9];
    ele[33][6] != ele[34][10];
    ele[33][6] != ele[34][11];
    ele[33][6] != ele[34][6];
    ele[33][6] != ele[34][7];
    ele[33][6] != ele[34][8];
    ele[33][6] != ele[34][9];
    ele[33][6] != ele[35][10];
    ele[33][6] != ele[35][11];
    ele[33][6] != ele[35][6];
    ele[33][6] != ele[35][7];
    ele[33][6] != ele[35][8];
    ele[33][6] != ele[35][9];
    ele[33][7] != ele[33][10];
    ele[33][7] != ele[33][11];
    ele[33][7] != ele[33][12];
    ele[33][7] != ele[33][13];
    ele[33][7] != ele[33][14];
    ele[33][7] != ele[33][15];
    ele[33][7] != ele[33][16];
    ele[33][7] != ele[33][17];
    ele[33][7] != ele[33][18];
    ele[33][7] != ele[33][19];
    ele[33][7] != ele[33][20];
    ele[33][7] != ele[33][21];
    ele[33][7] != ele[33][22];
    ele[33][7] != ele[33][23];
    ele[33][7] != ele[33][24];
    ele[33][7] != ele[33][25];
    ele[33][7] != ele[33][26];
    ele[33][7] != ele[33][27];
    ele[33][7] != ele[33][28];
    ele[33][7] != ele[33][29];
    ele[33][7] != ele[33][30];
    ele[33][7] != ele[33][31];
    ele[33][7] != ele[33][32];
    ele[33][7] != ele[33][33];
    ele[33][7] != ele[33][34];
    ele[33][7] != ele[33][35];
    ele[33][7] != ele[33][8];
    ele[33][7] != ele[33][9];
    ele[33][7] != ele[34][10];
    ele[33][7] != ele[34][11];
    ele[33][7] != ele[34][6];
    ele[33][7] != ele[34][7];
    ele[33][7] != ele[34][8];
    ele[33][7] != ele[34][9];
    ele[33][7] != ele[35][10];
    ele[33][7] != ele[35][11];
    ele[33][7] != ele[35][6];
    ele[33][7] != ele[35][7];
    ele[33][7] != ele[35][8];
    ele[33][7] != ele[35][9];
    ele[33][8] != ele[33][10];
    ele[33][8] != ele[33][11];
    ele[33][8] != ele[33][12];
    ele[33][8] != ele[33][13];
    ele[33][8] != ele[33][14];
    ele[33][8] != ele[33][15];
    ele[33][8] != ele[33][16];
    ele[33][8] != ele[33][17];
    ele[33][8] != ele[33][18];
    ele[33][8] != ele[33][19];
    ele[33][8] != ele[33][20];
    ele[33][8] != ele[33][21];
    ele[33][8] != ele[33][22];
    ele[33][8] != ele[33][23];
    ele[33][8] != ele[33][24];
    ele[33][8] != ele[33][25];
    ele[33][8] != ele[33][26];
    ele[33][8] != ele[33][27];
    ele[33][8] != ele[33][28];
    ele[33][8] != ele[33][29];
    ele[33][8] != ele[33][30];
    ele[33][8] != ele[33][31];
    ele[33][8] != ele[33][32];
    ele[33][8] != ele[33][33];
    ele[33][8] != ele[33][34];
    ele[33][8] != ele[33][35];
    ele[33][8] != ele[33][9];
    ele[33][8] != ele[34][10];
    ele[33][8] != ele[34][11];
    ele[33][8] != ele[34][6];
    ele[33][8] != ele[34][7];
    ele[33][8] != ele[34][8];
    ele[33][8] != ele[34][9];
    ele[33][8] != ele[35][10];
    ele[33][8] != ele[35][11];
    ele[33][8] != ele[35][6];
    ele[33][8] != ele[35][7];
    ele[33][8] != ele[35][8];
    ele[33][8] != ele[35][9];
    ele[33][9] != ele[33][10];
    ele[33][9] != ele[33][11];
    ele[33][9] != ele[33][12];
    ele[33][9] != ele[33][13];
    ele[33][9] != ele[33][14];
    ele[33][9] != ele[33][15];
    ele[33][9] != ele[33][16];
    ele[33][9] != ele[33][17];
    ele[33][9] != ele[33][18];
    ele[33][9] != ele[33][19];
    ele[33][9] != ele[33][20];
    ele[33][9] != ele[33][21];
    ele[33][9] != ele[33][22];
    ele[33][9] != ele[33][23];
    ele[33][9] != ele[33][24];
    ele[33][9] != ele[33][25];
    ele[33][9] != ele[33][26];
    ele[33][9] != ele[33][27];
    ele[33][9] != ele[33][28];
    ele[33][9] != ele[33][29];
    ele[33][9] != ele[33][30];
    ele[33][9] != ele[33][31];
    ele[33][9] != ele[33][32];
    ele[33][9] != ele[33][33];
    ele[33][9] != ele[33][34];
    ele[33][9] != ele[33][35];
    ele[33][9] != ele[34][10];
    ele[33][9] != ele[34][11];
    ele[33][9] != ele[34][6];
    ele[33][9] != ele[34][7];
    ele[33][9] != ele[34][8];
    ele[33][9] != ele[34][9];
    ele[33][9] != ele[35][10];
    ele[33][9] != ele[35][11];
    ele[33][9] != ele[35][6];
    ele[33][9] != ele[35][7];
    ele[33][9] != ele[35][8];
    ele[33][9] != ele[35][9];
    ele[34][0] != ele[34][1];
    ele[34][0] != ele[34][10];
    ele[34][0] != ele[34][11];
    ele[34][0] != ele[34][12];
    ele[34][0] != ele[34][13];
    ele[34][0] != ele[34][14];
    ele[34][0] != ele[34][15];
    ele[34][0] != ele[34][16];
    ele[34][0] != ele[34][17];
    ele[34][0] != ele[34][18];
    ele[34][0] != ele[34][19];
    ele[34][0] != ele[34][2];
    ele[34][0] != ele[34][20];
    ele[34][0] != ele[34][21];
    ele[34][0] != ele[34][22];
    ele[34][0] != ele[34][23];
    ele[34][0] != ele[34][24];
    ele[34][0] != ele[34][25];
    ele[34][0] != ele[34][26];
    ele[34][0] != ele[34][27];
    ele[34][0] != ele[34][28];
    ele[34][0] != ele[34][29];
    ele[34][0] != ele[34][3];
    ele[34][0] != ele[34][30];
    ele[34][0] != ele[34][31];
    ele[34][0] != ele[34][32];
    ele[34][0] != ele[34][33];
    ele[34][0] != ele[34][34];
    ele[34][0] != ele[34][35];
    ele[34][0] != ele[34][4];
    ele[34][0] != ele[34][5];
    ele[34][0] != ele[34][6];
    ele[34][0] != ele[34][7];
    ele[34][0] != ele[34][8];
    ele[34][0] != ele[34][9];
    ele[34][0] != ele[35][0];
    ele[34][0] != ele[35][1];
    ele[34][0] != ele[35][2];
    ele[34][0] != ele[35][3];
    ele[34][0] != ele[35][4];
    ele[34][0] != ele[35][5];
    ele[34][1] != ele[34][10];
    ele[34][1] != ele[34][11];
    ele[34][1] != ele[34][12];
    ele[34][1] != ele[34][13];
    ele[34][1] != ele[34][14];
    ele[34][1] != ele[34][15];
    ele[34][1] != ele[34][16];
    ele[34][1] != ele[34][17];
    ele[34][1] != ele[34][18];
    ele[34][1] != ele[34][19];
    ele[34][1] != ele[34][2];
    ele[34][1] != ele[34][20];
    ele[34][1] != ele[34][21];
    ele[34][1] != ele[34][22];
    ele[34][1] != ele[34][23];
    ele[34][1] != ele[34][24];
    ele[34][1] != ele[34][25];
    ele[34][1] != ele[34][26];
    ele[34][1] != ele[34][27];
    ele[34][1] != ele[34][28];
    ele[34][1] != ele[34][29];
    ele[34][1] != ele[34][3];
    ele[34][1] != ele[34][30];
    ele[34][1] != ele[34][31];
    ele[34][1] != ele[34][32];
    ele[34][1] != ele[34][33];
    ele[34][1] != ele[34][34];
    ele[34][1] != ele[34][35];
    ele[34][1] != ele[34][4];
    ele[34][1] != ele[34][5];
    ele[34][1] != ele[34][6];
    ele[34][1] != ele[34][7];
    ele[34][1] != ele[34][8];
    ele[34][1] != ele[34][9];
    ele[34][1] != ele[35][0];
    ele[34][1] != ele[35][1];
    ele[34][1] != ele[35][2];
    ele[34][1] != ele[35][3];
    ele[34][1] != ele[35][4];
    ele[34][1] != ele[35][5];
    ele[34][10] != ele[34][11];
    ele[34][10] != ele[34][12];
    ele[34][10] != ele[34][13];
    ele[34][10] != ele[34][14];
    ele[34][10] != ele[34][15];
    ele[34][10] != ele[34][16];
    ele[34][10] != ele[34][17];
    ele[34][10] != ele[34][18];
    ele[34][10] != ele[34][19];
    ele[34][10] != ele[34][20];
    ele[34][10] != ele[34][21];
    ele[34][10] != ele[34][22];
    ele[34][10] != ele[34][23];
    ele[34][10] != ele[34][24];
    ele[34][10] != ele[34][25];
    ele[34][10] != ele[34][26];
    ele[34][10] != ele[34][27];
    ele[34][10] != ele[34][28];
    ele[34][10] != ele[34][29];
    ele[34][10] != ele[34][30];
    ele[34][10] != ele[34][31];
    ele[34][10] != ele[34][32];
    ele[34][10] != ele[34][33];
    ele[34][10] != ele[34][34];
    ele[34][10] != ele[34][35];
    ele[34][10] != ele[35][10];
    ele[34][10] != ele[35][11];
    ele[34][10] != ele[35][6];
    ele[34][10] != ele[35][7];
    ele[34][10] != ele[35][8];
    ele[34][10] != ele[35][9];
    ele[34][11] != ele[34][12];
    ele[34][11] != ele[34][13];
    ele[34][11] != ele[34][14];
    ele[34][11] != ele[34][15];
    ele[34][11] != ele[34][16];
    ele[34][11] != ele[34][17];
    ele[34][11] != ele[34][18];
    ele[34][11] != ele[34][19];
    ele[34][11] != ele[34][20];
    ele[34][11] != ele[34][21];
    ele[34][11] != ele[34][22];
    ele[34][11] != ele[34][23];
    ele[34][11] != ele[34][24];
    ele[34][11] != ele[34][25];
    ele[34][11] != ele[34][26];
    ele[34][11] != ele[34][27];
    ele[34][11] != ele[34][28];
    ele[34][11] != ele[34][29];
    ele[34][11] != ele[34][30];
    ele[34][11] != ele[34][31];
    ele[34][11] != ele[34][32];
    ele[34][11] != ele[34][33];
    ele[34][11] != ele[34][34];
    ele[34][11] != ele[34][35];
    ele[34][11] != ele[35][10];
    ele[34][11] != ele[35][11];
    ele[34][11] != ele[35][6];
    ele[34][11] != ele[35][7];
    ele[34][11] != ele[35][8];
    ele[34][11] != ele[35][9];
    ele[34][12] != ele[34][13];
    ele[34][12] != ele[34][14];
    ele[34][12] != ele[34][15];
    ele[34][12] != ele[34][16];
    ele[34][12] != ele[34][17];
    ele[34][12] != ele[34][18];
    ele[34][12] != ele[34][19];
    ele[34][12] != ele[34][20];
    ele[34][12] != ele[34][21];
    ele[34][12] != ele[34][22];
    ele[34][12] != ele[34][23];
    ele[34][12] != ele[34][24];
    ele[34][12] != ele[34][25];
    ele[34][12] != ele[34][26];
    ele[34][12] != ele[34][27];
    ele[34][12] != ele[34][28];
    ele[34][12] != ele[34][29];
    ele[34][12] != ele[34][30];
    ele[34][12] != ele[34][31];
    ele[34][12] != ele[34][32];
    ele[34][12] != ele[34][33];
    ele[34][12] != ele[34][34];
    ele[34][12] != ele[34][35];
    ele[34][12] != ele[35][12];
    ele[34][12] != ele[35][13];
    ele[34][12] != ele[35][14];
    ele[34][12] != ele[35][15];
    ele[34][12] != ele[35][16];
    ele[34][12] != ele[35][17];
    ele[34][13] != ele[34][14];
    ele[34][13] != ele[34][15];
    ele[34][13] != ele[34][16];
    ele[34][13] != ele[34][17];
    ele[34][13] != ele[34][18];
    ele[34][13] != ele[34][19];
    ele[34][13] != ele[34][20];
    ele[34][13] != ele[34][21];
    ele[34][13] != ele[34][22];
    ele[34][13] != ele[34][23];
    ele[34][13] != ele[34][24];
    ele[34][13] != ele[34][25];
    ele[34][13] != ele[34][26];
    ele[34][13] != ele[34][27];
    ele[34][13] != ele[34][28];
    ele[34][13] != ele[34][29];
    ele[34][13] != ele[34][30];
    ele[34][13] != ele[34][31];
    ele[34][13] != ele[34][32];
    ele[34][13] != ele[34][33];
    ele[34][13] != ele[34][34];
    ele[34][13] != ele[34][35];
    ele[34][13] != ele[35][12];
    ele[34][13] != ele[35][13];
    ele[34][13] != ele[35][14];
    ele[34][13] != ele[35][15];
    ele[34][13] != ele[35][16];
    ele[34][13] != ele[35][17];
    ele[34][14] != ele[34][15];
    ele[34][14] != ele[34][16];
    ele[34][14] != ele[34][17];
    ele[34][14] != ele[34][18];
    ele[34][14] != ele[34][19];
    ele[34][14] != ele[34][20];
    ele[34][14] != ele[34][21];
    ele[34][14] != ele[34][22];
    ele[34][14] != ele[34][23];
    ele[34][14] != ele[34][24];
    ele[34][14] != ele[34][25];
    ele[34][14] != ele[34][26];
    ele[34][14] != ele[34][27];
    ele[34][14] != ele[34][28];
    ele[34][14] != ele[34][29];
    ele[34][14] != ele[34][30];
    ele[34][14] != ele[34][31];
    ele[34][14] != ele[34][32];
    ele[34][14] != ele[34][33];
    ele[34][14] != ele[34][34];
    ele[34][14] != ele[34][35];
    ele[34][14] != ele[35][12];
    ele[34][14] != ele[35][13];
    ele[34][14] != ele[35][14];
    ele[34][14] != ele[35][15];
    ele[34][14] != ele[35][16];
    ele[34][14] != ele[35][17];
    ele[34][15] != ele[34][16];
    ele[34][15] != ele[34][17];
    ele[34][15] != ele[34][18];
    ele[34][15] != ele[34][19];
    ele[34][15] != ele[34][20];
    ele[34][15] != ele[34][21];
    ele[34][15] != ele[34][22];
    ele[34][15] != ele[34][23];
    ele[34][15] != ele[34][24];
    ele[34][15] != ele[34][25];
    ele[34][15] != ele[34][26];
    ele[34][15] != ele[34][27];
    ele[34][15] != ele[34][28];
    ele[34][15] != ele[34][29];
    ele[34][15] != ele[34][30];
    ele[34][15] != ele[34][31];
    ele[34][15] != ele[34][32];
    ele[34][15] != ele[34][33];
    ele[34][15] != ele[34][34];
    ele[34][15] != ele[34][35];
    ele[34][15] != ele[35][12];
    ele[34][15] != ele[35][13];
    ele[34][15] != ele[35][14];
    ele[34][15] != ele[35][15];
    ele[34][15] != ele[35][16];
    ele[34][15] != ele[35][17];
    ele[34][16] != ele[34][17];
    ele[34][16] != ele[34][18];
    ele[34][16] != ele[34][19];
    ele[34][16] != ele[34][20];
    ele[34][16] != ele[34][21];
    ele[34][16] != ele[34][22];
    ele[34][16] != ele[34][23];
    ele[34][16] != ele[34][24];
    ele[34][16] != ele[34][25];
    ele[34][16] != ele[34][26];
    ele[34][16] != ele[34][27];
    ele[34][16] != ele[34][28];
    ele[34][16] != ele[34][29];
    ele[34][16] != ele[34][30];
    ele[34][16] != ele[34][31];
    ele[34][16] != ele[34][32];
    ele[34][16] != ele[34][33];
    ele[34][16] != ele[34][34];
    ele[34][16] != ele[34][35];
    ele[34][16] != ele[35][12];
    ele[34][16] != ele[35][13];
    ele[34][16] != ele[35][14];
    ele[34][16] != ele[35][15];
    ele[34][16] != ele[35][16];
    ele[34][16] != ele[35][17];
    ele[34][17] != ele[34][18];
    ele[34][17] != ele[34][19];
    ele[34][17] != ele[34][20];
    ele[34][17] != ele[34][21];
    ele[34][17] != ele[34][22];
    ele[34][17] != ele[34][23];
    ele[34][17] != ele[34][24];
    ele[34][17] != ele[34][25];
    ele[34][17] != ele[34][26];
    ele[34][17] != ele[34][27];
    ele[34][17] != ele[34][28];
    ele[34][17] != ele[34][29];
    ele[34][17] != ele[34][30];
    ele[34][17] != ele[34][31];
    ele[34][17] != ele[34][32];
    ele[34][17] != ele[34][33];
    ele[34][17] != ele[34][34];
    ele[34][17] != ele[34][35];
    ele[34][17] != ele[35][12];
    ele[34][17] != ele[35][13];
    ele[34][17] != ele[35][14];
    ele[34][17] != ele[35][15];
    ele[34][17] != ele[35][16];
    ele[34][17] != ele[35][17];
    ele[34][18] != ele[34][19];
    ele[34][18] != ele[34][20];
    ele[34][18] != ele[34][21];
    ele[34][18] != ele[34][22];
    ele[34][18] != ele[34][23];
    ele[34][18] != ele[34][24];
    ele[34][18] != ele[34][25];
    ele[34][18] != ele[34][26];
    ele[34][18] != ele[34][27];
    ele[34][18] != ele[34][28];
    ele[34][18] != ele[34][29];
    ele[34][18] != ele[34][30];
    ele[34][18] != ele[34][31];
    ele[34][18] != ele[34][32];
    ele[34][18] != ele[34][33];
    ele[34][18] != ele[34][34];
    ele[34][18] != ele[34][35];
    ele[34][18] != ele[35][18];
    ele[34][18] != ele[35][19];
    ele[34][18] != ele[35][20];
    ele[34][18] != ele[35][21];
    ele[34][18] != ele[35][22];
    ele[34][18] != ele[35][23];
    ele[34][19] != ele[34][20];
    ele[34][19] != ele[34][21];
    ele[34][19] != ele[34][22];
    ele[34][19] != ele[34][23];
    ele[34][19] != ele[34][24];
    ele[34][19] != ele[34][25];
    ele[34][19] != ele[34][26];
    ele[34][19] != ele[34][27];
    ele[34][19] != ele[34][28];
    ele[34][19] != ele[34][29];
    ele[34][19] != ele[34][30];
    ele[34][19] != ele[34][31];
    ele[34][19] != ele[34][32];
    ele[34][19] != ele[34][33];
    ele[34][19] != ele[34][34];
    ele[34][19] != ele[34][35];
    ele[34][19] != ele[35][18];
    ele[34][19] != ele[35][19];
    ele[34][19] != ele[35][20];
    ele[34][19] != ele[35][21];
    ele[34][19] != ele[35][22];
    ele[34][19] != ele[35][23];
    ele[34][2] != ele[34][10];
    ele[34][2] != ele[34][11];
    ele[34][2] != ele[34][12];
    ele[34][2] != ele[34][13];
    ele[34][2] != ele[34][14];
    ele[34][2] != ele[34][15];
    ele[34][2] != ele[34][16];
    ele[34][2] != ele[34][17];
    ele[34][2] != ele[34][18];
    ele[34][2] != ele[34][19];
    ele[34][2] != ele[34][20];
    ele[34][2] != ele[34][21];
    ele[34][2] != ele[34][22];
    ele[34][2] != ele[34][23];
    ele[34][2] != ele[34][24];
    ele[34][2] != ele[34][25];
    ele[34][2] != ele[34][26];
    ele[34][2] != ele[34][27];
    ele[34][2] != ele[34][28];
    ele[34][2] != ele[34][29];
    ele[34][2] != ele[34][3];
    ele[34][2] != ele[34][30];
    ele[34][2] != ele[34][31];
    ele[34][2] != ele[34][32];
    ele[34][2] != ele[34][33];
    ele[34][2] != ele[34][34];
    ele[34][2] != ele[34][35];
    ele[34][2] != ele[34][4];
    ele[34][2] != ele[34][5];
    ele[34][2] != ele[34][6];
    ele[34][2] != ele[34][7];
    ele[34][2] != ele[34][8];
    ele[34][2] != ele[34][9];
    ele[34][2] != ele[35][0];
    ele[34][2] != ele[35][1];
    ele[34][2] != ele[35][2];
    ele[34][2] != ele[35][3];
    ele[34][2] != ele[35][4];
    ele[34][2] != ele[35][5];
    ele[34][20] != ele[34][21];
    ele[34][20] != ele[34][22];
    ele[34][20] != ele[34][23];
    ele[34][20] != ele[34][24];
    ele[34][20] != ele[34][25];
    ele[34][20] != ele[34][26];
    ele[34][20] != ele[34][27];
    ele[34][20] != ele[34][28];
    ele[34][20] != ele[34][29];
    ele[34][20] != ele[34][30];
    ele[34][20] != ele[34][31];
    ele[34][20] != ele[34][32];
    ele[34][20] != ele[34][33];
    ele[34][20] != ele[34][34];
    ele[34][20] != ele[34][35];
    ele[34][20] != ele[35][18];
    ele[34][20] != ele[35][19];
    ele[34][20] != ele[35][20];
    ele[34][20] != ele[35][21];
    ele[34][20] != ele[35][22];
    ele[34][20] != ele[35][23];
    ele[34][21] != ele[34][22];
    ele[34][21] != ele[34][23];
    ele[34][21] != ele[34][24];
    ele[34][21] != ele[34][25];
    ele[34][21] != ele[34][26];
    ele[34][21] != ele[34][27];
    ele[34][21] != ele[34][28];
    ele[34][21] != ele[34][29];
    ele[34][21] != ele[34][30];
    ele[34][21] != ele[34][31];
    ele[34][21] != ele[34][32];
    ele[34][21] != ele[34][33];
    ele[34][21] != ele[34][34];
    ele[34][21] != ele[34][35];
    ele[34][21] != ele[35][18];
    ele[34][21] != ele[35][19];
    ele[34][21] != ele[35][20];
    ele[34][21] != ele[35][21];
    ele[34][21] != ele[35][22];
    ele[34][21] != ele[35][23];
    ele[34][22] != ele[34][23];
    ele[34][22] != ele[34][24];
    ele[34][22] != ele[34][25];
    ele[34][22] != ele[34][26];
    ele[34][22] != ele[34][27];
    ele[34][22] != ele[34][28];
    ele[34][22] != ele[34][29];
    ele[34][22] != ele[34][30];
    ele[34][22] != ele[34][31];
    ele[34][22] != ele[34][32];
    ele[34][22] != ele[34][33];
    ele[34][22] != ele[34][34];
    ele[34][22] != ele[34][35];
    ele[34][22] != ele[35][18];
    ele[34][22] != ele[35][19];
    ele[34][22] != ele[35][20];
    ele[34][22] != ele[35][21];
    ele[34][22] != ele[35][22];
    ele[34][22] != ele[35][23];
    ele[34][23] != ele[34][24];
    ele[34][23] != ele[34][25];
    ele[34][23] != ele[34][26];
    ele[34][23] != ele[34][27];
    ele[34][23] != ele[34][28];
    ele[34][23] != ele[34][29];
    ele[34][23] != ele[34][30];
    ele[34][23] != ele[34][31];
    ele[34][23] != ele[34][32];
    ele[34][23] != ele[34][33];
    ele[34][23] != ele[34][34];
    ele[34][23] != ele[34][35];
    ele[34][23] != ele[35][18];
    ele[34][23] != ele[35][19];
    ele[34][23] != ele[35][20];
    ele[34][23] != ele[35][21];
    ele[34][23] != ele[35][22];
    ele[34][23] != ele[35][23];
    ele[34][24] != ele[34][25];
    ele[34][24] != ele[34][26];
    ele[34][24] != ele[34][27];
    ele[34][24] != ele[34][28];
    ele[34][24] != ele[34][29];
    ele[34][24] != ele[34][30];
    ele[34][24] != ele[34][31];
    ele[34][24] != ele[34][32];
    ele[34][24] != ele[34][33];
    ele[34][24] != ele[34][34];
    ele[34][24] != ele[34][35];
    ele[34][24] != ele[35][24];
    ele[34][24] != ele[35][25];
    ele[34][24] != ele[35][26];
    ele[34][24] != ele[35][27];
    ele[34][24] != ele[35][28];
    ele[34][24] != ele[35][29];
    ele[34][25] != ele[34][26];
    ele[34][25] != ele[34][27];
    ele[34][25] != ele[34][28];
    ele[34][25] != ele[34][29];
    ele[34][25] != ele[34][30];
    ele[34][25] != ele[34][31];
    ele[34][25] != ele[34][32];
    ele[34][25] != ele[34][33];
    ele[34][25] != ele[34][34];
    ele[34][25] != ele[34][35];
    ele[34][25] != ele[35][24];
    ele[34][25] != ele[35][25];
    ele[34][25] != ele[35][26];
    ele[34][25] != ele[35][27];
    ele[34][25] != ele[35][28];
    ele[34][25] != ele[35][29];
    ele[34][26] != ele[34][27];
    ele[34][26] != ele[34][28];
    ele[34][26] != ele[34][29];
    ele[34][26] != ele[34][30];
    ele[34][26] != ele[34][31];
    ele[34][26] != ele[34][32];
    ele[34][26] != ele[34][33];
    ele[34][26] != ele[34][34];
    ele[34][26] != ele[34][35];
    ele[34][26] != ele[35][24];
    ele[34][26] != ele[35][25];
    ele[34][26] != ele[35][26];
    ele[34][26] != ele[35][27];
    ele[34][26] != ele[35][28];
    ele[34][26] != ele[35][29];
    ele[34][27] != ele[34][28];
    ele[34][27] != ele[34][29];
    ele[34][27] != ele[34][30];
    ele[34][27] != ele[34][31];
    ele[34][27] != ele[34][32];
    ele[34][27] != ele[34][33];
    ele[34][27] != ele[34][34];
    ele[34][27] != ele[34][35];
    ele[34][27] != ele[35][24];
    ele[34][27] != ele[35][25];
    ele[34][27] != ele[35][26];
    ele[34][27] != ele[35][27];
    ele[34][27] != ele[35][28];
    ele[34][27] != ele[35][29];
    ele[34][28] != ele[34][29];
    ele[34][28] != ele[34][30];
    ele[34][28] != ele[34][31];
    ele[34][28] != ele[34][32];
    ele[34][28] != ele[34][33];
    ele[34][28] != ele[34][34];
    ele[34][28] != ele[34][35];
    ele[34][28] != ele[35][24];
    ele[34][28] != ele[35][25];
    ele[34][28] != ele[35][26];
    ele[34][28] != ele[35][27];
    ele[34][28] != ele[35][28];
    ele[34][28] != ele[35][29];
    ele[34][29] != ele[34][30];
    ele[34][29] != ele[34][31];
    ele[34][29] != ele[34][32];
    ele[34][29] != ele[34][33];
    ele[34][29] != ele[34][34];
    ele[34][29] != ele[34][35];
    ele[34][29] != ele[35][24];
    ele[34][29] != ele[35][25];
    ele[34][29] != ele[35][26];
    ele[34][29] != ele[35][27];
    ele[34][29] != ele[35][28];
    ele[34][29] != ele[35][29];
    ele[34][3] != ele[34][10];
    ele[34][3] != ele[34][11];
    ele[34][3] != ele[34][12];
    ele[34][3] != ele[34][13];
    ele[34][3] != ele[34][14];
    ele[34][3] != ele[34][15];
    ele[34][3] != ele[34][16];
    ele[34][3] != ele[34][17];
    ele[34][3] != ele[34][18];
    ele[34][3] != ele[34][19];
    ele[34][3] != ele[34][20];
    ele[34][3] != ele[34][21];
    ele[34][3] != ele[34][22];
    ele[34][3] != ele[34][23];
    ele[34][3] != ele[34][24];
    ele[34][3] != ele[34][25];
    ele[34][3] != ele[34][26];
    ele[34][3] != ele[34][27];
    ele[34][3] != ele[34][28];
    ele[34][3] != ele[34][29];
    ele[34][3] != ele[34][30];
    ele[34][3] != ele[34][31];
    ele[34][3] != ele[34][32];
    ele[34][3] != ele[34][33];
    ele[34][3] != ele[34][34];
    ele[34][3] != ele[34][35];
    ele[34][3] != ele[34][4];
    ele[34][3] != ele[34][5];
    ele[34][3] != ele[34][6];
    ele[34][3] != ele[34][7];
    ele[34][3] != ele[34][8];
    ele[34][3] != ele[34][9];
    ele[34][3] != ele[35][0];
    ele[34][3] != ele[35][1];
    ele[34][3] != ele[35][2];
    ele[34][3] != ele[35][3];
    ele[34][3] != ele[35][4];
    ele[34][3] != ele[35][5];
    ele[34][30] != ele[34][31];
    ele[34][30] != ele[34][32];
    ele[34][30] != ele[34][33];
    ele[34][30] != ele[34][34];
    ele[34][30] != ele[34][35];
    ele[34][30] != ele[35][30];
    ele[34][30] != ele[35][31];
    ele[34][30] != ele[35][32];
    ele[34][30] != ele[35][33];
    ele[34][30] != ele[35][34];
    ele[34][30] != ele[35][35];
    ele[34][31] != ele[34][32];
    ele[34][31] != ele[34][33];
    ele[34][31] != ele[34][34];
    ele[34][31] != ele[34][35];
    ele[34][31] != ele[35][30];
    ele[34][31] != ele[35][31];
    ele[34][31] != ele[35][32];
    ele[34][31] != ele[35][33];
    ele[34][31] != ele[35][34];
    ele[34][31] != ele[35][35];
    ele[34][32] != ele[34][33];
    ele[34][32] != ele[34][34];
    ele[34][32] != ele[34][35];
    ele[34][32] != ele[35][30];
    ele[34][32] != ele[35][31];
    ele[34][32] != ele[35][32];
    ele[34][32] != ele[35][33];
    ele[34][32] != ele[35][34];
    ele[34][32] != ele[35][35];
    ele[34][33] != ele[34][34];
    ele[34][33] != ele[34][35];
    ele[34][33] != ele[35][30];
    ele[34][33] != ele[35][31];
    ele[34][33] != ele[35][32];
    ele[34][33] != ele[35][33];
    ele[34][33] != ele[35][34];
    ele[34][33] != ele[35][35];
    ele[34][34] != ele[34][35];
    ele[34][34] != ele[35][30];
    ele[34][34] != ele[35][31];
    ele[34][34] != ele[35][32];
    ele[34][34] != ele[35][33];
    ele[34][34] != ele[35][34];
    ele[34][34] != ele[35][35];
    ele[34][35] != ele[35][30];
    ele[34][35] != ele[35][31];
    ele[34][35] != ele[35][32];
    ele[34][35] != ele[35][33];
    ele[34][35] != ele[35][34];
    ele[34][35] != ele[35][35];
    ele[34][4] != ele[34][10];
    ele[34][4] != ele[34][11];
    ele[34][4] != ele[34][12];
    ele[34][4] != ele[34][13];
    ele[34][4] != ele[34][14];
    ele[34][4] != ele[34][15];
    ele[34][4] != ele[34][16];
    ele[34][4] != ele[34][17];
    ele[34][4] != ele[34][18];
    ele[34][4] != ele[34][19];
    ele[34][4] != ele[34][20];
    ele[34][4] != ele[34][21];
    ele[34][4] != ele[34][22];
    ele[34][4] != ele[34][23];
    ele[34][4] != ele[34][24];
    ele[34][4] != ele[34][25];
    ele[34][4] != ele[34][26];
    ele[34][4] != ele[34][27];
    ele[34][4] != ele[34][28];
    ele[34][4] != ele[34][29];
    ele[34][4] != ele[34][30];
    ele[34][4] != ele[34][31];
    ele[34][4] != ele[34][32];
    ele[34][4] != ele[34][33];
    ele[34][4] != ele[34][34];
    ele[34][4] != ele[34][35];
    ele[34][4] != ele[34][5];
    ele[34][4] != ele[34][6];
    ele[34][4] != ele[34][7];
    ele[34][4] != ele[34][8];
    ele[34][4] != ele[34][9];
    ele[34][4] != ele[35][0];
    ele[34][4] != ele[35][1];
    ele[34][4] != ele[35][2];
    ele[34][4] != ele[35][3];
    ele[34][4] != ele[35][4];
    ele[34][4] != ele[35][5];
    ele[34][5] != ele[34][10];
    ele[34][5] != ele[34][11];
    ele[34][5] != ele[34][12];
    ele[34][5] != ele[34][13];
    ele[34][5] != ele[34][14];
    ele[34][5] != ele[34][15];
    ele[34][5] != ele[34][16];
    ele[34][5] != ele[34][17];
    ele[34][5] != ele[34][18];
    ele[34][5] != ele[34][19];
    ele[34][5] != ele[34][20];
    ele[34][5] != ele[34][21];
    ele[34][5] != ele[34][22];
    ele[34][5] != ele[34][23];
    ele[34][5] != ele[34][24];
    ele[34][5] != ele[34][25];
    ele[34][5] != ele[34][26];
    ele[34][5] != ele[34][27];
    ele[34][5] != ele[34][28];
    ele[34][5] != ele[34][29];
    ele[34][5] != ele[34][30];
    ele[34][5] != ele[34][31];
    ele[34][5] != ele[34][32];
    ele[34][5] != ele[34][33];
    ele[34][5] != ele[34][34];
    ele[34][5] != ele[34][35];
    ele[34][5] != ele[34][6];
    ele[34][5] != ele[34][7];
    ele[34][5] != ele[34][8];
    ele[34][5] != ele[34][9];
    ele[34][5] != ele[35][0];
    ele[34][5] != ele[35][1];
    ele[34][5] != ele[35][2];
    ele[34][5] != ele[35][3];
    ele[34][5] != ele[35][4];
    ele[34][5] != ele[35][5];
    ele[34][6] != ele[34][10];
    ele[34][6] != ele[34][11];
    ele[34][6] != ele[34][12];
    ele[34][6] != ele[34][13];
    ele[34][6] != ele[34][14];
    ele[34][6] != ele[34][15];
    ele[34][6] != ele[34][16];
    ele[34][6] != ele[34][17];
    ele[34][6] != ele[34][18];
    ele[34][6] != ele[34][19];
    ele[34][6] != ele[34][20];
    ele[34][6] != ele[34][21];
    ele[34][6] != ele[34][22];
    ele[34][6] != ele[34][23];
    ele[34][6] != ele[34][24];
    ele[34][6] != ele[34][25];
    ele[34][6] != ele[34][26];
    ele[34][6] != ele[34][27];
    ele[34][6] != ele[34][28];
    ele[34][6] != ele[34][29];
    ele[34][6] != ele[34][30];
    ele[34][6] != ele[34][31];
    ele[34][6] != ele[34][32];
    ele[34][6] != ele[34][33];
    ele[34][6] != ele[34][34];
    ele[34][6] != ele[34][35];
    ele[34][6] != ele[34][7];
    ele[34][6] != ele[34][8];
    ele[34][6] != ele[34][9];
    ele[34][6] != ele[35][10];
    ele[34][6] != ele[35][11];
    ele[34][6] != ele[35][6];
    ele[34][6] != ele[35][7];
    ele[34][6] != ele[35][8];
    ele[34][6] != ele[35][9];
    ele[34][7] != ele[34][10];
    ele[34][7] != ele[34][11];
    ele[34][7] != ele[34][12];
    ele[34][7] != ele[34][13];
    ele[34][7] != ele[34][14];
    ele[34][7] != ele[34][15];
    ele[34][7] != ele[34][16];
    ele[34][7] != ele[34][17];
    ele[34][7] != ele[34][18];
    ele[34][7] != ele[34][19];
    ele[34][7] != ele[34][20];
    ele[34][7] != ele[34][21];
    ele[34][7] != ele[34][22];
    ele[34][7] != ele[34][23];
    ele[34][7] != ele[34][24];
    ele[34][7] != ele[34][25];
    ele[34][7] != ele[34][26];
    ele[34][7] != ele[34][27];
    ele[34][7] != ele[34][28];
    ele[34][7] != ele[34][29];
    ele[34][7] != ele[34][30];
    ele[34][7] != ele[34][31];
    ele[34][7] != ele[34][32];
    ele[34][7] != ele[34][33];
    ele[34][7] != ele[34][34];
    ele[34][7] != ele[34][35];
    ele[34][7] != ele[34][8];
    ele[34][7] != ele[34][9];
    ele[34][7] != ele[35][10];
    ele[34][7] != ele[35][11];
    ele[34][7] != ele[35][6];
    ele[34][7] != ele[35][7];
    ele[34][7] != ele[35][8];
    ele[34][7] != ele[35][9];
    ele[34][8] != ele[34][10];
    ele[34][8] != ele[34][11];
    ele[34][8] != ele[34][12];
    ele[34][8] != ele[34][13];
    ele[34][8] != ele[34][14];
    ele[34][8] != ele[34][15];
    ele[34][8] != ele[34][16];
    ele[34][8] != ele[34][17];
    ele[34][8] != ele[34][18];
    ele[34][8] != ele[34][19];
    ele[34][8] != ele[34][20];
    ele[34][8] != ele[34][21];
    ele[34][8] != ele[34][22];
    ele[34][8] != ele[34][23];
    ele[34][8] != ele[34][24];
    ele[34][8] != ele[34][25];
    ele[34][8] != ele[34][26];
    ele[34][8] != ele[34][27];
    ele[34][8] != ele[34][28];
    ele[34][8] != ele[34][29];
    ele[34][8] != ele[34][30];
    ele[34][8] != ele[34][31];
    ele[34][8] != ele[34][32];
    ele[34][8] != ele[34][33];
    ele[34][8] != ele[34][34];
    ele[34][8] != ele[34][35];
    ele[34][8] != ele[34][9];
    ele[34][8] != ele[35][10];
    ele[34][8] != ele[35][11];
    ele[34][8] != ele[35][6];
    ele[34][8] != ele[35][7];
    ele[34][8] != ele[35][8];
    ele[34][8] != ele[35][9];
    ele[34][9] != ele[34][10];
    ele[34][9] != ele[34][11];
    ele[34][9] != ele[34][12];
    ele[34][9] != ele[34][13];
    ele[34][9] != ele[34][14];
    ele[34][9] != ele[34][15];
    ele[34][9] != ele[34][16];
    ele[34][9] != ele[34][17];
    ele[34][9] != ele[34][18];
    ele[34][9] != ele[34][19];
    ele[34][9] != ele[34][20];
    ele[34][9] != ele[34][21];
    ele[34][9] != ele[34][22];
    ele[34][9] != ele[34][23];
    ele[34][9] != ele[34][24];
    ele[34][9] != ele[34][25];
    ele[34][9] != ele[34][26];
    ele[34][9] != ele[34][27];
    ele[34][9] != ele[34][28];
    ele[34][9] != ele[34][29];
    ele[34][9] != ele[34][30];
    ele[34][9] != ele[34][31];
    ele[34][9] != ele[34][32];
    ele[34][9] != ele[34][33];
    ele[34][9] != ele[34][34];
    ele[34][9] != ele[34][35];
    ele[34][9] != ele[35][10];
    ele[34][9] != ele[35][11];
    ele[34][9] != ele[35][6];
    ele[34][9] != ele[35][7];
    ele[34][9] != ele[35][8];
    ele[34][9] != ele[35][9];
    ele[35][0] != ele[35][1];
    ele[35][0] != ele[35][10];
    ele[35][0] != ele[35][11];
    ele[35][0] != ele[35][12];
    ele[35][0] != ele[35][13];
    ele[35][0] != ele[35][14];
    ele[35][0] != ele[35][15];
    ele[35][0] != ele[35][16];
    ele[35][0] != ele[35][17];
    ele[35][0] != ele[35][18];
    ele[35][0] != ele[35][19];
    ele[35][0] != ele[35][2];
    ele[35][0] != ele[35][20];
    ele[35][0] != ele[35][21];
    ele[35][0] != ele[35][22];
    ele[35][0] != ele[35][23];
    ele[35][0] != ele[35][24];
    ele[35][0] != ele[35][25];
    ele[35][0] != ele[35][26];
    ele[35][0] != ele[35][27];
    ele[35][0] != ele[35][28];
    ele[35][0] != ele[35][29];
    ele[35][0] != ele[35][3];
    ele[35][0] != ele[35][30];
    ele[35][0] != ele[35][31];
    ele[35][0] != ele[35][32];
    ele[35][0] != ele[35][33];
    ele[35][0] != ele[35][34];
    ele[35][0] != ele[35][35];
    ele[35][0] != ele[35][4];
    ele[35][0] != ele[35][5];
    ele[35][0] != ele[35][6];
    ele[35][0] != ele[35][7];
    ele[35][0] != ele[35][8];
    ele[35][0] != ele[35][9];
    ele[35][1] != ele[35][10];
    ele[35][1] != ele[35][11];
    ele[35][1] != ele[35][12];
    ele[35][1] != ele[35][13];
    ele[35][1] != ele[35][14];
    ele[35][1] != ele[35][15];
    ele[35][1] != ele[35][16];
    ele[35][1] != ele[35][17];
    ele[35][1] != ele[35][18];
    ele[35][1] != ele[35][19];
    ele[35][1] != ele[35][2];
    ele[35][1] != ele[35][20];
    ele[35][1] != ele[35][21];
    ele[35][1] != ele[35][22];
    ele[35][1] != ele[35][23];
    ele[35][1] != ele[35][24];
    ele[35][1] != ele[35][25];
    ele[35][1] != ele[35][26];
    ele[35][1] != ele[35][27];
    ele[35][1] != ele[35][28];
    ele[35][1] != ele[35][29];
    ele[35][1] != ele[35][3];
    ele[35][1] != ele[35][30];
    ele[35][1] != ele[35][31];
    ele[35][1] != ele[35][32];
    ele[35][1] != ele[35][33];
    ele[35][1] != ele[35][34];
    ele[35][1] != ele[35][35];
    ele[35][1] != ele[35][4];
    ele[35][1] != ele[35][5];
    ele[35][1] != ele[35][6];
    ele[35][1] != ele[35][7];
    ele[35][1] != ele[35][8];
    ele[35][1] != ele[35][9];
    ele[35][10] != ele[35][11];
    ele[35][10] != ele[35][12];
    ele[35][10] != ele[35][13];
    ele[35][10] != ele[35][14];
    ele[35][10] != ele[35][15];
    ele[35][10] != ele[35][16];
    ele[35][10] != ele[35][17];
    ele[35][10] != ele[35][18];
    ele[35][10] != ele[35][19];
    ele[35][10] != ele[35][20];
    ele[35][10] != ele[35][21];
    ele[35][10] != ele[35][22];
    ele[35][10] != ele[35][23];
    ele[35][10] != ele[35][24];
    ele[35][10] != ele[35][25];
    ele[35][10] != ele[35][26];
    ele[35][10] != ele[35][27];
    ele[35][10] != ele[35][28];
    ele[35][10] != ele[35][29];
    ele[35][10] != ele[35][30];
    ele[35][10] != ele[35][31];
    ele[35][10] != ele[35][32];
    ele[35][10] != ele[35][33];
    ele[35][10] != ele[35][34];
    ele[35][10] != ele[35][35];
    ele[35][11] != ele[35][12];
    ele[35][11] != ele[35][13];
    ele[35][11] != ele[35][14];
    ele[35][11] != ele[35][15];
    ele[35][11] != ele[35][16];
    ele[35][11] != ele[35][17];
    ele[35][11] != ele[35][18];
    ele[35][11] != ele[35][19];
    ele[35][11] != ele[35][20];
    ele[35][11] != ele[35][21];
    ele[35][11] != ele[35][22];
    ele[35][11] != ele[35][23];
    ele[35][11] != ele[35][24];
    ele[35][11] != ele[35][25];
    ele[35][11] != ele[35][26];
    ele[35][11] != ele[35][27];
    ele[35][11] != ele[35][28];
    ele[35][11] != ele[35][29];
    ele[35][11] != ele[35][30];
    ele[35][11] != ele[35][31];
    ele[35][11] != ele[35][32];
    ele[35][11] != ele[35][33];
    ele[35][11] != ele[35][34];
    ele[35][11] != ele[35][35];
    ele[35][12] != ele[35][13];
    ele[35][12] != ele[35][14];
    ele[35][12] != ele[35][15];
    ele[35][12] != ele[35][16];
    ele[35][12] != ele[35][17];
    ele[35][12] != ele[35][18];
    ele[35][12] != ele[35][19];
    ele[35][12] != ele[35][20];
    ele[35][12] != ele[35][21];
    ele[35][12] != ele[35][22];
    ele[35][12] != ele[35][23];
    ele[35][12] != ele[35][24];
    ele[35][12] != ele[35][25];
    ele[35][12] != ele[35][26];
    ele[35][12] != ele[35][27];
    ele[35][12] != ele[35][28];
    ele[35][12] != ele[35][29];
    ele[35][12] != ele[35][30];
    ele[35][12] != ele[35][31];
    ele[35][12] != ele[35][32];
    ele[35][12] != ele[35][33];
    ele[35][12] != ele[35][34];
    ele[35][12] != ele[35][35];
    ele[35][13] != ele[35][14];
    ele[35][13] != ele[35][15];
    ele[35][13] != ele[35][16];
    ele[35][13] != ele[35][17];
    ele[35][13] != ele[35][18];
    ele[35][13] != ele[35][19];
    ele[35][13] != ele[35][20];
    ele[35][13] != ele[35][21];
    ele[35][13] != ele[35][22];
    ele[35][13] != ele[35][23];
    ele[35][13] != ele[35][24];
    ele[35][13] != ele[35][25];
    ele[35][13] != ele[35][26];
    ele[35][13] != ele[35][27];
    ele[35][13] != ele[35][28];
    ele[35][13] != ele[35][29];
    ele[35][13] != ele[35][30];
    ele[35][13] != ele[35][31];
    ele[35][13] != ele[35][32];
    ele[35][13] != ele[35][33];
    ele[35][13] != ele[35][34];
    ele[35][13] != ele[35][35];
    ele[35][14] != ele[35][15];
    ele[35][14] != ele[35][16];
    ele[35][14] != ele[35][17];
    ele[35][14] != ele[35][18];
    ele[35][14] != ele[35][19];
    ele[35][14] != ele[35][20];
    ele[35][14] != ele[35][21];
    ele[35][14] != ele[35][22];
    ele[35][14] != ele[35][23];
    ele[35][14] != ele[35][24];
    ele[35][14] != ele[35][25];
    ele[35][14] != ele[35][26];
    ele[35][14] != ele[35][27];
    ele[35][14] != ele[35][28];
    ele[35][14] != ele[35][29];
    ele[35][14] != ele[35][30];
    ele[35][14] != ele[35][31];
    ele[35][14] != ele[35][32];
    ele[35][14] != ele[35][33];
    ele[35][14] != ele[35][34];
    ele[35][14] != ele[35][35];
    ele[35][15] != ele[35][16];
    ele[35][15] != ele[35][17];
    ele[35][15] != ele[35][18];
    ele[35][15] != ele[35][19];
    ele[35][15] != ele[35][20];
    ele[35][15] != ele[35][21];
    ele[35][15] != ele[35][22];
    ele[35][15] != ele[35][23];
    ele[35][15] != ele[35][24];
    ele[35][15] != ele[35][25];
    ele[35][15] != ele[35][26];
    ele[35][15] != ele[35][27];
    ele[35][15] != ele[35][28];
    ele[35][15] != ele[35][29];
    ele[35][15] != ele[35][30];
    ele[35][15] != ele[35][31];
    ele[35][15] != ele[35][32];
    ele[35][15] != ele[35][33];
    ele[35][15] != ele[35][34];
    ele[35][15] != ele[35][35];
    ele[35][16] != ele[35][17];
    ele[35][16] != ele[35][18];
    ele[35][16] != ele[35][19];
    ele[35][16] != ele[35][20];
    ele[35][16] != ele[35][21];
    ele[35][16] != ele[35][22];
    ele[35][16] != ele[35][23];
    ele[35][16] != ele[35][24];
    ele[35][16] != ele[35][25];
    ele[35][16] != ele[35][26];
    ele[35][16] != ele[35][27];
    ele[35][16] != ele[35][28];
    ele[35][16] != ele[35][29];
    ele[35][16] != ele[35][30];
    ele[35][16] != ele[35][31];
    ele[35][16] != ele[35][32];
    ele[35][16] != ele[35][33];
    ele[35][16] != ele[35][34];
    ele[35][16] != ele[35][35];
    ele[35][17] != ele[35][18];
    ele[35][17] != ele[35][19];
    ele[35][17] != ele[35][20];
    ele[35][17] != ele[35][21];
    ele[35][17] != ele[35][22];
    ele[35][17] != ele[35][23];
    ele[35][17] != ele[35][24];
    ele[35][17] != ele[35][25];
    ele[35][17] != ele[35][26];
    ele[35][17] != ele[35][27];
    ele[35][17] != ele[35][28];
    ele[35][17] != ele[35][29];
    ele[35][17] != ele[35][30];
    ele[35][17] != ele[35][31];
    ele[35][17] != ele[35][32];
    ele[35][17] != ele[35][33];
    ele[35][17] != ele[35][34];
    ele[35][17] != ele[35][35];
    ele[35][18] != ele[35][19];
    ele[35][18] != ele[35][20];
    ele[35][18] != ele[35][21];
    ele[35][18] != ele[35][22];
    ele[35][18] != ele[35][23];
    ele[35][18] != ele[35][24];
    ele[35][18] != ele[35][25];
    ele[35][18] != ele[35][26];
    ele[35][18] != ele[35][27];
    ele[35][18] != ele[35][28];
    ele[35][18] != ele[35][29];
    ele[35][18] != ele[35][30];
    ele[35][18] != ele[35][31];
    ele[35][18] != ele[35][32];
    ele[35][18] != ele[35][33];
    ele[35][18] != ele[35][34];
    ele[35][18] != ele[35][35];
    ele[35][19] != ele[35][20];
    ele[35][19] != ele[35][21];
    ele[35][19] != ele[35][22];
    ele[35][19] != ele[35][23];
    ele[35][19] != ele[35][24];
    ele[35][19] != ele[35][25];
    ele[35][19] != ele[35][26];
    ele[35][19] != ele[35][27];
    ele[35][19] != ele[35][28];
    ele[35][19] != ele[35][29];
    ele[35][19] != ele[35][30];
    ele[35][19] != ele[35][31];
    ele[35][19] != ele[35][32];
    ele[35][19] != ele[35][33];
    ele[35][19] != ele[35][34];
    ele[35][19] != ele[35][35];
    ele[35][2] != ele[35][10];
    ele[35][2] != ele[35][11];
    ele[35][2] != ele[35][12];
    ele[35][2] != ele[35][13];
    ele[35][2] != ele[35][14];
    ele[35][2] != ele[35][15];
    ele[35][2] != ele[35][16];
    ele[35][2] != ele[35][17];
    ele[35][2] != ele[35][18];
    ele[35][2] != ele[35][19];
    ele[35][2] != ele[35][20];
    ele[35][2] != ele[35][21];
    ele[35][2] != ele[35][22];
    ele[35][2] != ele[35][23];
    ele[35][2] != ele[35][24];
    ele[35][2] != ele[35][25];
    ele[35][2] != ele[35][26];
    ele[35][2] != ele[35][27];
    ele[35][2] != ele[35][28];
    ele[35][2] != ele[35][29];
    ele[35][2] != ele[35][3];
    ele[35][2] != ele[35][30];
    ele[35][2] != ele[35][31];
    ele[35][2] != ele[35][32];
    ele[35][2] != ele[35][33];
    ele[35][2] != ele[35][34];
    ele[35][2] != ele[35][35];
    ele[35][2] != ele[35][4];
    ele[35][2] != ele[35][5];
    ele[35][2] != ele[35][6];
    ele[35][2] != ele[35][7];
    ele[35][2] != ele[35][8];
    ele[35][2] != ele[35][9];
    ele[35][20] != ele[35][21];
    ele[35][20] != ele[35][22];
    ele[35][20] != ele[35][23];
    ele[35][20] != ele[35][24];
    ele[35][20] != ele[35][25];
    ele[35][20] != ele[35][26];
    ele[35][20] != ele[35][27];
    ele[35][20] != ele[35][28];
    ele[35][20] != ele[35][29];
    ele[35][20] != ele[35][30];
    ele[35][20] != ele[35][31];
    ele[35][20] != ele[35][32];
    ele[35][20] != ele[35][33];
    ele[35][20] != ele[35][34];
    ele[35][20] != ele[35][35];
    ele[35][21] != ele[35][22];
    ele[35][21] != ele[35][23];
    ele[35][21] != ele[35][24];
    ele[35][21] != ele[35][25];
    ele[35][21] != ele[35][26];
    ele[35][21] != ele[35][27];
    ele[35][21] != ele[35][28];
    ele[35][21] != ele[35][29];
    ele[35][21] != ele[35][30];
    ele[35][21] != ele[35][31];
    ele[35][21] != ele[35][32];
    ele[35][21] != ele[35][33];
    ele[35][21] != ele[35][34];
    ele[35][21] != ele[35][35];
    ele[35][22] != ele[35][23];
    ele[35][22] != ele[35][24];
    ele[35][22] != ele[35][25];
    ele[35][22] != ele[35][26];
    ele[35][22] != ele[35][27];
    ele[35][22] != ele[35][28];
    ele[35][22] != ele[35][29];
    ele[35][22] != ele[35][30];
    ele[35][22] != ele[35][31];
    ele[35][22] != ele[35][32];
    ele[35][22] != ele[35][33];
    ele[35][22] != ele[35][34];
    ele[35][22] != ele[35][35];
    ele[35][23] != ele[35][24];
    ele[35][23] != ele[35][25];
    ele[35][23] != ele[35][26];
    ele[35][23] != ele[35][27];
    ele[35][23] != ele[35][28];
    ele[35][23] != ele[35][29];
    ele[35][23] != ele[35][30];
    ele[35][23] != ele[35][31];
    ele[35][23] != ele[35][32];
    ele[35][23] != ele[35][33];
    ele[35][23] != ele[35][34];
    ele[35][23] != ele[35][35];
    ele[35][24] != ele[35][25];
    ele[35][24] != ele[35][26];
    ele[35][24] != ele[35][27];
    ele[35][24] != ele[35][28];
    ele[35][24] != ele[35][29];
    ele[35][24] != ele[35][30];
    ele[35][24] != ele[35][31];
    ele[35][24] != ele[35][32];
    ele[35][24] != ele[35][33];
    ele[35][24] != ele[35][34];
    ele[35][24] != ele[35][35];
    ele[35][25] != ele[35][26];
    ele[35][25] != ele[35][27];
    ele[35][25] != ele[35][28];
    ele[35][25] != ele[35][29];
    ele[35][25] != ele[35][30];
    ele[35][25] != ele[35][31];
    ele[35][25] != ele[35][32];
    ele[35][25] != ele[35][33];
    ele[35][25] != ele[35][34];
    ele[35][25] != ele[35][35];
    ele[35][26] != ele[35][27];
    ele[35][26] != ele[35][28];
    ele[35][26] != ele[35][29];
    ele[35][26] != ele[35][30];
    ele[35][26] != ele[35][31];
    ele[35][26] != ele[35][32];
    ele[35][26] != ele[35][33];
    ele[35][26] != ele[35][34];
    ele[35][26] != ele[35][35];
    ele[35][27] != ele[35][28];
    ele[35][27] != ele[35][29];
    ele[35][27] != ele[35][30];
    ele[35][27] != ele[35][31];
    ele[35][27] != ele[35][32];
    ele[35][27] != ele[35][33];
    ele[35][27] != ele[35][34];
    ele[35][27] != ele[35][35];
    ele[35][28] != ele[35][29];
    ele[35][28] != ele[35][30];
    ele[35][28] != ele[35][31];
    ele[35][28] != ele[35][32];
    ele[35][28] != ele[35][33];
    ele[35][28] != ele[35][34];
    ele[35][28] != ele[35][35];
    ele[35][29] != ele[35][30];
    ele[35][29] != ele[35][31];
    ele[35][29] != ele[35][32];
    ele[35][29] != ele[35][33];
    ele[35][29] != ele[35][34];
    ele[35][29] != ele[35][35];
    ele[35][3] != ele[35][10];
    ele[35][3] != ele[35][11];
    ele[35][3] != ele[35][12];
    ele[35][3] != ele[35][13];
    ele[35][3] != ele[35][14];
    ele[35][3] != ele[35][15];
    ele[35][3] != ele[35][16];
    ele[35][3] != ele[35][17];
    ele[35][3] != ele[35][18];
    ele[35][3] != ele[35][19];
    ele[35][3] != ele[35][20];
    ele[35][3] != ele[35][21];
    ele[35][3] != ele[35][22];
    ele[35][3] != ele[35][23];
    ele[35][3] != ele[35][24];
    ele[35][3] != ele[35][25];
    ele[35][3] != ele[35][26];
    ele[35][3] != ele[35][27];
    ele[35][3] != ele[35][28];
    ele[35][3] != ele[35][29];
    ele[35][3] != ele[35][30];
    ele[35][3] != ele[35][31];
    ele[35][3] != ele[35][32];
    ele[35][3] != ele[35][33];
    ele[35][3] != ele[35][34];
    ele[35][3] != ele[35][35];
    ele[35][3] != ele[35][4];
    ele[35][3] != ele[35][5];
    ele[35][3] != ele[35][6];
    ele[35][3] != ele[35][7];
    ele[35][3] != ele[35][8];
    ele[35][3] != ele[35][9];
    ele[35][30] != ele[35][31];
    ele[35][30] != ele[35][32];
    ele[35][30] != ele[35][33];
    ele[35][30] != ele[35][34];
    ele[35][30] != ele[35][35];
    ele[35][31] != ele[35][32];
    ele[35][31] != ele[35][33];
    ele[35][31] != ele[35][34];
    ele[35][31] != ele[35][35];
    ele[35][32] != ele[35][33];
    ele[35][32] != ele[35][34];
    ele[35][32] != ele[35][35];
    ele[35][33] != ele[35][34];
    ele[35][33] != ele[35][35];
    ele[35][34] != ele[35][35];
    ele[35][4] != ele[35][10];
    ele[35][4] != ele[35][11];
    ele[35][4] != ele[35][12];
    ele[35][4] != ele[35][13];
    ele[35][4] != ele[35][14];
    ele[35][4] != ele[35][15];
    ele[35][4] != ele[35][16];
    ele[35][4] != ele[35][17];
    ele[35][4] != ele[35][18];
    ele[35][4] != ele[35][19];
    ele[35][4] != ele[35][20];
    ele[35][4] != ele[35][21];
    ele[35][4] != ele[35][22];
    ele[35][4] != ele[35][23];
    ele[35][4] != ele[35][24];
    ele[35][4] != ele[35][25];
    ele[35][4] != ele[35][26];
    ele[35][4] != ele[35][27];
    ele[35][4] != ele[35][28];
    ele[35][4] != ele[35][29];
    ele[35][4] != ele[35][30];
    ele[35][4] != ele[35][31];
    ele[35][4] != ele[35][32];
    ele[35][4] != ele[35][33];
    ele[35][4] != ele[35][34];
    ele[35][4] != ele[35][35];
    ele[35][4] != ele[35][5];
    ele[35][4] != ele[35][6];
    ele[35][4] != ele[35][7];
    ele[35][4] != ele[35][8];
    ele[35][4] != ele[35][9];
    ele[35][5] != ele[35][10];
    ele[35][5] != ele[35][11];
    ele[35][5] != ele[35][12];
    ele[35][5] != ele[35][13];
    ele[35][5] != ele[35][14];
    ele[35][5] != ele[35][15];
    ele[35][5] != ele[35][16];
    ele[35][5] != ele[35][17];
    ele[35][5] != ele[35][18];
    ele[35][5] != ele[35][19];
    ele[35][5] != ele[35][20];
    ele[35][5] != ele[35][21];
    ele[35][5] != ele[35][22];
    ele[35][5] != ele[35][23];
    ele[35][5] != ele[35][24];
    ele[35][5] != ele[35][25];
    ele[35][5] != ele[35][26];
    ele[35][5] != ele[35][27];
    ele[35][5] != ele[35][28];
    ele[35][5] != ele[35][29];
    ele[35][5] != ele[35][30];
    ele[35][5] != ele[35][31];
    ele[35][5] != ele[35][32];
    ele[35][5] != ele[35][33];
    ele[35][5] != ele[35][34];
    ele[35][5] != ele[35][35];
    ele[35][5] != ele[35][6];
    ele[35][5] != ele[35][7];
    ele[35][5] != ele[35][8];
    ele[35][5] != ele[35][9];
    ele[35][6] != ele[35][10];
    ele[35][6] != ele[35][11];
    ele[35][6] != ele[35][12];
    ele[35][6] != ele[35][13];
    ele[35][6] != ele[35][14];
    ele[35][6] != ele[35][15];
    ele[35][6] != ele[35][16];
    ele[35][6] != ele[35][17];
    ele[35][6] != ele[35][18];
    ele[35][6] != ele[35][19];
    ele[35][6] != ele[35][20];
    ele[35][6] != ele[35][21];
    ele[35][6] != ele[35][22];
    ele[35][6] != ele[35][23];
    ele[35][6] != ele[35][24];
    ele[35][6] != ele[35][25];
    ele[35][6] != ele[35][26];
    ele[35][6] != ele[35][27];
    ele[35][6] != ele[35][28];
    ele[35][6] != ele[35][29];
    ele[35][6] != ele[35][30];
    ele[35][6] != ele[35][31];
    ele[35][6] != ele[35][32];
    ele[35][6] != ele[35][33];
    ele[35][6] != ele[35][34];
    ele[35][6] != ele[35][35];
    ele[35][6] != ele[35][7];
    ele[35][6] != ele[35][8];
    ele[35][6] != ele[35][9];
    ele[35][7] != ele[35][10];
    ele[35][7] != ele[35][11];
    ele[35][7] != ele[35][12];
    ele[35][7] != ele[35][13];
    ele[35][7] != ele[35][14];
    ele[35][7] != ele[35][15];
    ele[35][7] != ele[35][16];
    ele[35][7] != ele[35][17];
    ele[35][7] != ele[35][18];
    ele[35][7] != ele[35][19];
    ele[35][7] != ele[35][20];
    ele[35][7] != ele[35][21];
    ele[35][7] != ele[35][22];
    ele[35][7] != ele[35][23];
    ele[35][7] != ele[35][24];
    ele[35][7] != ele[35][25];
    ele[35][7] != ele[35][26];
    ele[35][7] != ele[35][27];
    ele[35][7] != ele[35][28];
    ele[35][7] != ele[35][29];
    ele[35][7] != ele[35][30];
    ele[35][7] != ele[35][31];
    ele[35][7] != ele[35][32];
    ele[35][7] != ele[35][33];
    ele[35][7] != ele[35][34];
    ele[35][7] != ele[35][35];
    ele[35][7] != ele[35][8];
    ele[35][7] != ele[35][9];
    ele[35][8] != ele[35][10];
    ele[35][8] != ele[35][11];
    ele[35][8] != ele[35][12];
    ele[35][8] != ele[35][13];
    ele[35][8] != ele[35][14];
    ele[35][8] != ele[35][15];
    ele[35][8] != ele[35][16];
    ele[35][8] != ele[35][17];
    ele[35][8] != ele[35][18];
    ele[35][8] != ele[35][19];
    ele[35][8] != ele[35][20];
    ele[35][8] != ele[35][21];
    ele[35][8] != ele[35][22];
    ele[35][8] != ele[35][23];
    ele[35][8] != ele[35][24];
    ele[35][8] != ele[35][25];
    ele[35][8] != ele[35][26];
    ele[35][8] != ele[35][27];
    ele[35][8] != ele[35][28];
    ele[35][8] != ele[35][29];
    ele[35][8] != ele[35][30];
    ele[35][8] != ele[35][31];
    ele[35][8] != ele[35][32];
    ele[35][8] != ele[35][33];
    ele[35][8] != ele[35][34];
    ele[35][8] != ele[35][35];
    ele[35][8] != ele[35][9];
    ele[35][9] != ele[35][10];
    ele[35][9] != ele[35][11];
    ele[35][9] != ele[35][12];
    ele[35][9] != ele[35][13];
    ele[35][9] != ele[35][14];
    ele[35][9] != ele[35][15];
    ele[35][9] != ele[35][16];
    ele[35][9] != ele[35][17];
    ele[35][9] != ele[35][18];
    ele[35][9] != ele[35][19];
    ele[35][9] != ele[35][20];
    ele[35][9] != ele[35][21];
    ele[35][9] != ele[35][22];
    ele[35][9] != ele[35][23];
    ele[35][9] != ele[35][24];
    ele[35][9] != ele[35][25];
    ele[35][9] != ele[35][26];
    ele[35][9] != ele[35][27];
    ele[35][9] != ele[35][28];
    ele[35][9] != ele[35][29];
    ele[35][9] != ele[35][30];
    ele[35][9] != ele[35][31];
    ele[35][9] != ele[35][32];
    ele[35][9] != ele[35][33];
    ele[35][9] != ele[35][34];
    ele[35][9] != ele[35][35];
    ele[4][0] != ele[10][0];
    ele[4][0] != ele[11][0];
    ele[4][0] != ele[12][0];
    ele[4][0] != ele[13][0];
    ele[4][0] != ele[14][0];
    ele[4][0] != ele[15][0];
    ele[4][0] != ele[16][0];
    ele[4][0] != ele[17][0];
    ele[4][0] != ele[18][0];
    ele[4][0] != ele[19][0];
    ele[4][0] != ele[20][0];
    ele[4][0] != ele[21][0];
    ele[4][0] != ele[22][0];
    ele[4][0] != ele[23][0];
    ele[4][0] != ele[24][0];
    ele[4][0] != ele[25][0];
    ele[4][0] != ele[26][0];
    ele[4][0] != ele[27][0];
    ele[4][0] != ele[28][0];
    ele[4][0] != ele[29][0];
    ele[4][0] != ele[30][0];
    ele[4][0] != ele[31][0];
    ele[4][0] != ele[32][0];
    ele[4][0] != ele[33][0];
    ele[4][0] != ele[34][0];
    ele[4][0] != ele[35][0];
    ele[4][0] != ele[4][1];
    ele[4][0] != ele[4][10];
    ele[4][0] != ele[4][11];
    ele[4][0] != ele[4][12];
    ele[4][0] != ele[4][13];
    ele[4][0] != ele[4][14];
    ele[4][0] != ele[4][15];
    ele[4][0] != ele[4][16];
    ele[4][0] != ele[4][17];
    ele[4][0] != ele[4][18];
    ele[4][0] != ele[4][19];
    ele[4][0] != ele[4][2];
    ele[4][0] != ele[4][20];
    ele[4][0] != ele[4][21];
    ele[4][0] != ele[4][22];
    ele[4][0] != ele[4][23];
    ele[4][0] != ele[4][24];
    ele[4][0] != ele[4][25];
    ele[4][0] != ele[4][26];
    ele[4][0] != ele[4][27];
    ele[4][0] != ele[4][28];
    ele[4][0] != ele[4][29];
    ele[4][0] != ele[4][3];
    ele[4][0] != ele[4][30];
    ele[4][0] != ele[4][31];
    ele[4][0] != ele[4][32];
    ele[4][0] != ele[4][33];
    ele[4][0] != ele[4][34];
    ele[4][0] != ele[4][35];
    ele[4][0] != ele[4][4];
    ele[4][0] != ele[4][5];
    ele[4][0] != ele[4][6];
    ele[4][0] != ele[4][7];
    ele[4][0] != ele[4][8];
    ele[4][0] != ele[4][9];
    ele[4][0] != ele[5][0];
    ele[4][0] != ele[5][1];
    ele[4][0] != ele[5][2];
    ele[4][0] != ele[5][3];
    ele[4][0] != ele[5][4];
    ele[4][0] != ele[5][5];
    ele[4][0] != ele[6][0];
    ele[4][0] != ele[7][0];
    ele[4][0] != ele[8][0];
    ele[4][0] != ele[9][0];
    ele[4][1] != ele[10][1];
    ele[4][1] != ele[11][1];
    ele[4][1] != ele[12][1];
    ele[4][1] != ele[13][1];
    ele[4][1] != ele[14][1];
    ele[4][1] != ele[15][1];
    ele[4][1] != ele[16][1];
    ele[4][1] != ele[17][1];
    ele[4][1] != ele[18][1];
    ele[4][1] != ele[19][1];
    ele[4][1] != ele[20][1];
    ele[4][1] != ele[21][1];
    ele[4][1] != ele[22][1];
    ele[4][1] != ele[23][1];
    ele[4][1] != ele[24][1];
    ele[4][1] != ele[25][1];
    ele[4][1] != ele[26][1];
    ele[4][1] != ele[27][1];
    ele[4][1] != ele[28][1];
    ele[4][1] != ele[29][1];
    ele[4][1] != ele[30][1];
    ele[4][1] != ele[31][1];
    ele[4][1] != ele[32][1];
    ele[4][1] != ele[33][1];
    ele[4][1] != ele[34][1];
    ele[4][1] != ele[35][1];
    ele[4][1] != ele[4][10];
    ele[4][1] != ele[4][11];
    ele[4][1] != ele[4][12];
    ele[4][1] != ele[4][13];
    ele[4][1] != ele[4][14];
    ele[4][1] != ele[4][15];
    ele[4][1] != ele[4][16];
    ele[4][1] != ele[4][17];
    ele[4][1] != ele[4][18];
    ele[4][1] != ele[4][19];
    ele[4][1] != ele[4][2];
    ele[4][1] != ele[4][20];
    ele[4][1] != ele[4][21];
    ele[4][1] != ele[4][22];
    ele[4][1] != ele[4][23];
    ele[4][1] != ele[4][24];
    ele[4][1] != ele[4][25];
    ele[4][1] != ele[4][26];
    ele[4][1] != ele[4][27];
    ele[4][1] != ele[4][28];
    ele[4][1] != ele[4][29];
    ele[4][1] != ele[4][3];
    ele[4][1] != ele[4][30];
    ele[4][1] != ele[4][31];
    ele[4][1] != ele[4][32];
    ele[4][1] != ele[4][33];
    ele[4][1] != ele[4][34];
    ele[4][1] != ele[4][35];
    ele[4][1] != ele[4][4];
    ele[4][1] != ele[4][5];
    ele[4][1] != ele[4][6];
    ele[4][1] != ele[4][7];
    ele[4][1] != ele[4][8];
    ele[4][1] != ele[4][9];
    ele[4][1] != ele[5][0];
    ele[4][1] != ele[5][1];
    ele[4][1] != ele[5][2];
    ele[4][1] != ele[5][3];
    ele[4][1] != ele[5][4];
    ele[4][1] != ele[5][5];
    ele[4][1] != ele[6][1];
    ele[4][1] != ele[7][1];
    ele[4][1] != ele[8][1];
    ele[4][1] != ele[9][1];
    ele[4][10] != ele[10][10];
    ele[4][10] != ele[11][10];
    ele[4][10] != ele[12][10];
    ele[4][10] != ele[13][10];
    ele[4][10] != ele[14][10];
    ele[4][10] != ele[15][10];
    ele[4][10] != ele[16][10];
    ele[4][10] != ele[17][10];
    ele[4][10] != ele[18][10];
    ele[4][10] != ele[19][10];
    ele[4][10] != ele[20][10];
    ele[4][10] != ele[21][10];
    ele[4][10] != ele[22][10];
    ele[4][10] != ele[23][10];
    ele[4][10] != ele[24][10];
    ele[4][10] != ele[25][10];
    ele[4][10] != ele[26][10];
    ele[4][10] != ele[27][10];
    ele[4][10] != ele[28][10];
    ele[4][10] != ele[29][10];
    ele[4][10] != ele[30][10];
    ele[4][10] != ele[31][10];
    ele[4][10] != ele[32][10];
    ele[4][10] != ele[33][10];
    ele[4][10] != ele[34][10];
    ele[4][10] != ele[35][10];
    ele[4][10] != ele[4][11];
    ele[4][10] != ele[4][12];
    ele[4][10] != ele[4][13];
    ele[4][10] != ele[4][14];
    ele[4][10] != ele[4][15];
    ele[4][10] != ele[4][16];
    ele[4][10] != ele[4][17];
    ele[4][10] != ele[4][18];
    ele[4][10] != ele[4][19];
    ele[4][10] != ele[4][20];
    ele[4][10] != ele[4][21];
    ele[4][10] != ele[4][22];
    ele[4][10] != ele[4][23];
    ele[4][10] != ele[4][24];
    ele[4][10] != ele[4][25];
    ele[4][10] != ele[4][26];
    ele[4][10] != ele[4][27];
    ele[4][10] != ele[4][28];
    ele[4][10] != ele[4][29];
    ele[4][10] != ele[4][30];
    ele[4][10] != ele[4][31];
    ele[4][10] != ele[4][32];
    ele[4][10] != ele[4][33];
    ele[4][10] != ele[4][34];
    ele[4][10] != ele[4][35];
    ele[4][10] != ele[5][10];
    ele[4][10] != ele[5][11];
    ele[4][10] != ele[5][6];
    ele[4][10] != ele[5][7];
    ele[4][10] != ele[5][8];
    ele[4][10] != ele[5][9];
    ele[4][10] != ele[6][10];
    ele[4][10] != ele[7][10];
    ele[4][10] != ele[8][10];
    ele[4][10] != ele[9][10];
    ele[4][11] != ele[10][11];
    ele[4][11] != ele[11][11];
    ele[4][11] != ele[12][11];
    ele[4][11] != ele[13][11];
    ele[4][11] != ele[14][11];
    ele[4][11] != ele[15][11];
    ele[4][11] != ele[16][11];
    ele[4][11] != ele[17][11];
    ele[4][11] != ele[18][11];
    ele[4][11] != ele[19][11];
    ele[4][11] != ele[20][11];
    ele[4][11] != ele[21][11];
    ele[4][11] != ele[22][11];
    ele[4][11] != ele[23][11];
    ele[4][11] != ele[24][11];
    ele[4][11] != ele[25][11];
    ele[4][11] != ele[26][11];
    ele[4][11] != ele[27][11];
    ele[4][11] != ele[28][11];
    ele[4][11] != ele[29][11];
    ele[4][11] != ele[30][11];
    ele[4][11] != ele[31][11];
    ele[4][11] != ele[32][11];
    ele[4][11] != ele[33][11];
    ele[4][11] != ele[34][11];
    ele[4][11] != ele[35][11];
    ele[4][11] != ele[4][12];
    ele[4][11] != ele[4][13];
    ele[4][11] != ele[4][14];
    ele[4][11] != ele[4][15];
    ele[4][11] != ele[4][16];
    ele[4][11] != ele[4][17];
    ele[4][11] != ele[4][18];
    ele[4][11] != ele[4][19];
    ele[4][11] != ele[4][20];
    ele[4][11] != ele[4][21];
    ele[4][11] != ele[4][22];
    ele[4][11] != ele[4][23];
    ele[4][11] != ele[4][24];
    ele[4][11] != ele[4][25];
    ele[4][11] != ele[4][26];
    ele[4][11] != ele[4][27];
    ele[4][11] != ele[4][28];
    ele[4][11] != ele[4][29];
    ele[4][11] != ele[4][30];
    ele[4][11] != ele[4][31];
    ele[4][11] != ele[4][32];
    ele[4][11] != ele[4][33];
    ele[4][11] != ele[4][34];
    ele[4][11] != ele[4][35];
    ele[4][11] != ele[5][10];
    ele[4][11] != ele[5][11];
    ele[4][11] != ele[5][6];
    ele[4][11] != ele[5][7];
    ele[4][11] != ele[5][8];
    ele[4][11] != ele[5][9];
    ele[4][11] != ele[6][11];
    ele[4][11] != ele[7][11];
    ele[4][11] != ele[8][11];
    ele[4][11] != ele[9][11];
    ele[4][12] != ele[10][12];
    ele[4][12] != ele[11][12];
    ele[4][12] != ele[12][12];
    ele[4][12] != ele[13][12];
    ele[4][12] != ele[14][12];
    ele[4][12] != ele[15][12];
    ele[4][12] != ele[16][12];
    ele[4][12] != ele[17][12];
    ele[4][12] != ele[18][12];
    ele[4][12] != ele[19][12];
    ele[4][12] != ele[20][12];
    ele[4][12] != ele[21][12];
    ele[4][12] != ele[22][12];
    ele[4][12] != ele[23][12];
    ele[4][12] != ele[24][12];
    ele[4][12] != ele[25][12];
    ele[4][12] != ele[26][12];
    ele[4][12] != ele[27][12];
    ele[4][12] != ele[28][12];
    ele[4][12] != ele[29][12];
    ele[4][12] != ele[30][12];
    ele[4][12] != ele[31][12];
    ele[4][12] != ele[32][12];
    ele[4][12] != ele[33][12];
    ele[4][12] != ele[34][12];
    ele[4][12] != ele[35][12];
    ele[4][12] != ele[4][13];
    ele[4][12] != ele[4][14];
    ele[4][12] != ele[4][15];
    ele[4][12] != ele[4][16];
    ele[4][12] != ele[4][17];
    ele[4][12] != ele[4][18];
    ele[4][12] != ele[4][19];
    ele[4][12] != ele[4][20];
    ele[4][12] != ele[4][21];
    ele[4][12] != ele[4][22];
    ele[4][12] != ele[4][23];
    ele[4][12] != ele[4][24];
    ele[4][12] != ele[4][25];
    ele[4][12] != ele[4][26];
    ele[4][12] != ele[4][27];
    ele[4][12] != ele[4][28];
    ele[4][12] != ele[4][29];
    ele[4][12] != ele[4][30];
    ele[4][12] != ele[4][31];
    ele[4][12] != ele[4][32];
    ele[4][12] != ele[4][33];
    ele[4][12] != ele[4][34];
    ele[4][12] != ele[4][35];
    ele[4][12] != ele[5][12];
    ele[4][12] != ele[5][13];
    ele[4][12] != ele[5][14];
    ele[4][12] != ele[5][15];
    ele[4][12] != ele[5][16];
    ele[4][12] != ele[5][17];
    ele[4][12] != ele[6][12];
    ele[4][12] != ele[7][12];
    ele[4][12] != ele[8][12];
    ele[4][12] != ele[9][12];
    ele[4][13] != ele[10][13];
    ele[4][13] != ele[11][13];
    ele[4][13] != ele[12][13];
    ele[4][13] != ele[13][13];
    ele[4][13] != ele[14][13];
    ele[4][13] != ele[15][13];
    ele[4][13] != ele[16][13];
    ele[4][13] != ele[17][13];
    ele[4][13] != ele[18][13];
    ele[4][13] != ele[19][13];
    ele[4][13] != ele[20][13];
    ele[4][13] != ele[21][13];
    ele[4][13] != ele[22][13];
    ele[4][13] != ele[23][13];
    ele[4][13] != ele[24][13];
    ele[4][13] != ele[25][13];
    ele[4][13] != ele[26][13];
    ele[4][13] != ele[27][13];
    ele[4][13] != ele[28][13];
    ele[4][13] != ele[29][13];
    ele[4][13] != ele[30][13];
    ele[4][13] != ele[31][13];
    ele[4][13] != ele[32][13];
    ele[4][13] != ele[33][13];
    ele[4][13] != ele[34][13];
    ele[4][13] != ele[35][13];
    ele[4][13] != ele[4][14];
    ele[4][13] != ele[4][15];
    ele[4][13] != ele[4][16];
    ele[4][13] != ele[4][17];
    ele[4][13] != ele[4][18];
    ele[4][13] != ele[4][19];
    ele[4][13] != ele[4][20];
    ele[4][13] != ele[4][21];
    ele[4][13] != ele[4][22];
    ele[4][13] != ele[4][23];
    ele[4][13] != ele[4][24];
    ele[4][13] != ele[4][25];
    ele[4][13] != ele[4][26];
    ele[4][13] != ele[4][27];
    ele[4][13] != ele[4][28];
    ele[4][13] != ele[4][29];
    ele[4][13] != ele[4][30];
    ele[4][13] != ele[4][31];
    ele[4][13] != ele[4][32];
    ele[4][13] != ele[4][33];
    ele[4][13] != ele[4][34];
    ele[4][13] != ele[4][35];
    ele[4][13] != ele[5][12];
    ele[4][13] != ele[5][13];
    ele[4][13] != ele[5][14];
    ele[4][13] != ele[5][15];
    ele[4][13] != ele[5][16];
    ele[4][13] != ele[5][17];
    ele[4][13] != ele[6][13];
    ele[4][13] != ele[7][13];
    ele[4][13] != ele[8][13];
    ele[4][13] != ele[9][13];
    ele[4][14] != ele[10][14];
    ele[4][14] != ele[11][14];
    ele[4][14] != ele[12][14];
    ele[4][14] != ele[13][14];
    ele[4][14] != ele[14][14];
    ele[4][14] != ele[15][14];
    ele[4][14] != ele[16][14];
    ele[4][14] != ele[17][14];
    ele[4][14] != ele[18][14];
    ele[4][14] != ele[19][14];
    ele[4][14] != ele[20][14];
    ele[4][14] != ele[21][14];
    ele[4][14] != ele[22][14];
    ele[4][14] != ele[23][14];
    ele[4][14] != ele[24][14];
    ele[4][14] != ele[25][14];
    ele[4][14] != ele[26][14];
    ele[4][14] != ele[27][14];
    ele[4][14] != ele[28][14];
    ele[4][14] != ele[29][14];
    ele[4][14] != ele[30][14];
    ele[4][14] != ele[31][14];
    ele[4][14] != ele[32][14];
    ele[4][14] != ele[33][14];
    ele[4][14] != ele[34][14];
    ele[4][14] != ele[35][14];
    ele[4][14] != ele[4][15];
    ele[4][14] != ele[4][16];
    ele[4][14] != ele[4][17];
    ele[4][14] != ele[4][18];
    ele[4][14] != ele[4][19];
    ele[4][14] != ele[4][20];
    ele[4][14] != ele[4][21];
    ele[4][14] != ele[4][22];
    ele[4][14] != ele[4][23];
    ele[4][14] != ele[4][24];
    ele[4][14] != ele[4][25];
    ele[4][14] != ele[4][26];
    ele[4][14] != ele[4][27];
    ele[4][14] != ele[4][28];
    ele[4][14] != ele[4][29];
    ele[4][14] != ele[4][30];
    ele[4][14] != ele[4][31];
    ele[4][14] != ele[4][32];
    ele[4][14] != ele[4][33];
    ele[4][14] != ele[4][34];
    ele[4][14] != ele[4][35];
    ele[4][14] != ele[5][12];
    ele[4][14] != ele[5][13];
    ele[4][14] != ele[5][14];
    ele[4][14] != ele[5][15];
    ele[4][14] != ele[5][16];
    ele[4][14] != ele[5][17];
    ele[4][14] != ele[6][14];
    ele[4][14] != ele[7][14];
    ele[4][14] != ele[8][14];
    ele[4][14] != ele[9][14];
    ele[4][15] != ele[10][15];
    ele[4][15] != ele[11][15];
    ele[4][15] != ele[12][15];
    ele[4][15] != ele[13][15];
    ele[4][15] != ele[14][15];
    ele[4][15] != ele[15][15];
    ele[4][15] != ele[16][15];
    ele[4][15] != ele[17][15];
    ele[4][15] != ele[18][15];
    ele[4][15] != ele[19][15];
    ele[4][15] != ele[20][15];
    ele[4][15] != ele[21][15];
    ele[4][15] != ele[22][15];
    ele[4][15] != ele[23][15];
    ele[4][15] != ele[24][15];
    ele[4][15] != ele[25][15];
    ele[4][15] != ele[26][15];
    ele[4][15] != ele[27][15];
    ele[4][15] != ele[28][15];
    ele[4][15] != ele[29][15];
    ele[4][15] != ele[30][15];
    ele[4][15] != ele[31][15];
    ele[4][15] != ele[32][15];
    ele[4][15] != ele[33][15];
    ele[4][15] != ele[34][15];
    ele[4][15] != ele[35][15];
    ele[4][15] != ele[4][16];
    ele[4][15] != ele[4][17];
    ele[4][15] != ele[4][18];
    ele[4][15] != ele[4][19];
    ele[4][15] != ele[4][20];
    ele[4][15] != ele[4][21];
    ele[4][15] != ele[4][22];
    ele[4][15] != ele[4][23];
    ele[4][15] != ele[4][24];
    ele[4][15] != ele[4][25];
    ele[4][15] != ele[4][26];
    ele[4][15] != ele[4][27];
    ele[4][15] != ele[4][28];
    ele[4][15] != ele[4][29];
    ele[4][15] != ele[4][30];
    ele[4][15] != ele[4][31];
    ele[4][15] != ele[4][32];
    ele[4][15] != ele[4][33];
    ele[4][15] != ele[4][34];
    ele[4][15] != ele[4][35];
    ele[4][15] != ele[5][12];
    ele[4][15] != ele[5][13];
    ele[4][15] != ele[5][14];
    ele[4][15] != ele[5][15];
    ele[4][15] != ele[5][16];
    ele[4][15] != ele[5][17];
    ele[4][15] != ele[6][15];
    ele[4][15] != ele[7][15];
    ele[4][15] != ele[8][15];
    ele[4][15] != ele[9][15];
    ele[4][16] != ele[10][16];
    ele[4][16] != ele[11][16];
    ele[4][16] != ele[12][16];
    ele[4][16] != ele[13][16];
    ele[4][16] != ele[14][16];
    ele[4][16] != ele[15][16];
    ele[4][16] != ele[16][16];
    ele[4][16] != ele[17][16];
    ele[4][16] != ele[18][16];
    ele[4][16] != ele[19][16];
    ele[4][16] != ele[20][16];
    ele[4][16] != ele[21][16];
    ele[4][16] != ele[22][16];
    ele[4][16] != ele[23][16];
    ele[4][16] != ele[24][16];
    ele[4][16] != ele[25][16];
    ele[4][16] != ele[26][16];
    ele[4][16] != ele[27][16];
    ele[4][16] != ele[28][16];
    ele[4][16] != ele[29][16];
    ele[4][16] != ele[30][16];
    ele[4][16] != ele[31][16];
    ele[4][16] != ele[32][16];
    ele[4][16] != ele[33][16];
    ele[4][16] != ele[34][16];
    ele[4][16] != ele[35][16];
    ele[4][16] != ele[4][17];
    ele[4][16] != ele[4][18];
    ele[4][16] != ele[4][19];
    ele[4][16] != ele[4][20];
    ele[4][16] != ele[4][21];
    ele[4][16] != ele[4][22];
    ele[4][16] != ele[4][23];
    ele[4][16] != ele[4][24];
    ele[4][16] != ele[4][25];
    ele[4][16] != ele[4][26];
    ele[4][16] != ele[4][27];
    ele[4][16] != ele[4][28];
    ele[4][16] != ele[4][29];
    ele[4][16] != ele[4][30];
    ele[4][16] != ele[4][31];
    ele[4][16] != ele[4][32];
    ele[4][16] != ele[4][33];
    ele[4][16] != ele[4][34];
    ele[4][16] != ele[4][35];
    ele[4][16] != ele[5][12];
    ele[4][16] != ele[5][13];
    ele[4][16] != ele[5][14];
    ele[4][16] != ele[5][15];
    ele[4][16] != ele[5][16];
    ele[4][16] != ele[5][17];
    ele[4][16] != ele[6][16];
    ele[4][16] != ele[7][16];
    ele[4][16] != ele[8][16];
    ele[4][16] != ele[9][16];
    ele[4][17] != ele[10][17];
    ele[4][17] != ele[11][17];
    ele[4][17] != ele[12][17];
    ele[4][17] != ele[13][17];
    ele[4][17] != ele[14][17];
    ele[4][17] != ele[15][17];
    ele[4][17] != ele[16][17];
    ele[4][17] != ele[17][17];
    ele[4][17] != ele[18][17];
    ele[4][17] != ele[19][17];
    ele[4][17] != ele[20][17];
    ele[4][17] != ele[21][17];
    ele[4][17] != ele[22][17];
    ele[4][17] != ele[23][17];
    ele[4][17] != ele[24][17];
    ele[4][17] != ele[25][17];
    ele[4][17] != ele[26][17];
    ele[4][17] != ele[27][17];
    ele[4][17] != ele[28][17];
    ele[4][17] != ele[29][17];
    ele[4][17] != ele[30][17];
    ele[4][17] != ele[31][17];
    ele[4][17] != ele[32][17];
    ele[4][17] != ele[33][17];
    ele[4][17] != ele[34][17];
    ele[4][17] != ele[35][17];
    ele[4][17] != ele[4][18];
    ele[4][17] != ele[4][19];
    ele[4][17] != ele[4][20];
    ele[4][17] != ele[4][21];
    ele[4][17] != ele[4][22];
    ele[4][17] != ele[4][23];
    ele[4][17] != ele[4][24];
    ele[4][17] != ele[4][25];
    ele[4][17] != ele[4][26];
    ele[4][17] != ele[4][27];
    ele[4][17] != ele[4][28];
    ele[4][17] != ele[4][29];
    ele[4][17] != ele[4][30];
    ele[4][17] != ele[4][31];
    ele[4][17] != ele[4][32];
    ele[4][17] != ele[4][33];
    ele[4][17] != ele[4][34];
    ele[4][17] != ele[4][35];
    ele[4][17] != ele[5][12];
    ele[4][17] != ele[5][13];
    ele[4][17] != ele[5][14];
    ele[4][17] != ele[5][15];
    ele[4][17] != ele[5][16];
    ele[4][17] != ele[5][17];
    ele[4][17] != ele[6][17];
    ele[4][17] != ele[7][17];
    ele[4][17] != ele[8][17];
    ele[4][17] != ele[9][17];
    ele[4][18] != ele[10][18];
    ele[4][18] != ele[11][18];
    ele[4][18] != ele[12][18];
    ele[4][18] != ele[13][18];
    ele[4][18] != ele[14][18];
    ele[4][18] != ele[15][18];
    ele[4][18] != ele[16][18];
    ele[4][18] != ele[17][18];
    ele[4][18] != ele[18][18];
    ele[4][18] != ele[19][18];
    ele[4][18] != ele[20][18];
    ele[4][18] != ele[21][18];
    ele[4][18] != ele[22][18];
    ele[4][18] != ele[23][18];
    ele[4][18] != ele[24][18];
    ele[4][18] != ele[25][18];
    ele[4][18] != ele[26][18];
    ele[4][18] != ele[27][18];
    ele[4][18] != ele[28][18];
    ele[4][18] != ele[29][18];
    ele[4][18] != ele[30][18];
    ele[4][18] != ele[31][18];
    ele[4][18] != ele[32][18];
    ele[4][18] != ele[33][18];
    ele[4][18] != ele[34][18];
    ele[4][18] != ele[35][18];
    ele[4][18] != ele[4][19];
    ele[4][18] != ele[4][20];
    ele[4][18] != ele[4][21];
    ele[4][18] != ele[4][22];
    ele[4][18] != ele[4][23];
    ele[4][18] != ele[4][24];
    ele[4][18] != ele[4][25];
    ele[4][18] != ele[4][26];
    ele[4][18] != ele[4][27];
    ele[4][18] != ele[4][28];
    ele[4][18] != ele[4][29];
    ele[4][18] != ele[4][30];
    ele[4][18] != ele[4][31];
    ele[4][18] != ele[4][32];
    ele[4][18] != ele[4][33];
    ele[4][18] != ele[4][34];
    ele[4][18] != ele[4][35];
    ele[4][18] != ele[5][18];
    ele[4][18] != ele[5][19];
    ele[4][18] != ele[5][20];
    ele[4][18] != ele[5][21];
    ele[4][18] != ele[5][22];
    ele[4][18] != ele[5][23];
    ele[4][18] != ele[6][18];
    ele[4][18] != ele[7][18];
    ele[4][18] != ele[8][18];
    ele[4][18] != ele[9][18];
    ele[4][19] != ele[10][19];
    ele[4][19] != ele[11][19];
    ele[4][19] != ele[12][19];
    ele[4][19] != ele[13][19];
    ele[4][19] != ele[14][19];
    ele[4][19] != ele[15][19];
    ele[4][19] != ele[16][19];
    ele[4][19] != ele[17][19];
    ele[4][19] != ele[18][19];
    ele[4][19] != ele[19][19];
    ele[4][19] != ele[20][19];
    ele[4][19] != ele[21][19];
    ele[4][19] != ele[22][19];
    ele[4][19] != ele[23][19];
    ele[4][19] != ele[24][19];
    ele[4][19] != ele[25][19];
    ele[4][19] != ele[26][19];
    ele[4][19] != ele[27][19];
    ele[4][19] != ele[28][19];
    ele[4][19] != ele[29][19];
    ele[4][19] != ele[30][19];
    ele[4][19] != ele[31][19];
    ele[4][19] != ele[32][19];
    ele[4][19] != ele[33][19];
    ele[4][19] != ele[34][19];
    ele[4][19] != ele[35][19];
    ele[4][19] != ele[4][20];
    ele[4][19] != ele[4][21];
    ele[4][19] != ele[4][22];
    ele[4][19] != ele[4][23];
    ele[4][19] != ele[4][24];
    ele[4][19] != ele[4][25];
    ele[4][19] != ele[4][26];
    ele[4][19] != ele[4][27];
    ele[4][19] != ele[4][28];
    ele[4][19] != ele[4][29];
    ele[4][19] != ele[4][30];
    ele[4][19] != ele[4][31];
    ele[4][19] != ele[4][32];
    ele[4][19] != ele[4][33];
    ele[4][19] != ele[4][34];
    ele[4][19] != ele[4][35];
    ele[4][19] != ele[5][18];
    ele[4][19] != ele[5][19];
    ele[4][19] != ele[5][20];
    ele[4][19] != ele[5][21];
    ele[4][19] != ele[5][22];
    ele[4][19] != ele[5][23];
    ele[4][19] != ele[6][19];
    ele[4][19] != ele[7][19];
    ele[4][19] != ele[8][19];
    ele[4][19] != ele[9][19];
    ele[4][2] != ele[10][2];
    ele[4][2] != ele[11][2];
    ele[4][2] != ele[12][2];
    ele[4][2] != ele[13][2];
    ele[4][2] != ele[14][2];
    ele[4][2] != ele[15][2];
    ele[4][2] != ele[16][2];
    ele[4][2] != ele[17][2];
    ele[4][2] != ele[18][2];
    ele[4][2] != ele[19][2];
    ele[4][2] != ele[20][2];
    ele[4][2] != ele[21][2];
    ele[4][2] != ele[22][2];
    ele[4][2] != ele[23][2];
    ele[4][2] != ele[24][2];
    ele[4][2] != ele[25][2];
    ele[4][2] != ele[26][2];
    ele[4][2] != ele[27][2];
    ele[4][2] != ele[28][2];
    ele[4][2] != ele[29][2];
    ele[4][2] != ele[30][2];
    ele[4][2] != ele[31][2];
    ele[4][2] != ele[32][2];
    ele[4][2] != ele[33][2];
    ele[4][2] != ele[34][2];
    ele[4][2] != ele[35][2];
    ele[4][2] != ele[4][10];
    ele[4][2] != ele[4][11];
    ele[4][2] != ele[4][12];
    ele[4][2] != ele[4][13];
    ele[4][2] != ele[4][14];
    ele[4][2] != ele[4][15];
    ele[4][2] != ele[4][16];
    ele[4][2] != ele[4][17];
    ele[4][2] != ele[4][18];
    ele[4][2] != ele[4][19];
    ele[4][2] != ele[4][20];
    ele[4][2] != ele[4][21];
    ele[4][2] != ele[4][22];
    ele[4][2] != ele[4][23];
    ele[4][2] != ele[4][24];
    ele[4][2] != ele[4][25];
    ele[4][2] != ele[4][26];
    ele[4][2] != ele[4][27];
    ele[4][2] != ele[4][28];
    ele[4][2] != ele[4][29];
    ele[4][2] != ele[4][3];
    ele[4][2] != ele[4][30];
    ele[4][2] != ele[4][31];
    ele[4][2] != ele[4][32];
    ele[4][2] != ele[4][33];
    ele[4][2] != ele[4][34];
    ele[4][2] != ele[4][35];
    ele[4][2] != ele[4][4];
    ele[4][2] != ele[4][5];
    ele[4][2] != ele[4][6];
    ele[4][2] != ele[4][7];
    ele[4][2] != ele[4][8];
    ele[4][2] != ele[4][9];
    ele[4][2] != ele[5][0];
    ele[4][2] != ele[5][1];
    ele[4][2] != ele[5][2];
    ele[4][2] != ele[5][3];
    ele[4][2] != ele[5][4];
    ele[4][2] != ele[5][5];
    ele[4][2] != ele[6][2];
    ele[4][2] != ele[7][2];
    ele[4][2] != ele[8][2];
    ele[4][2] != ele[9][2];
    ele[4][20] != ele[10][20];
    ele[4][20] != ele[11][20];
    ele[4][20] != ele[12][20];
    ele[4][20] != ele[13][20];
    ele[4][20] != ele[14][20];
    ele[4][20] != ele[15][20];
    ele[4][20] != ele[16][20];
    ele[4][20] != ele[17][20];
    ele[4][20] != ele[18][20];
    ele[4][20] != ele[19][20];
    ele[4][20] != ele[20][20];
    ele[4][20] != ele[21][20];
    ele[4][20] != ele[22][20];
    ele[4][20] != ele[23][20];
    ele[4][20] != ele[24][20];
    ele[4][20] != ele[25][20];
    ele[4][20] != ele[26][20];
    ele[4][20] != ele[27][20];
    ele[4][20] != ele[28][20];
    ele[4][20] != ele[29][20];
    ele[4][20] != ele[30][20];
    ele[4][20] != ele[31][20];
    ele[4][20] != ele[32][20];
    ele[4][20] != ele[33][20];
    ele[4][20] != ele[34][20];
    ele[4][20] != ele[35][20];
    ele[4][20] != ele[4][21];
    ele[4][20] != ele[4][22];
    ele[4][20] != ele[4][23];
    ele[4][20] != ele[4][24];
    ele[4][20] != ele[4][25];
    ele[4][20] != ele[4][26];
    ele[4][20] != ele[4][27];
    ele[4][20] != ele[4][28];
    ele[4][20] != ele[4][29];
    ele[4][20] != ele[4][30];
    ele[4][20] != ele[4][31];
    ele[4][20] != ele[4][32];
    ele[4][20] != ele[4][33];
    ele[4][20] != ele[4][34];
    ele[4][20] != ele[4][35];
    ele[4][20] != ele[5][18];
    ele[4][20] != ele[5][19];
    ele[4][20] != ele[5][20];
    ele[4][20] != ele[5][21];
    ele[4][20] != ele[5][22];
    ele[4][20] != ele[5][23];
    ele[4][20] != ele[6][20];
    ele[4][20] != ele[7][20];
    ele[4][20] != ele[8][20];
    ele[4][20] != ele[9][20];
    ele[4][21] != ele[10][21];
    ele[4][21] != ele[11][21];
    ele[4][21] != ele[12][21];
    ele[4][21] != ele[13][21];
    ele[4][21] != ele[14][21];
    ele[4][21] != ele[15][21];
    ele[4][21] != ele[16][21];
    ele[4][21] != ele[17][21];
    ele[4][21] != ele[18][21];
    ele[4][21] != ele[19][21];
    ele[4][21] != ele[20][21];
    ele[4][21] != ele[21][21];
    ele[4][21] != ele[22][21];
    ele[4][21] != ele[23][21];
    ele[4][21] != ele[24][21];
    ele[4][21] != ele[25][21];
    ele[4][21] != ele[26][21];
    ele[4][21] != ele[27][21];
    ele[4][21] != ele[28][21];
    ele[4][21] != ele[29][21];
    ele[4][21] != ele[30][21];
    ele[4][21] != ele[31][21];
    ele[4][21] != ele[32][21];
    ele[4][21] != ele[33][21];
    ele[4][21] != ele[34][21];
    ele[4][21] != ele[35][21];
    ele[4][21] != ele[4][22];
    ele[4][21] != ele[4][23];
    ele[4][21] != ele[4][24];
    ele[4][21] != ele[4][25];
    ele[4][21] != ele[4][26];
    ele[4][21] != ele[4][27];
    ele[4][21] != ele[4][28];
    ele[4][21] != ele[4][29];
    ele[4][21] != ele[4][30];
    ele[4][21] != ele[4][31];
    ele[4][21] != ele[4][32];
    ele[4][21] != ele[4][33];
    ele[4][21] != ele[4][34];
    ele[4][21] != ele[4][35];
    ele[4][21] != ele[5][18];
    ele[4][21] != ele[5][19];
    ele[4][21] != ele[5][20];
    ele[4][21] != ele[5][21];
    ele[4][21] != ele[5][22];
    ele[4][21] != ele[5][23];
    ele[4][21] != ele[6][21];
    ele[4][21] != ele[7][21];
    ele[4][21] != ele[8][21];
    ele[4][21] != ele[9][21];
    ele[4][22] != ele[10][22];
    ele[4][22] != ele[11][22];
    ele[4][22] != ele[12][22];
    ele[4][22] != ele[13][22];
    ele[4][22] != ele[14][22];
    ele[4][22] != ele[15][22];
    ele[4][22] != ele[16][22];
    ele[4][22] != ele[17][22];
    ele[4][22] != ele[18][22];
    ele[4][22] != ele[19][22];
    ele[4][22] != ele[20][22];
    ele[4][22] != ele[21][22];
    ele[4][22] != ele[22][22];
    ele[4][22] != ele[23][22];
    ele[4][22] != ele[24][22];
    ele[4][22] != ele[25][22];
    ele[4][22] != ele[26][22];
    ele[4][22] != ele[27][22];
    ele[4][22] != ele[28][22];
    ele[4][22] != ele[29][22];
    ele[4][22] != ele[30][22];
    ele[4][22] != ele[31][22];
    ele[4][22] != ele[32][22];
    ele[4][22] != ele[33][22];
    ele[4][22] != ele[34][22];
    ele[4][22] != ele[35][22];
    ele[4][22] != ele[4][23];
    ele[4][22] != ele[4][24];
    ele[4][22] != ele[4][25];
    ele[4][22] != ele[4][26];
    ele[4][22] != ele[4][27];
    ele[4][22] != ele[4][28];
    ele[4][22] != ele[4][29];
    ele[4][22] != ele[4][30];
    ele[4][22] != ele[4][31];
    ele[4][22] != ele[4][32];
    ele[4][22] != ele[4][33];
    ele[4][22] != ele[4][34];
    ele[4][22] != ele[4][35];
    ele[4][22] != ele[5][18];
    ele[4][22] != ele[5][19];
    ele[4][22] != ele[5][20];
    ele[4][22] != ele[5][21];
    ele[4][22] != ele[5][22];
    ele[4][22] != ele[5][23];
    ele[4][22] != ele[6][22];
    ele[4][22] != ele[7][22];
    ele[4][22] != ele[8][22];
    ele[4][22] != ele[9][22];
    ele[4][23] != ele[10][23];
    ele[4][23] != ele[11][23];
    ele[4][23] != ele[12][23];
    ele[4][23] != ele[13][23];
    ele[4][23] != ele[14][23];
    ele[4][23] != ele[15][23];
    ele[4][23] != ele[16][23];
    ele[4][23] != ele[17][23];
    ele[4][23] != ele[18][23];
    ele[4][23] != ele[19][23];
    ele[4][23] != ele[20][23];
    ele[4][23] != ele[21][23];
    ele[4][23] != ele[22][23];
    ele[4][23] != ele[23][23];
    ele[4][23] != ele[24][23];
    ele[4][23] != ele[25][23];
    ele[4][23] != ele[26][23];
    ele[4][23] != ele[27][23];
    ele[4][23] != ele[28][23];
    ele[4][23] != ele[29][23];
    ele[4][23] != ele[30][23];
    ele[4][23] != ele[31][23];
    ele[4][23] != ele[32][23];
    ele[4][23] != ele[33][23];
    ele[4][23] != ele[34][23];
    ele[4][23] != ele[35][23];
    ele[4][23] != ele[4][24];
    ele[4][23] != ele[4][25];
    ele[4][23] != ele[4][26];
    ele[4][23] != ele[4][27];
    ele[4][23] != ele[4][28];
    ele[4][23] != ele[4][29];
    ele[4][23] != ele[4][30];
    ele[4][23] != ele[4][31];
    ele[4][23] != ele[4][32];
    ele[4][23] != ele[4][33];
    ele[4][23] != ele[4][34];
    ele[4][23] != ele[4][35];
    ele[4][23] != ele[5][18];
    ele[4][23] != ele[5][19];
    ele[4][23] != ele[5][20];
    ele[4][23] != ele[5][21];
    ele[4][23] != ele[5][22];
    ele[4][23] != ele[5][23];
    ele[4][23] != ele[6][23];
    ele[4][23] != ele[7][23];
    ele[4][23] != ele[8][23];
    ele[4][23] != ele[9][23];
    ele[4][24] != ele[10][24];
    ele[4][24] != ele[11][24];
    ele[4][24] != ele[12][24];
    ele[4][24] != ele[13][24];
    ele[4][24] != ele[14][24];
    ele[4][24] != ele[15][24];
    ele[4][24] != ele[16][24];
    ele[4][24] != ele[17][24];
    ele[4][24] != ele[18][24];
    ele[4][24] != ele[19][24];
    ele[4][24] != ele[20][24];
    ele[4][24] != ele[21][24];
    ele[4][24] != ele[22][24];
    ele[4][24] != ele[23][24];
    ele[4][24] != ele[24][24];
    ele[4][24] != ele[25][24];
    ele[4][24] != ele[26][24];
    ele[4][24] != ele[27][24];
    ele[4][24] != ele[28][24];
    ele[4][24] != ele[29][24];
    ele[4][24] != ele[30][24];
    ele[4][24] != ele[31][24];
    ele[4][24] != ele[32][24];
    ele[4][24] != ele[33][24];
    ele[4][24] != ele[34][24];
    ele[4][24] != ele[35][24];
    ele[4][24] != ele[4][25];
    ele[4][24] != ele[4][26];
    ele[4][24] != ele[4][27];
    ele[4][24] != ele[4][28];
    ele[4][24] != ele[4][29];
    ele[4][24] != ele[4][30];
    ele[4][24] != ele[4][31];
    ele[4][24] != ele[4][32];
    ele[4][24] != ele[4][33];
    ele[4][24] != ele[4][34];
    ele[4][24] != ele[4][35];
    ele[4][24] != ele[5][24];
    ele[4][24] != ele[5][25];
    ele[4][24] != ele[5][26];
    ele[4][24] != ele[5][27];
    ele[4][24] != ele[5][28];
    ele[4][24] != ele[5][29];
    ele[4][24] != ele[6][24];
    ele[4][24] != ele[7][24];
    ele[4][24] != ele[8][24];
    ele[4][24] != ele[9][24];
    ele[4][25] != ele[10][25];
    ele[4][25] != ele[11][25];
    ele[4][25] != ele[12][25];
    ele[4][25] != ele[13][25];
    ele[4][25] != ele[14][25];
    ele[4][25] != ele[15][25];
    ele[4][25] != ele[16][25];
    ele[4][25] != ele[17][25];
    ele[4][25] != ele[18][25];
    ele[4][25] != ele[19][25];
    ele[4][25] != ele[20][25];
    ele[4][25] != ele[21][25];
    ele[4][25] != ele[22][25];
    ele[4][25] != ele[23][25];
    ele[4][25] != ele[24][25];
    ele[4][25] != ele[25][25];
    ele[4][25] != ele[26][25];
    ele[4][25] != ele[27][25];
    ele[4][25] != ele[28][25];
    ele[4][25] != ele[29][25];
    ele[4][25] != ele[30][25];
    ele[4][25] != ele[31][25];
    ele[4][25] != ele[32][25];
    ele[4][25] != ele[33][25];
    ele[4][25] != ele[34][25];
    ele[4][25] != ele[35][25];
    ele[4][25] != ele[4][26];
    ele[4][25] != ele[4][27];
    ele[4][25] != ele[4][28];
    ele[4][25] != ele[4][29];
    ele[4][25] != ele[4][30];
    ele[4][25] != ele[4][31];
    ele[4][25] != ele[4][32];
    ele[4][25] != ele[4][33];
    ele[4][25] != ele[4][34];
    ele[4][25] != ele[4][35];
    ele[4][25] != ele[5][24];
    ele[4][25] != ele[5][25];
    ele[4][25] != ele[5][26];
    ele[4][25] != ele[5][27];
    ele[4][25] != ele[5][28];
    ele[4][25] != ele[5][29];
    ele[4][25] != ele[6][25];
    ele[4][25] != ele[7][25];
    ele[4][25] != ele[8][25];
    ele[4][25] != ele[9][25];
    ele[4][26] != ele[10][26];
    ele[4][26] != ele[11][26];
    ele[4][26] != ele[12][26];
    ele[4][26] != ele[13][26];
    ele[4][26] != ele[14][26];
    ele[4][26] != ele[15][26];
    ele[4][26] != ele[16][26];
    ele[4][26] != ele[17][26];
    ele[4][26] != ele[18][26];
    ele[4][26] != ele[19][26];
    ele[4][26] != ele[20][26];
    ele[4][26] != ele[21][26];
    ele[4][26] != ele[22][26];
    ele[4][26] != ele[23][26];
    ele[4][26] != ele[24][26];
    ele[4][26] != ele[25][26];
    ele[4][26] != ele[26][26];
    ele[4][26] != ele[27][26];
    ele[4][26] != ele[28][26];
    ele[4][26] != ele[29][26];
    ele[4][26] != ele[30][26];
    ele[4][26] != ele[31][26];
    ele[4][26] != ele[32][26];
    ele[4][26] != ele[33][26];
    ele[4][26] != ele[34][26];
    ele[4][26] != ele[35][26];
    ele[4][26] != ele[4][27];
    ele[4][26] != ele[4][28];
    ele[4][26] != ele[4][29];
    ele[4][26] != ele[4][30];
    ele[4][26] != ele[4][31];
    ele[4][26] != ele[4][32];
    ele[4][26] != ele[4][33];
    ele[4][26] != ele[4][34];
    ele[4][26] != ele[4][35];
    ele[4][26] != ele[5][24];
    ele[4][26] != ele[5][25];
    ele[4][26] != ele[5][26];
    ele[4][26] != ele[5][27];
    ele[4][26] != ele[5][28];
    ele[4][26] != ele[5][29];
    ele[4][26] != ele[6][26];
    ele[4][26] != ele[7][26];
    ele[4][26] != ele[8][26];
    ele[4][26] != ele[9][26];
    ele[4][27] != ele[10][27];
    ele[4][27] != ele[11][27];
    ele[4][27] != ele[12][27];
    ele[4][27] != ele[13][27];
    ele[4][27] != ele[14][27];
    ele[4][27] != ele[15][27];
    ele[4][27] != ele[16][27];
    ele[4][27] != ele[17][27];
    ele[4][27] != ele[18][27];
    ele[4][27] != ele[19][27];
    ele[4][27] != ele[20][27];
    ele[4][27] != ele[21][27];
    ele[4][27] != ele[22][27];
    ele[4][27] != ele[23][27];
    ele[4][27] != ele[24][27];
    ele[4][27] != ele[25][27];
    ele[4][27] != ele[26][27];
    ele[4][27] != ele[27][27];
    ele[4][27] != ele[28][27];
    ele[4][27] != ele[29][27];
    ele[4][27] != ele[30][27];
    ele[4][27] != ele[31][27];
    ele[4][27] != ele[32][27];
    ele[4][27] != ele[33][27];
    ele[4][27] != ele[34][27];
    ele[4][27] != ele[35][27];
    ele[4][27] != ele[4][28];
    ele[4][27] != ele[4][29];
    ele[4][27] != ele[4][30];
    ele[4][27] != ele[4][31];
    ele[4][27] != ele[4][32];
    ele[4][27] != ele[4][33];
    ele[4][27] != ele[4][34];
    ele[4][27] != ele[4][35];
    ele[4][27] != ele[5][24];
    ele[4][27] != ele[5][25];
    ele[4][27] != ele[5][26];
    ele[4][27] != ele[5][27];
    ele[4][27] != ele[5][28];
    ele[4][27] != ele[5][29];
    ele[4][27] != ele[6][27];
    ele[4][27] != ele[7][27];
    ele[4][27] != ele[8][27];
    ele[4][27] != ele[9][27];
    ele[4][28] != ele[10][28];
    ele[4][28] != ele[11][28];
    ele[4][28] != ele[12][28];
    ele[4][28] != ele[13][28];
    ele[4][28] != ele[14][28];
    ele[4][28] != ele[15][28];
    ele[4][28] != ele[16][28];
    ele[4][28] != ele[17][28];
    ele[4][28] != ele[18][28];
    ele[4][28] != ele[19][28];
    ele[4][28] != ele[20][28];
    ele[4][28] != ele[21][28];
    ele[4][28] != ele[22][28];
    ele[4][28] != ele[23][28];
    ele[4][28] != ele[24][28];
    ele[4][28] != ele[25][28];
    ele[4][28] != ele[26][28];
    ele[4][28] != ele[27][28];
    ele[4][28] != ele[28][28];
    ele[4][28] != ele[29][28];
    ele[4][28] != ele[30][28];
    ele[4][28] != ele[31][28];
    ele[4][28] != ele[32][28];
    ele[4][28] != ele[33][28];
    ele[4][28] != ele[34][28];
    ele[4][28] != ele[35][28];
    ele[4][28] != ele[4][29];
    ele[4][28] != ele[4][30];
    ele[4][28] != ele[4][31];
    ele[4][28] != ele[4][32];
    ele[4][28] != ele[4][33];
    ele[4][28] != ele[4][34];
    ele[4][28] != ele[4][35];
    ele[4][28] != ele[5][24];
    ele[4][28] != ele[5][25];
    ele[4][28] != ele[5][26];
    ele[4][28] != ele[5][27];
    ele[4][28] != ele[5][28];
    ele[4][28] != ele[5][29];
    ele[4][28] != ele[6][28];
    ele[4][28] != ele[7][28];
    ele[4][28] != ele[8][28];
    ele[4][28] != ele[9][28];
    ele[4][29] != ele[10][29];
    ele[4][29] != ele[11][29];
    ele[4][29] != ele[12][29];
    ele[4][29] != ele[13][29];
    ele[4][29] != ele[14][29];
    ele[4][29] != ele[15][29];
    ele[4][29] != ele[16][29];
    ele[4][29] != ele[17][29];
    ele[4][29] != ele[18][29];
    ele[4][29] != ele[19][29];
    ele[4][29] != ele[20][29];
    ele[4][29] != ele[21][29];
    ele[4][29] != ele[22][29];
    ele[4][29] != ele[23][29];
    ele[4][29] != ele[24][29];
    ele[4][29] != ele[25][29];
    ele[4][29] != ele[26][29];
    ele[4][29] != ele[27][29];
    ele[4][29] != ele[28][29];
    ele[4][29] != ele[29][29];
    ele[4][29] != ele[30][29];
    ele[4][29] != ele[31][29];
    ele[4][29] != ele[32][29];
    ele[4][29] != ele[33][29];
    ele[4][29] != ele[34][29];
    ele[4][29] != ele[35][29];
    ele[4][29] != ele[4][30];
    ele[4][29] != ele[4][31];
    ele[4][29] != ele[4][32];
    ele[4][29] != ele[4][33];
    ele[4][29] != ele[4][34];
    ele[4][29] != ele[4][35];
    ele[4][29] != ele[5][24];
    ele[4][29] != ele[5][25];
    ele[4][29] != ele[5][26];
    ele[4][29] != ele[5][27];
    ele[4][29] != ele[5][28];
    ele[4][29] != ele[5][29];
    ele[4][29] != ele[6][29];
    ele[4][29] != ele[7][29];
    ele[4][29] != ele[8][29];
    ele[4][29] != ele[9][29];
    ele[4][3] != ele[10][3];
    ele[4][3] != ele[11][3];
    ele[4][3] != ele[12][3];
    ele[4][3] != ele[13][3];
    ele[4][3] != ele[14][3];
    ele[4][3] != ele[15][3];
    ele[4][3] != ele[16][3];
    ele[4][3] != ele[17][3];
    ele[4][3] != ele[18][3];
    ele[4][3] != ele[19][3];
    ele[4][3] != ele[20][3];
    ele[4][3] != ele[21][3];
    ele[4][3] != ele[22][3];
    ele[4][3] != ele[23][3];
    ele[4][3] != ele[24][3];
    ele[4][3] != ele[25][3];
    ele[4][3] != ele[26][3];
    ele[4][3] != ele[27][3];
    ele[4][3] != ele[28][3];
    ele[4][3] != ele[29][3];
    ele[4][3] != ele[30][3];
    ele[4][3] != ele[31][3];
    ele[4][3] != ele[32][3];
    ele[4][3] != ele[33][3];
    ele[4][3] != ele[34][3];
    ele[4][3] != ele[35][3];
    ele[4][3] != ele[4][10];
    ele[4][3] != ele[4][11];
    ele[4][3] != ele[4][12];
    ele[4][3] != ele[4][13];
    ele[4][3] != ele[4][14];
    ele[4][3] != ele[4][15];
    ele[4][3] != ele[4][16];
    ele[4][3] != ele[4][17];
    ele[4][3] != ele[4][18];
    ele[4][3] != ele[4][19];
    ele[4][3] != ele[4][20];
    ele[4][3] != ele[4][21];
    ele[4][3] != ele[4][22];
    ele[4][3] != ele[4][23];
    ele[4][3] != ele[4][24];
    ele[4][3] != ele[4][25];
    ele[4][3] != ele[4][26];
    ele[4][3] != ele[4][27];
    ele[4][3] != ele[4][28];
    ele[4][3] != ele[4][29];
    ele[4][3] != ele[4][30];
    ele[4][3] != ele[4][31];
    ele[4][3] != ele[4][32];
    ele[4][3] != ele[4][33];
    ele[4][3] != ele[4][34];
    ele[4][3] != ele[4][35];
    ele[4][3] != ele[4][4];
    ele[4][3] != ele[4][5];
    ele[4][3] != ele[4][6];
    ele[4][3] != ele[4][7];
    ele[4][3] != ele[4][8];
    ele[4][3] != ele[4][9];
    ele[4][3] != ele[5][0];
    ele[4][3] != ele[5][1];
    ele[4][3] != ele[5][2];
    ele[4][3] != ele[5][3];
    ele[4][3] != ele[5][4];
    ele[4][3] != ele[5][5];
    ele[4][3] != ele[6][3];
    ele[4][3] != ele[7][3];
    ele[4][3] != ele[8][3];
    ele[4][3] != ele[9][3];
    ele[4][30] != ele[10][30];
    ele[4][30] != ele[11][30];
    ele[4][30] != ele[12][30];
    ele[4][30] != ele[13][30];
    ele[4][30] != ele[14][30];
    ele[4][30] != ele[15][30];
    ele[4][30] != ele[16][30];
    ele[4][30] != ele[17][30];
    ele[4][30] != ele[18][30];
    ele[4][30] != ele[19][30];
    ele[4][30] != ele[20][30];
    ele[4][30] != ele[21][30];
    ele[4][30] != ele[22][30];
    ele[4][30] != ele[23][30];
    ele[4][30] != ele[24][30];
    ele[4][30] != ele[25][30];
    ele[4][30] != ele[26][30];
    ele[4][30] != ele[27][30];
    ele[4][30] != ele[28][30];
    ele[4][30] != ele[29][30];
    ele[4][30] != ele[30][30];
    ele[4][30] != ele[31][30];
    ele[4][30] != ele[32][30];
    ele[4][30] != ele[33][30];
    ele[4][30] != ele[34][30];
    ele[4][30] != ele[35][30];
    ele[4][30] != ele[4][31];
    ele[4][30] != ele[4][32];
    ele[4][30] != ele[4][33];
    ele[4][30] != ele[4][34];
    ele[4][30] != ele[4][35];
    ele[4][30] != ele[5][30];
    ele[4][30] != ele[5][31];
    ele[4][30] != ele[5][32];
    ele[4][30] != ele[5][33];
    ele[4][30] != ele[5][34];
    ele[4][30] != ele[5][35];
    ele[4][30] != ele[6][30];
    ele[4][30] != ele[7][30];
    ele[4][30] != ele[8][30];
    ele[4][30] != ele[9][30];
    ele[4][31] != ele[10][31];
    ele[4][31] != ele[11][31];
    ele[4][31] != ele[12][31];
    ele[4][31] != ele[13][31];
    ele[4][31] != ele[14][31];
    ele[4][31] != ele[15][31];
    ele[4][31] != ele[16][31];
    ele[4][31] != ele[17][31];
    ele[4][31] != ele[18][31];
    ele[4][31] != ele[19][31];
    ele[4][31] != ele[20][31];
    ele[4][31] != ele[21][31];
    ele[4][31] != ele[22][31];
    ele[4][31] != ele[23][31];
    ele[4][31] != ele[24][31];
    ele[4][31] != ele[25][31];
    ele[4][31] != ele[26][31];
    ele[4][31] != ele[27][31];
    ele[4][31] != ele[28][31];
    ele[4][31] != ele[29][31];
    ele[4][31] != ele[30][31];
    ele[4][31] != ele[31][31];
    ele[4][31] != ele[32][31];
    ele[4][31] != ele[33][31];
    ele[4][31] != ele[34][31];
    ele[4][31] != ele[35][31];
    ele[4][31] != ele[4][32];
    ele[4][31] != ele[4][33];
    ele[4][31] != ele[4][34];
    ele[4][31] != ele[4][35];
    ele[4][31] != ele[5][30];
    ele[4][31] != ele[5][31];
    ele[4][31] != ele[5][32];
    ele[4][31] != ele[5][33];
    ele[4][31] != ele[5][34];
    ele[4][31] != ele[5][35];
    ele[4][31] != ele[6][31];
    ele[4][31] != ele[7][31];
    ele[4][31] != ele[8][31];
    ele[4][31] != ele[9][31];
    ele[4][32] != ele[10][32];
    ele[4][32] != ele[11][32];
    ele[4][32] != ele[12][32];
    ele[4][32] != ele[13][32];
    ele[4][32] != ele[14][32];
    ele[4][32] != ele[15][32];
    ele[4][32] != ele[16][32];
    ele[4][32] != ele[17][32];
    ele[4][32] != ele[18][32];
    ele[4][32] != ele[19][32];
    ele[4][32] != ele[20][32];
    ele[4][32] != ele[21][32];
    ele[4][32] != ele[22][32];
    ele[4][32] != ele[23][32];
    ele[4][32] != ele[24][32];
    ele[4][32] != ele[25][32];
    ele[4][32] != ele[26][32];
    ele[4][32] != ele[27][32];
    ele[4][32] != ele[28][32];
    ele[4][32] != ele[29][32];
    ele[4][32] != ele[30][32];
    ele[4][32] != ele[31][32];
    ele[4][32] != ele[32][32];
    ele[4][32] != ele[33][32];
    ele[4][32] != ele[34][32];
    ele[4][32] != ele[35][32];
    ele[4][32] != ele[4][33];
    ele[4][32] != ele[4][34];
    ele[4][32] != ele[4][35];
    ele[4][32] != ele[5][30];
    ele[4][32] != ele[5][31];
    ele[4][32] != ele[5][32];
    ele[4][32] != ele[5][33];
    ele[4][32] != ele[5][34];
    ele[4][32] != ele[5][35];
    ele[4][32] != ele[6][32];
    ele[4][32] != ele[7][32];
    ele[4][32] != ele[8][32];
    ele[4][32] != ele[9][32];
    ele[4][33] != ele[10][33];
    ele[4][33] != ele[11][33];
    ele[4][33] != ele[12][33];
    ele[4][33] != ele[13][33];
    ele[4][33] != ele[14][33];
    ele[4][33] != ele[15][33];
    ele[4][33] != ele[16][33];
    ele[4][33] != ele[17][33];
    ele[4][33] != ele[18][33];
    ele[4][33] != ele[19][33];
    ele[4][33] != ele[20][33];
    ele[4][33] != ele[21][33];
    ele[4][33] != ele[22][33];
    ele[4][33] != ele[23][33];
    ele[4][33] != ele[24][33];
    ele[4][33] != ele[25][33];
    ele[4][33] != ele[26][33];
    ele[4][33] != ele[27][33];
    ele[4][33] != ele[28][33];
    ele[4][33] != ele[29][33];
    ele[4][33] != ele[30][33];
    ele[4][33] != ele[31][33];
    ele[4][33] != ele[32][33];
    ele[4][33] != ele[33][33];
    ele[4][33] != ele[34][33];
    ele[4][33] != ele[35][33];
    ele[4][33] != ele[4][34];
    ele[4][33] != ele[4][35];
    ele[4][33] != ele[5][30];
    ele[4][33] != ele[5][31];
    ele[4][33] != ele[5][32];
    ele[4][33] != ele[5][33];
    ele[4][33] != ele[5][34];
    ele[4][33] != ele[5][35];
    ele[4][33] != ele[6][33];
    ele[4][33] != ele[7][33];
    ele[4][33] != ele[8][33];
    ele[4][33] != ele[9][33];
    ele[4][34] != ele[10][34];
    ele[4][34] != ele[11][34];
    ele[4][34] != ele[12][34];
    ele[4][34] != ele[13][34];
    ele[4][34] != ele[14][34];
    ele[4][34] != ele[15][34];
    ele[4][34] != ele[16][34];
    ele[4][34] != ele[17][34];
    ele[4][34] != ele[18][34];
    ele[4][34] != ele[19][34];
    ele[4][34] != ele[20][34];
    ele[4][34] != ele[21][34];
    ele[4][34] != ele[22][34];
    ele[4][34] != ele[23][34];
    ele[4][34] != ele[24][34];
    ele[4][34] != ele[25][34];
    ele[4][34] != ele[26][34];
    ele[4][34] != ele[27][34];
    ele[4][34] != ele[28][34];
    ele[4][34] != ele[29][34];
    ele[4][34] != ele[30][34];
    ele[4][34] != ele[31][34];
    ele[4][34] != ele[32][34];
    ele[4][34] != ele[33][34];
    ele[4][34] != ele[34][34];
    ele[4][34] != ele[35][34];
    ele[4][34] != ele[4][35];
    ele[4][34] != ele[5][30];
    ele[4][34] != ele[5][31];
    ele[4][34] != ele[5][32];
    ele[4][34] != ele[5][33];
    ele[4][34] != ele[5][34];
    ele[4][34] != ele[5][35];
    ele[4][34] != ele[6][34];
    ele[4][34] != ele[7][34];
    ele[4][34] != ele[8][34];
    ele[4][34] != ele[9][34];
    ele[4][35] != ele[10][35];
    ele[4][35] != ele[11][35];
    ele[4][35] != ele[12][35];
    ele[4][35] != ele[13][35];
    ele[4][35] != ele[14][35];
    ele[4][35] != ele[15][35];
    ele[4][35] != ele[16][35];
    ele[4][35] != ele[17][35];
    ele[4][35] != ele[18][35];
    ele[4][35] != ele[19][35];
    ele[4][35] != ele[20][35];
    ele[4][35] != ele[21][35];
    ele[4][35] != ele[22][35];
    ele[4][35] != ele[23][35];
    ele[4][35] != ele[24][35];
    ele[4][35] != ele[25][35];
    ele[4][35] != ele[26][35];
    ele[4][35] != ele[27][35];
    ele[4][35] != ele[28][35];
    ele[4][35] != ele[29][35];
    ele[4][35] != ele[30][35];
    ele[4][35] != ele[31][35];
    ele[4][35] != ele[32][35];
    ele[4][35] != ele[33][35];
    ele[4][35] != ele[34][35];
    ele[4][35] != ele[35][35];
    ele[4][35] != ele[5][30];
    ele[4][35] != ele[5][31];
    ele[4][35] != ele[5][32];
    ele[4][35] != ele[5][33];
    ele[4][35] != ele[5][34];
    ele[4][35] != ele[5][35];
    ele[4][35] != ele[6][35];
    ele[4][35] != ele[7][35];
    ele[4][35] != ele[8][35];
    ele[4][35] != ele[9][35];
    ele[4][4] != ele[10][4];
    ele[4][4] != ele[11][4];
    ele[4][4] != ele[12][4];
    ele[4][4] != ele[13][4];
    ele[4][4] != ele[14][4];
    ele[4][4] != ele[15][4];
    ele[4][4] != ele[16][4];
    ele[4][4] != ele[17][4];
    ele[4][4] != ele[18][4];
    ele[4][4] != ele[19][4];
    ele[4][4] != ele[20][4];
    ele[4][4] != ele[21][4];
    ele[4][4] != ele[22][4];
    ele[4][4] != ele[23][4];
    ele[4][4] != ele[24][4];
    ele[4][4] != ele[25][4];
    ele[4][4] != ele[26][4];
    ele[4][4] != ele[27][4];
    ele[4][4] != ele[28][4];
    ele[4][4] != ele[29][4];
    ele[4][4] != ele[30][4];
    ele[4][4] != ele[31][4];
    ele[4][4] != ele[32][4];
    ele[4][4] != ele[33][4];
    ele[4][4] != ele[34][4];
    ele[4][4] != ele[35][4];
    ele[4][4] != ele[4][10];
    ele[4][4] != ele[4][11];
    ele[4][4] != ele[4][12];
    ele[4][4] != ele[4][13];
    ele[4][4] != ele[4][14];
    ele[4][4] != ele[4][15];
    ele[4][4] != ele[4][16];
    ele[4][4] != ele[4][17];
    ele[4][4] != ele[4][18];
    ele[4][4] != ele[4][19];
    ele[4][4] != ele[4][20];
    ele[4][4] != ele[4][21];
    ele[4][4] != ele[4][22];
    ele[4][4] != ele[4][23];
    ele[4][4] != ele[4][24];
    ele[4][4] != ele[4][25];
    ele[4][4] != ele[4][26];
    ele[4][4] != ele[4][27];
    ele[4][4] != ele[4][28];
    ele[4][4] != ele[4][29];
    ele[4][4] != ele[4][30];
    ele[4][4] != ele[4][31];
    ele[4][4] != ele[4][32];
    ele[4][4] != ele[4][33];
    ele[4][4] != ele[4][34];
    ele[4][4] != ele[4][35];
    ele[4][4] != ele[4][5];
    ele[4][4] != ele[4][6];
    ele[4][4] != ele[4][7];
    ele[4][4] != ele[4][8];
    ele[4][4] != ele[4][9];
    ele[4][4] != ele[5][0];
    ele[4][4] != ele[5][1];
    ele[4][4] != ele[5][2];
    ele[4][4] != ele[5][3];
    ele[4][4] != ele[5][4];
    ele[4][4] != ele[5][5];
    ele[4][4] != ele[6][4];
    ele[4][4] != ele[7][4];
    ele[4][4] != ele[8][4];
    ele[4][4] != ele[9][4];
    ele[4][5] != ele[10][5];
    ele[4][5] != ele[11][5];
    ele[4][5] != ele[12][5];
    ele[4][5] != ele[13][5];
    ele[4][5] != ele[14][5];
    ele[4][5] != ele[15][5];
    ele[4][5] != ele[16][5];
    ele[4][5] != ele[17][5];
    ele[4][5] != ele[18][5];
    ele[4][5] != ele[19][5];
    ele[4][5] != ele[20][5];
    ele[4][5] != ele[21][5];
    ele[4][5] != ele[22][5];
    ele[4][5] != ele[23][5];
    ele[4][5] != ele[24][5];
    ele[4][5] != ele[25][5];
    ele[4][5] != ele[26][5];
    ele[4][5] != ele[27][5];
    ele[4][5] != ele[28][5];
    ele[4][5] != ele[29][5];
    ele[4][5] != ele[30][5];
    ele[4][5] != ele[31][5];
    ele[4][5] != ele[32][5];
    ele[4][5] != ele[33][5];
    ele[4][5] != ele[34][5];
    ele[4][5] != ele[35][5];
    ele[4][5] != ele[4][10];
    ele[4][5] != ele[4][11];
    ele[4][5] != ele[4][12];
    ele[4][5] != ele[4][13];
    ele[4][5] != ele[4][14];
    ele[4][5] != ele[4][15];
    ele[4][5] != ele[4][16];
    ele[4][5] != ele[4][17];
    ele[4][5] != ele[4][18];
    ele[4][5] != ele[4][19];
    ele[4][5] != ele[4][20];
    ele[4][5] != ele[4][21];
    ele[4][5] != ele[4][22];
    ele[4][5] != ele[4][23];
    ele[4][5] != ele[4][24];
    ele[4][5] != ele[4][25];
    ele[4][5] != ele[4][26];
    ele[4][5] != ele[4][27];
    ele[4][5] != ele[4][28];
    ele[4][5] != ele[4][29];
    ele[4][5] != ele[4][30];
    ele[4][5] != ele[4][31];
    ele[4][5] != ele[4][32];
    ele[4][5] != ele[4][33];
    ele[4][5] != ele[4][34];
    ele[4][5] != ele[4][35];
    ele[4][5] != ele[4][6];
    ele[4][5] != ele[4][7];
    ele[4][5] != ele[4][8];
    ele[4][5] != ele[4][9];
    ele[4][5] != ele[5][0];
    ele[4][5] != ele[5][1];
    ele[4][5] != ele[5][2];
    ele[4][5] != ele[5][3];
    ele[4][5] != ele[5][4];
    ele[4][5] != ele[5][5];
    ele[4][5] != ele[6][5];
    ele[4][5] != ele[7][5];
    ele[4][5] != ele[8][5];
    ele[4][5] != ele[9][5];
    ele[4][6] != ele[10][6];
    ele[4][6] != ele[11][6];
    ele[4][6] != ele[12][6];
    ele[4][6] != ele[13][6];
    ele[4][6] != ele[14][6];
    ele[4][6] != ele[15][6];
    ele[4][6] != ele[16][6];
    ele[4][6] != ele[17][6];
    ele[4][6] != ele[18][6];
    ele[4][6] != ele[19][6];
    ele[4][6] != ele[20][6];
    ele[4][6] != ele[21][6];
    ele[4][6] != ele[22][6];
    ele[4][6] != ele[23][6];
    ele[4][6] != ele[24][6];
    ele[4][6] != ele[25][6];
    ele[4][6] != ele[26][6];
    ele[4][6] != ele[27][6];
    ele[4][6] != ele[28][6];
    ele[4][6] != ele[29][6];
    ele[4][6] != ele[30][6];
    ele[4][6] != ele[31][6];
    ele[4][6] != ele[32][6];
    ele[4][6] != ele[33][6];
    ele[4][6] != ele[34][6];
    ele[4][6] != ele[35][6];
    ele[4][6] != ele[4][10];
    ele[4][6] != ele[4][11];
    ele[4][6] != ele[4][12];
    ele[4][6] != ele[4][13];
    ele[4][6] != ele[4][14];
    ele[4][6] != ele[4][15];
    ele[4][6] != ele[4][16];
    ele[4][6] != ele[4][17];
    ele[4][6] != ele[4][18];
    ele[4][6] != ele[4][19];
    ele[4][6] != ele[4][20];
    ele[4][6] != ele[4][21];
    ele[4][6] != ele[4][22];
    ele[4][6] != ele[4][23];
    ele[4][6] != ele[4][24];
    ele[4][6] != ele[4][25];
    ele[4][6] != ele[4][26];
    ele[4][6] != ele[4][27];
    ele[4][6] != ele[4][28];
    ele[4][6] != ele[4][29];
    ele[4][6] != ele[4][30];
    ele[4][6] != ele[4][31];
    ele[4][6] != ele[4][32];
    ele[4][6] != ele[4][33];
    ele[4][6] != ele[4][34];
    ele[4][6] != ele[4][35];
    ele[4][6] != ele[4][7];
    ele[4][6] != ele[4][8];
    ele[4][6] != ele[4][9];
    ele[4][6] != ele[5][10];
    ele[4][6] != ele[5][11];
    ele[4][6] != ele[5][6];
    ele[4][6] != ele[5][7];
    ele[4][6] != ele[5][8];
    ele[4][6] != ele[5][9];
    ele[4][6] != ele[6][6];
    ele[4][6] != ele[7][6];
    ele[4][6] != ele[8][6];
    ele[4][6] != ele[9][6];
    ele[4][7] != ele[10][7];
    ele[4][7] != ele[11][7];
    ele[4][7] != ele[12][7];
    ele[4][7] != ele[13][7];
    ele[4][7] != ele[14][7];
    ele[4][7] != ele[15][7];
    ele[4][7] != ele[16][7];
    ele[4][7] != ele[17][7];
    ele[4][7] != ele[18][7];
    ele[4][7] != ele[19][7];
    ele[4][7] != ele[20][7];
    ele[4][7] != ele[21][7];
    ele[4][7] != ele[22][7];
    ele[4][7] != ele[23][7];
    ele[4][7] != ele[24][7];
    ele[4][7] != ele[25][7];
    ele[4][7] != ele[26][7];
    ele[4][7] != ele[27][7];
    ele[4][7] != ele[28][7];
    ele[4][7] != ele[29][7];
    ele[4][7] != ele[30][7];
    ele[4][7] != ele[31][7];
    ele[4][7] != ele[32][7];
    ele[4][7] != ele[33][7];
    ele[4][7] != ele[34][7];
    ele[4][7] != ele[35][7];
    ele[4][7] != ele[4][10];
    ele[4][7] != ele[4][11];
    ele[4][7] != ele[4][12];
    ele[4][7] != ele[4][13];
    ele[4][7] != ele[4][14];
    ele[4][7] != ele[4][15];
    ele[4][7] != ele[4][16];
    ele[4][7] != ele[4][17];
    ele[4][7] != ele[4][18];
    ele[4][7] != ele[4][19];
    ele[4][7] != ele[4][20];
    ele[4][7] != ele[4][21];
    ele[4][7] != ele[4][22];
    ele[4][7] != ele[4][23];
    ele[4][7] != ele[4][24];
    ele[4][7] != ele[4][25];
    ele[4][7] != ele[4][26];
    ele[4][7] != ele[4][27];
    ele[4][7] != ele[4][28];
    ele[4][7] != ele[4][29];
    ele[4][7] != ele[4][30];
    ele[4][7] != ele[4][31];
    ele[4][7] != ele[4][32];
    ele[4][7] != ele[4][33];
    ele[4][7] != ele[4][34];
    ele[4][7] != ele[4][35];
    ele[4][7] != ele[4][8];
    ele[4][7] != ele[4][9];
    ele[4][7] != ele[5][10];
    ele[4][7] != ele[5][11];
    ele[4][7] != ele[5][6];
    ele[4][7] != ele[5][7];
    ele[4][7] != ele[5][8];
    ele[4][7] != ele[5][9];
    ele[4][7] != ele[6][7];
    ele[4][7] != ele[7][7];
    ele[4][7] != ele[8][7];
    ele[4][7] != ele[9][7];
    ele[4][8] != ele[10][8];
    ele[4][8] != ele[11][8];
    ele[4][8] != ele[12][8];
    ele[4][8] != ele[13][8];
    ele[4][8] != ele[14][8];
    ele[4][8] != ele[15][8];
    ele[4][8] != ele[16][8];
    ele[4][8] != ele[17][8];
    ele[4][8] != ele[18][8];
    ele[4][8] != ele[19][8];
    ele[4][8] != ele[20][8];
    ele[4][8] != ele[21][8];
    ele[4][8] != ele[22][8];
    ele[4][8] != ele[23][8];
    ele[4][8] != ele[24][8];
    ele[4][8] != ele[25][8];
    ele[4][8] != ele[26][8];
    ele[4][8] != ele[27][8];
    ele[4][8] != ele[28][8];
    ele[4][8] != ele[29][8];
    ele[4][8] != ele[30][8];
    ele[4][8] != ele[31][8];
    ele[4][8] != ele[32][8];
    ele[4][8] != ele[33][8];
    ele[4][8] != ele[34][8];
    ele[4][8] != ele[35][8];
    ele[4][8] != ele[4][10];
    ele[4][8] != ele[4][11];
    ele[4][8] != ele[4][12];
    ele[4][8] != ele[4][13];
    ele[4][8] != ele[4][14];
    ele[4][8] != ele[4][15];
    ele[4][8] != ele[4][16];
    ele[4][8] != ele[4][17];
    ele[4][8] != ele[4][18];
    ele[4][8] != ele[4][19];
    ele[4][8] != ele[4][20];
    ele[4][8] != ele[4][21];
    ele[4][8] != ele[4][22];
    ele[4][8] != ele[4][23];
    ele[4][8] != ele[4][24];
    ele[4][8] != ele[4][25];
    ele[4][8] != ele[4][26];
    ele[4][8] != ele[4][27];
    ele[4][8] != ele[4][28];
    ele[4][8] != ele[4][29];
    ele[4][8] != ele[4][30];
    ele[4][8] != ele[4][31];
    ele[4][8] != ele[4][32];
    ele[4][8] != ele[4][33];
    ele[4][8] != ele[4][34];
    ele[4][8] != ele[4][35];
    ele[4][8] != ele[4][9];
    ele[4][8] != ele[5][10];
    ele[4][8] != ele[5][11];
    ele[4][8] != ele[5][6];
    ele[4][8] != ele[5][7];
    ele[4][8] != ele[5][8];
    ele[4][8] != ele[5][9];
    ele[4][8] != ele[6][8];
    ele[4][8] != ele[7][8];
    ele[4][8] != ele[8][8];
    ele[4][8] != ele[9][8];
    ele[4][9] != ele[10][9];
    ele[4][9] != ele[11][9];
    ele[4][9] != ele[12][9];
    ele[4][9] != ele[13][9];
    ele[4][9] != ele[14][9];
    ele[4][9] != ele[15][9];
    ele[4][9] != ele[16][9];
    ele[4][9] != ele[17][9];
    ele[4][9] != ele[18][9];
    ele[4][9] != ele[19][9];
    ele[4][9] != ele[20][9];
    ele[4][9] != ele[21][9];
    ele[4][9] != ele[22][9];
    ele[4][9] != ele[23][9];
    ele[4][9] != ele[24][9];
    ele[4][9] != ele[25][9];
    ele[4][9] != ele[26][9];
    ele[4][9] != ele[27][9];
    ele[4][9] != ele[28][9];
    ele[4][9] != ele[29][9];
    ele[4][9] != ele[30][9];
    ele[4][9] != ele[31][9];
    ele[4][9] != ele[32][9];
    ele[4][9] != ele[33][9];
    ele[4][9] != ele[34][9];
    ele[4][9] != ele[35][9];
    ele[4][9] != ele[4][10];
    ele[4][9] != ele[4][11];
    ele[4][9] != ele[4][12];
    ele[4][9] != ele[4][13];
    ele[4][9] != ele[4][14];
    ele[4][9] != ele[4][15];
    ele[4][9] != ele[4][16];
    ele[4][9] != ele[4][17];
    ele[4][9] != ele[4][18];
    ele[4][9] != ele[4][19];
    ele[4][9] != ele[4][20];
    ele[4][9] != ele[4][21];
    ele[4][9] != ele[4][22];
    ele[4][9] != ele[4][23];
    ele[4][9] != ele[4][24];
    ele[4][9] != ele[4][25];
    ele[4][9] != ele[4][26];
    ele[4][9] != ele[4][27];
    ele[4][9] != ele[4][28];
    ele[4][9] != ele[4][29];
    ele[4][9] != ele[4][30];
    ele[4][9] != ele[4][31];
    ele[4][9] != ele[4][32];
    ele[4][9] != ele[4][33];
    ele[4][9] != ele[4][34];
    ele[4][9] != ele[4][35];
    ele[4][9] != ele[5][10];
    ele[4][9] != ele[5][11];
    ele[4][9] != ele[5][6];
    ele[4][9] != ele[5][7];
    ele[4][9] != ele[5][8];
    ele[4][9] != ele[5][9];
    ele[4][9] != ele[6][9];
    ele[4][9] != ele[7][9];
    ele[4][9] != ele[8][9];
    ele[4][9] != ele[9][9];
    ele[5][0] != ele[10][0];
    ele[5][0] != ele[11][0];
    ele[5][0] != ele[12][0];
    ele[5][0] != ele[13][0];
    ele[5][0] != ele[14][0];
    ele[5][0] != ele[15][0];
    ele[5][0] != ele[16][0];
    ele[5][0] != ele[17][0];
    ele[5][0] != ele[18][0];
    ele[5][0] != ele[19][0];
    ele[5][0] != ele[20][0];
    ele[5][0] != ele[21][0];
    ele[5][0] != ele[22][0];
    ele[5][0] != ele[23][0];
    ele[5][0] != ele[24][0];
    ele[5][0] != ele[25][0];
    ele[5][0] != ele[26][0];
    ele[5][0] != ele[27][0];
    ele[5][0] != ele[28][0];
    ele[5][0] != ele[29][0];
    ele[5][0] != ele[30][0];
    ele[5][0] != ele[31][0];
    ele[5][0] != ele[32][0];
    ele[5][0] != ele[33][0];
    ele[5][0] != ele[34][0];
    ele[5][0] != ele[35][0];
    ele[5][0] != ele[5][1];
    ele[5][0] != ele[5][10];
    ele[5][0] != ele[5][11];
    ele[5][0] != ele[5][12];
    ele[5][0] != ele[5][13];
    ele[5][0] != ele[5][14];
    ele[5][0] != ele[5][15];
    ele[5][0] != ele[5][16];
    ele[5][0] != ele[5][17];
    ele[5][0] != ele[5][18];
    ele[5][0] != ele[5][19];
    ele[5][0] != ele[5][2];
    ele[5][0] != ele[5][20];
    ele[5][0] != ele[5][21];
    ele[5][0] != ele[5][22];
    ele[5][0] != ele[5][23];
    ele[5][0] != ele[5][24];
    ele[5][0] != ele[5][25];
    ele[5][0] != ele[5][26];
    ele[5][0] != ele[5][27];
    ele[5][0] != ele[5][28];
    ele[5][0] != ele[5][29];
    ele[5][0] != ele[5][3];
    ele[5][0] != ele[5][30];
    ele[5][0] != ele[5][31];
    ele[5][0] != ele[5][32];
    ele[5][0] != ele[5][33];
    ele[5][0] != ele[5][34];
    ele[5][0] != ele[5][35];
    ele[5][0] != ele[5][4];
    ele[5][0] != ele[5][5];
    ele[5][0] != ele[5][6];
    ele[5][0] != ele[5][7];
    ele[5][0] != ele[5][8];
    ele[5][0] != ele[5][9];
    ele[5][0] != ele[6][0];
    ele[5][0] != ele[7][0];
    ele[5][0] != ele[8][0];
    ele[5][0] != ele[9][0];
    ele[5][1] != ele[10][1];
    ele[5][1] != ele[11][1];
    ele[5][1] != ele[12][1];
    ele[5][1] != ele[13][1];
    ele[5][1] != ele[14][1];
    ele[5][1] != ele[15][1];
    ele[5][1] != ele[16][1];
    ele[5][1] != ele[17][1];
    ele[5][1] != ele[18][1];
    ele[5][1] != ele[19][1];
    ele[5][1] != ele[20][1];
    ele[5][1] != ele[21][1];
    ele[5][1] != ele[22][1];
    ele[5][1] != ele[23][1];
    ele[5][1] != ele[24][1];
    ele[5][1] != ele[25][1];
    ele[5][1] != ele[26][1];
    ele[5][1] != ele[27][1];
    ele[5][1] != ele[28][1];
    ele[5][1] != ele[29][1];
    ele[5][1] != ele[30][1];
    ele[5][1] != ele[31][1];
    ele[5][1] != ele[32][1];
    ele[5][1] != ele[33][1];
    ele[5][1] != ele[34][1];
    ele[5][1] != ele[35][1];
    ele[5][1] != ele[5][10];
    ele[5][1] != ele[5][11];
    ele[5][1] != ele[5][12];
    ele[5][1] != ele[5][13];
    ele[5][1] != ele[5][14];
    ele[5][1] != ele[5][15];
    ele[5][1] != ele[5][16];
    ele[5][1] != ele[5][17];
    ele[5][1] != ele[5][18];
    ele[5][1] != ele[5][19];
    ele[5][1] != ele[5][2];
    ele[5][1] != ele[5][20];
    ele[5][1] != ele[5][21];
    ele[5][1] != ele[5][22];
    ele[5][1] != ele[5][23];
    ele[5][1] != ele[5][24];
    ele[5][1] != ele[5][25];
    ele[5][1] != ele[5][26];
    ele[5][1] != ele[5][27];
    ele[5][1] != ele[5][28];
    ele[5][1] != ele[5][29];
    ele[5][1] != ele[5][3];
    ele[5][1] != ele[5][30];
    ele[5][1] != ele[5][31];
    ele[5][1] != ele[5][32];
    ele[5][1] != ele[5][33];
    ele[5][1] != ele[5][34];
    ele[5][1] != ele[5][35];
    ele[5][1] != ele[5][4];
    ele[5][1] != ele[5][5];
    ele[5][1] != ele[5][6];
    ele[5][1] != ele[5][7];
    ele[5][1] != ele[5][8];
    ele[5][1] != ele[5][9];
    ele[5][1] != ele[6][1];
    ele[5][1] != ele[7][1];
    ele[5][1] != ele[8][1];
    ele[5][1] != ele[9][1];
    ele[5][10] != ele[10][10];
    ele[5][10] != ele[11][10];
    ele[5][10] != ele[12][10];
    ele[5][10] != ele[13][10];
    ele[5][10] != ele[14][10];
    ele[5][10] != ele[15][10];
    ele[5][10] != ele[16][10];
    ele[5][10] != ele[17][10];
    ele[5][10] != ele[18][10];
    ele[5][10] != ele[19][10];
    ele[5][10] != ele[20][10];
    ele[5][10] != ele[21][10];
    ele[5][10] != ele[22][10];
    ele[5][10] != ele[23][10];
    ele[5][10] != ele[24][10];
    ele[5][10] != ele[25][10];
    ele[5][10] != ele[26][10];
    ele[5][10] != ele[27][10];
    ele[5][10] != ele[28][10];
    ele[5][10] != ele[29][10];
    ele[5][10] != ele[30][10];
    ele[5][10] != ele[31][10];
    ele[5][10] != ele[32][10];
    ele[5][10] != ele[33][10];
    ele[5][10] != ele[34][10];
    ele[5][10] != ele[35][10];
    ele[5][10] != ele[5][11];
    ele[5][10] != ele[5][12];
    ele[5][10] != ele[5][13];
    ele[5][10] != ele[5][14];
    ele[5][10] != ele[5][15];
    ele[5][10] != ele[5][16];
    ele[5][10] != ele[5][17];
    ele[5][10] != ele[5][18];
    ele[5][10] != ele[5][19];
    ele[5][10] != ele[5][20];
    ele[5][10] != ele[5][21];
    ele[5][10] != ele[5][22];
    ele[5][10] != ele[5][23];
    ele[5][10] != ele[5][24];
    ele[5][10] != ele[5][25];
    ele[5][10] != ele[5][26];
    ele[5][10] != ele[5][27];
    ele[5][10] != ele[5][28];
    ele[5][10] != ele[5][29];
    ele[5][10] != ele[5][30];
    ele[5][10] != ele[5][31];
    ele[5][10] != ele[5][32];
    ele[5][10] != ele[5][33];
    ele[5][10] != ele[5][34];
    ele[5][10] != ele[5][35];
    ele[5][10] != ele[6][10];
    ele[5][10] != ele[7][10];
    ele[5][10] != ele[8][10];
    ele[5][10] != ele[9][10];
    ele[5][11] != ele[10][11];
    ele[5][11] != ele[11][11];
    ele[5][11] != ele[12][11];
    ele[5][11] != ele[13][11];
    ele[5][11] != ele[14][11];
    ele[5][11] != ele[15][11];
    ele[5][11] != ele[16][11];
    ele[5][11] != ele[17][11];
    ele[5][11] != ele[18][11];
    ele[5][11] != ele[19][11];
    ele[5][11] != ele[20][11];
    ele[5][11] != ele[21][11];
    ele[5][11] != ele[22][11];
    ele[5][11] != ele[23][11];
    ele[5][11] != ele[24][11];
    ele[5][11] != ele[25][11];
    ele[5][11] != ele[26][11];
    ele[5][11] != ele[27][11];
    ele[5][11] != ele[28][11];
    ele[5][11] != ele[29][11];
    ele[5][11] != ele[30][11];
    ele[5][11] != ele[31][11];
    ele[5][11] != ele[32][11];
    ele[5][11] != ele[33][11];
    ele[5][11] != ele[34][11];
    ele[5][11] != ele[35][11];
    ele[5][11] != ele[5][12];
    ele[5][11] != ele[5][13];
    ele[5][11] != ele[5][14];
    ele[5][11] != ele[5][15];
    ele[5][11] != ele[5][16];
    ele[5][11] != ele[5][17];
    ele[5][11] != ele[5][18];
    ele[5][11] != ele[5][19];
    ele[5][11] != ele[5][20];
    ele[5][11] != ele[5][21];
    ele[5][11] != ele[5][22];
    ele[5][11] != ele[5][23];
    ele[5][11] != ele[5][24];
    ele[5][11] != ele[5][25];
    ele[5][11] != ele[5][26];
    ele[5][11] != ele[5][27];
    ele[5][11] != ele[5][28];
    ele[5][11] != ele[5][29];
    ele[5][11] != ele[5][30];
    ele[5][11] != ele[5][31];
    ele[5][11] != ele[5][32];
    ele[5][11] != ele[5][33];
    ele[5][11] != ele[5][34];
    ele[5][11] != ele[5][35];
    ele[5][11] != ele[6][11];
    ele[5][11] != ele[7][11];
    ele[5][11] != ele[8][11];
    ele[5][11] != ele[9][11];
    ele[5][12] != ele[10][12];
    ele[5][12] != ele[11][12];
    ele[5][12] != ele[12][12];
    ele[5][12] != ele[13][12];
    ele[5][12] != ele[14][12];
    ele[5][12] != ele[15][12];
    ele[5][12] != ele[16][12];
    ele[5][12] != ele[17][12];
    ele[5][12] != ele[18][12];
    ele[5][12] != ele[19][12];
    ele[5][12] != ele[20][12];
    ele[5][12] != ele[21][12];
    ele[5][12] != ele[22][12];
    ele[5][12] != ele[23][12];
    ele[5][12] != ele[24][12];
    ele[5][12] != ele[25][12];
    ele[5][12] != ele[26][12];
    ele[5][12] != ele[27][12];
    ele[5][12] != ele[28][12];
    ele[5][12] != ele[29][12];
    ele[5][12] != ele[30][12];
    ele[5][12] != ele[31][12];
    ele[5][12] != ele[32][12];
    ele[5][12] != ele[33][12];
    ele[5][12] != ele[34][12];
    ele[5][12] != ele[35][12];
    ele[5][12] != ele[5][13];
    ele[5][12] != ele[5][14];
    ele[5][12] != ele[5][15];
    ele[5][12] != ele[5][16];
    ele[5][12] != ele[5][17];
    ele[5][12] != ele[5][18];
    ele[5][12] != ele[5][19];
    ele[5][12] != ele[5][20];
    ele[5][12] != ele[5][21];
    ele[5][12] != ele[5][22];
    ele[5][12] != ele[5][23];
    ele[5][12] != ele[5][24];
    ele[5][12] != ele[5][25];
    ele[5][12] != ele[5][26];
    ele[5][12] != ele[5][27];
    ele[5][12] != ele[5][28];
    ele[5][12] != ele[5][29];
    ele[5][12] != ele[5][30];
    ele[5][12] != ele[5][31];
    ele[5][12] != ele[5][32];
    ele[5][12] != ele[5][33];
    ele[5][12] != ele[5][34];
    ele[5][12] != ele[5][35];
    ele[5][12] != ele[6][12];
    ele[5][12] != ele[7][12];
    ele[5][12] != ele[8][12];
    ele[5][12] != ele[9][12];
    ele[5][13] != ele[10][13];
    ele[5][13] != ele[11][13];
    ele[5][13] != ele[12][13];
    ele[5][13] != ele[13][13];
    ele[5][13] != ele[14][13];
    ele[5][13] != ele[15][13];
    ele[5][13] != ele[16][13];
    ele[5][13] != ele[17][13];
    ele[5][13] != ele[18][13];
    ele[5][13] != ele[19][13];
    ele[5][13] != ele[20][13];
    ele[5][13] != ele[21][13];
    ele[5][13] != ele[22][13];
    ele[5][13] != ele[23][13];
    ele[5][13] != ele[24][13];
    ele[5][13] != ele[25][13];
    ele[5][13] != ele[26][13];
    ele[5][13] != ele[27][13];
    ele[5][13] != ele[28][13];
    ele[5][13] != ele[29][13];
    ele[5][13] != ele[30][13];
    ele[5][13] != ele[31][13];
    ele[5][13] != ele[32][13];
    ele[5][13] != ele[33][13];
    ele[5][13] != ele[34][13];
    ele[5][13] != ele[35][13];
    ele[5][13] != ele[5][14];
    ele[5][13] != ele[5][15];
    ele[5][13] != ele[5][16];
    ele[5][13] != ele[5][17];
    ele[5][13] != ele[5][18];
    ele[5][13] != ele[5][19];
    ele[5][13] != ele[5][20];
    ele[5][13] != ele[5][21];
    ele[5][13] != ele[5][22];
    ele[5][13] != ele[5][23];
    ele[5][13] != ele[5][24];
    ele[5][13] != ele[5][25];
    ele[5][13] != ele[5][26];
    ele[5][13] != ele[5][27];
    ele[5][13] != ele[5][28];
    ele[5][13] != ele[5][29];
    ele[5][13] != ele[5][30];
    ele[5][13] != ele[5][31];
    ele[5][13] != ele[5][32];
    ele[5][13] != ele[5][33];
    ele[5][13] != ele[5][34];
    ele[5][13] != ele[5][35];
    ele[5][13] != ele[6][13];
    ele[5][13] != ele[7][13];
    ele[5][13] != ele[8][13];
    ele[5][13] != ele[9][13];
    ele[5][14] != ele[10][14];
    ele[5][14] != ele[11][14];
    ele[5][14] != ele[12][14];
    ele[5][14] != ele[13][14];
    ele[5][14] != ele[14][14];
    ele[5][14] != ele[15][14];
    ele[5][14] != ele[16][14];
    ele[5][14] != ele[17][14];
    ele[5][14] != ele[18][14];
    ele[5][14] != ele[19][14];
    ele[5][14] != ele[20][14];
    ele[5][14] != ele[21][14];
    ele[5][14] != ele[22][14];
    ele[5][14] != ele[23][14];
    ele[5][14] != ele[24][14];
    ele[5][14] != ele[25][14];
    ele[5][14] != ele[26][14];
    ele[5][14] != ele[27][14];
    ele[5][14] != ele[28][14];
    ele[5][14] != ele[29][14];
    ele[5][14] != ele[30][14];
    ele[5][14] != ele[31][14];
    ele[5][14] != ele[32][14];
    ele[5][14] != ele[33][14];
    ele[5][14] != ele[34][14];
    ele[5][14] != ele[35][14];
    ele[5][14] != ele[5][15];
    ele[5][14] != ele[5][16];
    ele[5][14] != ele[5][17];
    ele[5][14] != ele[5][18];
    ele[5][14] != ele[5][19];
    ele[5][14] != ele[5][20];
    ele[5][14] != ele[5][21];
    ele[5][14] != ele[5][22];
    ele[5][14] != ele[5][23];
    ele[5][14] != ele[5][24];
    ele[5][14] != ele[5][25];
    ele[5][14] != ele[5][26];
    ele[5][14] != ele[5][27];
    ele[5][14] != ele[5][28];
    ele[5][14] != ele[5][29];
    ele[5][14] != ele[5][30];
    ele[5][14] != ele[5][31];
    ele[5][14] != ele[5][32];
    ele[5][14] != ele[5][33];
    ele[5][14] != ele[5][34];
    ele[5][14] != ele[5][35];
    ele[5][14] != ele[6][14];
    ele[5][14] != ele[7][14];
    ele[5][14] != ele[8][14];
    ele[5][14] != ele[9][14];
    ele[5][15] != ele[10][15];
    ele[5][15] != ele[11][15];
    ele[5][15] != ele[12][15];
    ele[5][15] != ele[13][15];
    ele[5][15] != ele[14][15];
    ele[5][15] != ele[15][15];
    ele[5][15] != ele[16][15];
    ele[5][15] != ele[17][15];
    ele[5][15] != ele[18][15];
    ele[5][15] != ele[19][15];
    ele[5][15] != ele[20][15];
    ele[5][15] != ele[21][15];
    ele[5][15] != ele[22][15];
    ele[5][15] != ele[23][15];
    ele[5][15] != ele[24][15];
    ele[5][15] != ele[25][15];
    ele[5][15] != ele[26][15];
    ele[5][15] != ele[27][15];
    ele[5][15] != ele[28][15];
    ele[5][15] != ele[29][15];
    ele[5][15] != ele[30][15];
    ele[5][15] != ele[31][15];
    ele[5][15] != ele[32][15];
    ele[5][15] != ele[33][15];
    ele[5][15] != ele[34][15];
    ele[5][15] != ele[35][15];
    ele[5][15] != ele[5][16];
    ele[5][15] != ele[5][17];
    ele[5][15] != ele[5][18];
    ele[5][15] != ele[5][19];
    ele[5][15] != ele[5][20];
    ele[5][15] != ele[5][21];
    ele[5][15] != ele[5][22];
    ele[5][15] != ele[5][23];
    ele[5][15] != ele[5][24];
    ele[5][15] != ele[5][25];
    ele[5][15] != ele[5][26];
    ele[5][15] != ele[5][27];
    ele[5][15] != ele[5][28];
    ele[5][15] != ele[5][29];
    ele[5][15] != ele[5][30];
    ele[5][15] != ele[5][31];
    ele[5][15] != ele[5][32];
    ele[5][15] != ele[5][33];
    ele[5][15] != ele[5][34];
    ele[5][15] != ele[5][35];
    ele[5][15] != ele[6][15];
    ele[5][15] != ele[7][15];
    ele[5][15] != ele[8][15];
    ele[5][15] != ele[9][15];
    ele[5][16] != ele[10][16];
    ele[5][16] != ele[11][16];
    ele[5][16] != ele[12][16];
    ele[5][16] != ele[13][16];
    ele[5][16] != ele[14][16];
    ele[5][16] != ele[15][16];
    ele[5][16] != ele[16][16];
    ele[5][16] != ele[17][16];
    ele[5][16] != ele[18][16];
    ele[5][16] != ele[19][16];
    ele[5][16] != ele[20][16];
    ele[5][16] != ele[21][16];
    ele[5][16] != ele[22][16];
    ele[5][16] != ele[23][16];
    ele[5][16] != ele[24][16];
    ele[5][16] != ele[25][16];
    ele[5][16] != ele[26][16];
    ele[5][16] != ele[27][16];
    ele[5][16] != ele[28][16];
    ele[5][16] != ele[29][16];
    ele[5][16] != ele[30][16];
    ele[5][16] != ele[31][16];
    ele[5][16] != ele[32][16];
    ele[5][16] != ele[33][16];
    ele[5][16] != ele[34][16];
    ele[5][16] != ele[35][16];
    ele[5][16] != ele[5][17];
    ele[5][16] != ele[5][18];
    ele[5][16] != ele[5][19];
    ele[5][16] != ele[5][20];
    ele[5][16] != ele[5][21];
    ele[5][16] != ele[5][22];
    ele[5][16] != ele[5][23];
    ele[5][16] != ele[5][24];
    ele[5][16] != ele[5][25];
    ele[5][16] != ele[5][26];
    ele[5][16] != ele[5][27];
    ele[5][16] != ele[5][28];
    ele[5][16] != ele[5][29];
    ele[5][16] != ele[5][30];
    ele[5][16] != ele[5][31];
    ele[5][16] != ele[5][32];
    ele[5][16] != ele[5][33];
    ele[5][16] != ele[5][34];
    ele[5][16] != ele[5][35];
    ele[5][16] != ele[6][16];
    ele[5][16] != ele[7][16];
    ele[5][16] != ele[8][16];
    ele[5][16] != ele[9][16];
    ele[5][17] != ele[10][17];
    ele[5][17] != ele[11][17];
    ele[5][17] != ele[12][17];
    ele[5][17] != ele[13][17];
    ele[5][17] != ele[14][17];
    ele[5][17] != ele[15][17];
    ele[5][17] != ele[16][17];
    ele[5][17] != ele[17][17];
    ele[5][17] != ele[18][17];
    ele[5][17] != ele[19][17];
    ele[5][17] != ele[20][17];
    ele[5][17] != ele[21][17];
    ele[5][17] != ele[22][17];
    ele[5][17] != ele[23][17];
    ele[5][17] != ele[24][17];
    ele[5][17] != ele[25][17];
    ele[5][17] != ele[26][17];
    ele[5][17] != ele[27][17];
    ele[5][17] != ele[28][17];
    ele[5][17] != ele[29][17];
    ele[5][17] != ele[30][17];
    ele[5][17] != ele[31][17];
    ele[5][17] != ele[32][17];
    ele[5][17] != ele[33][17];
    ele[5][17] != ele[34][17];
    ele[5][17] != ele[35][17];
    ele[5][17] != ele[5][18];
    ele[5][17] != ele[5][19];
    ele[5][17] != ele[5][20];
    ele[5][17] != ele[5][21];
    ele[5][17] != ele[5][22];
    ele[5][17] != ele[5][23];
    ele[5][17] != ele[5][24];
    ele[5][17] != ele[5][25];
    ele[5][17] != ele[5][26];
    ele[5][17] != ele[5][27];
    ele[5][17] != ele[5][28];
    ele[5][17] != ele[5][29];
    ele[5][17] != ele[5][30];
    ele[5][17] != ele[5][31];
    ele[5][17] != ele[5][32];
    ele[5][17] != ele[5][33];
    ele[5][17] != ele[5][34];
    ele[5][17] != ele[5][35];
    ele[5][17] != ele[6][17];
    ele[5][17] != ele[7][17];
    ele[5][17] != ele[8][17];
    ele[5][17] != ele[9][17];
    ele[5][18] != ele[10][18];
    ele[5][18] != ele[11][18];
    ele[5][18] != ele[12][18];
    ele[5][18] != ele[13][18];
    ele[5][18] != ele[14][18];
    ele[5][18] != ele[15][18];
    ele[5][18] != ele[16][18];
    ele[5][18] != ele[17][18];
    ele[5][18] != ele[18][18];
    ele[5][18] != ele[19][18];
    ele[5][18] != ele[20][18];
    ele[5][18] != ele[21][18];
    ele[5][18] != ele[22][18];
    ele[5][18] != ele[23][18];
    ele[5][18] != ele[24][18];
    ele[5][18] != ele[25][18];
    ele[5][18] != ele[26][18];
    ele[5][18] != ele[27][18];
    ele[5][18] != ele[28][18];
    ele[5][18] != ele[29][18];
    ele[5][18] != ele[30][18];
    ele[5][18] != ele[31][18];
    ele[5][18] != ele[32][18];
    ele[5][18] != ele[33][18];
    ele[5][18] != ele[34][18];
    ele[5][18] != ele[35][18];
    ele[5][18] != ele[5][19];
    ele[5][18] != ele[5][20];
    ele[5][18] != ele[5][21];
    ele[5][18] != ele[5][22];
    ele[5][18] != ele[5][23];
    ele[5][18] != ele[5][24];
    ele[5][18] != ele[5][25];
    ele[5][18] != ele[5][26];
    ele[5][18] != ele[5][27];
    ele[5][18] != ele[5][28];
    ele[5][18] != ele[5][29];
    ele[5][18] != ele[5][30];
    ele[5][18] != ele[5][31];
    ele[5][18] != ele[5][32];
    ele[5][18] != ele[5][33];
    ele[5][18] != ele[5][34];
    ele[5][18] != ele[5][35];
    ele[5][18] != ele[6][18];
    ele[5][18] != ele[7][18];
    ele[5][18] != ele[8][18];
    ele[5][18] != ele[9][18];
    ele[5][19] != ele[10][19];
    ele[5][19] != ele[11][19];
    ele[5][19] != ele[12][19];
    ele[5][19] != ele[13][19];
    ele[5][19] != ele[14][19];
    ele[5][19] != ele[15][19];
    ele[5][19] != ele[16][19];
    ele[5][19] != ele[17][19];
    ele[5][19] != ele[18][19];
    ele[5][19] != ele[19][19];
    ele[5][19] != ele[20][19];
    ele[5][19] != ele[21][19];
    ele[5][19] != ele[22][19];
    ele[5][19] != ele[23][19];
    ele[5][19] != ele[24][19];
    ele[5][19] != ele[25][19];
    ele[5][19] != ele[26][19];
    ele[5][19] != ele[27][19];
    ele[5][19] != ele[28][19];
    ele[5][19] != ele[29][19];
    ele[5][19] != ele[30][19];
    ele[5][19] != ele[31][19];
    ele[5][19] != ele[32][19];
    ele[5][19] != ele[33][19];
    ele[5][19] != ele[34][19];
    ele[5][19] != ele[35][19];
    ele[5][19] != ele[5][20];
    ele[5][19] != ele[5][21];
    ele[5][19] != ele[5][22];
    ele[5][19] != ele[5][23];
    ele[5][19] != ele[5][24];
    ele[5][19] != ele[5][25];
    ele[5][19] != ele[5][26];
    ele[5][19] != ele[5][27];
    ele[5][19] != ele[5][28];
    ele[5][19] != ele[5][29];
    ele[5][19] != ele[5][30];
    ele[5][19] != ele[5][31];
    ele[5][19] != ele[5][32];
    ele[5][19] != ele[5][33];
    ele[5][19] != ele[5][34];
    ele[5][19] != ele[5][35];
    ele[5][19] != ele[6][19];
    ele[5][19] != ele[7][19];
    ele[5][19] != ele[8][19];
    ele[5][19] != ele[9][19];
    ele[5][2] != ele[10][2];
    ele[5][2] != ele[11][2];
    ele[5][2] != ele[12][2];
    ele[5][2] != ele[13][2];
    ele[5][2] != ele[14][2];
    ele[5][2] != ele[15][2];
    ele[5][2] != ele[16][2];
    ele[5][2] != ele[17][2];
    ele[5][2] != ele[18][2];
    ele[5][2] != ele[19][2];
    ele[5][2] != ele[20][2];
    ele[5][2] != ele[21][2];
    ele[5][2] != ele[22][2];
    ele[5][2] != ele[23][2];
    ele[5][2] != ele[24][2];
    ele[5][2] != ele[25][2];
    ele[5][2] != ele[26][2];
    ele[5][2] != ele[27][2];
    ele[5][2] != ele[28][2];
    ele[5][2] != ele[29][2];
    ele[5][2] != ele[30][2];
    ele[5][2] != ele[31][2];
    ele[5][2] != ele[32][2];
    ele[5][2] != ele[33][2];
    ele[5][2] != ele[34][2];
    ele[5][2] != ele[35][2];
    ele[5][2] != ele[5][10];
    ele[5][2] != ele[5][11];
    ele[5][2] != ele[5][12];
    ele[5][2] != ele[5][13];
    ele[5][2] != ele[5][14];
    ele[5][2] != ele[5][15];
    ele[5][2] != ele[5][16];
    ele[5][2] != ele[5][17];
    ele[5][2] != ele[5][18];
    ele[5][2] != ele[5][19];
    ele[5][2] != ele[5][20];
    ele[5][2] != ele[5][21];
    ele[5][2] != ele[5][22];
    ele[5][2] != ele[5][23];
    ele[5][2] != ele[5][24];
    ele[5][2] != ele[5][25];
    ele[5][2] != ele[5][26];
    ele[5][2] != ele[5][27];
    ele[5][2] != ele[5][28];
    ele[5][2] != ele[5][29];
    ele[5][2] != ele[5][3];
    ele[5][2] != ele[5][30];
    ele[5][2] != ele[5][31];
    ele[5][2] != ele[5][32];
    ele[5][2] != ele[5][33];
    ele[5][2] != ele[5][34];
    ele[5][2] != ele[5][35];
    ele[5][2] != ele[5][4];
    ele[5][2] != ele[5][5];
    ele[5][2] != ele[5][6];
    ele[5][2] != ele[5][7];
    ele[5][2] != ele[5][8];
    ele[5][2] != ele[5][9];
    ele[5][2] != ele[6][2];
    ele[5][2] != ele[7][2];
    ele[5][2] != ele[8][2];
    ele[5][2] != ele[9][2];
    ele[5][20] != ele[10][20];
    ele[5][20] != ele[11][20];
    ele[5][20] != ele[12][20];
    ele[5][20] != ele[13][20];
    ele[5][20] != ele[14][20];
    ele[5][20] != ele[15][20];
    ele[5][20] != ele[16][20];
    ele[5][20] != ele[17][20];
    ele[5][20] != ele[18][20];
    ele[5][20] != ele[19][20];
    ele[5][20] != ele[20][20];
    ele[5][20] != ele[21][20];
    ele[5][20] != ele[22][20];
    ele[5][20] != ele[23][20];
    ele[5][20] != ele[24][20];
    ele[5][20] != ele[25][20];
    ele[5][20] != ele[26][20];
    ele[5][20] != ele[27][20];
    ele[5][20] != ele[28][20];
    ele[5][20] != ele[29][20];
    ele[5][20] != ele[30][20];
    ele[5][20] != ele[31][20];
    ele[5][20] != ele[32][20];
    ele[5][20] != ele[33][20];
    ele[5][20] != ele[34][20];
    ele[5][20] != ele[35][20];
    ele[5][20] != ele[5][21];
    ele[5][20] != ele[5][22];
    ele[5][20] != ele[5][23];
    ele[5][20] != ele[5][24];
    ele[5][20] != ele[5][25];
    ele[5][20] != ele[5][26];
    ele[5][20] != ele[5][27];
    ele[5][20] != ele[5][28];
    ele[5][20] != ele[5][29];
    ele[5][20] != ele[5][30];
    ele[5][20] != ele[5][31];
    ele[5][20] != ele[5][32];
    ele[5][20] != ele[5][33];
    ele[5][20] != ele[5][34];
    ele[5][20] != ele[5][35];
    ele[5][20] != ele[6][20];
    ele[5][20] != ele[7][20];
    ele[5][20] != ele[8][20];
    ele[5][20] != ele[9][20];
    ele[5][21] != ele[10][21];
    ele[5][21] != ele[11][21];
    ele[5][21] != ele[12][21];
    ele[5][21] != ele[13][21];
    ele[5][21] != ele[14][21];
    ele[5][21] != ele[15][21];
    ele[5][21] != ele[16][21];
    ele[5][21] != ele[17][21];
    ele[5][21] != ele[18][21];
    ele[5][21] != ele[19][21];
    ele[5][21] != ele[20][21];
    ele[5][21] != ele[21][21];
    ele[5][21] != ele[22][21];
    ele[5][21] != ele[23][21];
    ele[5][21] != ele[24][21];
    ele[5][21] != ele[25][21];
    ele[5][21] != ele[26][21];
    ele[5][21] != ele[27][21];
    ele[5][21] != ele[28][21];
    ele[5][21] != ele[29][21];
    ele[5][21] != ele[30][21];
    ele[5][21] != ele[31][21];
    ele[5][21] != ele[32][21];
    ele[5][21] != ele[33][21];
    ele[5][21] != ele[34][21];
    ele[5][21] != ele[35][21];
    ele[5][21] != ele[5][22];
    ele[5][21] != ele[5][23];
    ele[5][21] != ele[5][24];
    ele[5][21] != ele[5][25];
    ele[5][21] != ele[5][26];
    ele[5][21] != ele[5][27];
    ele[5][21] != ele[5][28];
    ele[5][21] != ele[5][29];
    ele[5][21] != ele[5][30];
    ele[5][21] != ele[5][31];
    ele[5][21] != ele[5][32];
    ele[5][21] != ele[5][33];
    ele[5][21] != ele[5][34];
    ele[5][21] != ele[5][35];
    ele[5][21] != ele[6][21];
    ele[5][21] != ele[7][21];
    ele[5][21] != ele[8][21];
    ele[5][21] != ele[9][21];
    ele[5][22] != ele[10][22];
    ele[5][22] != ele[11][22];
    ele[5][22] != ele[12][22];
    ele[5][22] != ele[13][22];
    ele[5][22] != ele[14][22];
    ele[5][22] != ele[15][22];
    ele[5][22] != ele[16][22];
    ele[5][22] != ele[17][22];
    ele[5][22] != ele[18][22];
    ele[5][22] != ele[19][22];
    ele[5][22] != ele[20][22];
    ele[5][22] != ele[21][22];
    ele[5][22] != ele[22][22];
    ele[5][22] != ele[23][22];
    ele[5][22] != ele[24][22];
    ele[5][22] != ele[25][22];
    ele[5][22] != ele[26][22];
    ele[5][22] != ele[27][22];
    ele[5][22] != ele[28][22];
    ele[5][22] != ele[29][22];
    ele[5][22] != ele[30][22];
    ele[5][22] != ele[31][22];
    ele[5][22] != ele[32][22];
    ele[5][22] != ele[33][22];
    ele[5][22] != ele[34][22];
    ele[5][22] != ele[35][22];
    ele[5][22] != ele[5][23];
    ele[5][22] != ele[5][24];
    ele[5][22] != ele[5][25];
    ele[5][22] != ele[5][26];
    ele[5][22] != ele[5][27];
    ele[5][22] != ele[5][28];
    ele[5][22] != ele[5][29];
    ele[5][22] != ele[5][30];
    ele[5][22] != ele[5][31];
    ele[5][22] != ele[5][32];
    ele[5][22] != ele[5][33];
    ele[5][22] != ele[5][34];
    ele[5][22] != ele[5][35];
    ele[5][22] != ele[6][22];
    ele[5][22] != ele[7][22];
    ele[5][22] != ele[8][22];
    ele[5][22] != ele[9][22];
    ele[5][23] != ele[10][23];
    ele[5][23] != ele[11][23];
    ele[5][23] != ele[12][23];
    ele[5][23] != ele[13][23];
    ele[5][23] != ele[14][23];
    ele[5][23] != ele[15][23];
    ele[5][23] != ele[16][23];
    ele[5][23] != ele[17][23];
    ele[5][23] != ele[18][23];
    ele[5][23] != ele[19][23];
    ele[5][23] != ele[20][23];
    ele[5][23] != ele[21][23];
    ele[5][23] != ele[22][23];
    ele[5][23] != ele[23][23];
    ele[5][23] != ele[24][23];
    ele[5][23] != ele[25][23];
    ele[5][23] != ele[26][23];
    ele[5][23] != ele[27][23];
    ele[5][23] != ele[28][23];
    ele[5][23] != ele[29][23];
    ele[5][23] != ele[30][23];
    ele[5][23] != ele[31][23];
    ele[5][23] != ele[32][23];
    ele[5][23] != ele[33][23];
    ele[5][23] != ele[34][23];
    ele[5][23] != ele[35][23];
    ele[5][23] != ele[5][24];
    ele[5][23] != ele[5][25];
    ele[5][23] != ele[5][26];
    ele[5][23] != ele[5][27];
    ele[5][23] != ele[5][28];
    ele[5][23] != ele[5][29];
    ele[5][23] != ele[5][30];
    ele[5][23] != ele[5][31];
    ele[5][23] != ele[5][32];
    ele[5][23] != ele[5][33];
    ele[5][23] != ele[5][34];
    ele[5][23] != ele[5][35];
    ele[5][23] != ele[6][23];
    ele[5][23] != ele[7][23];
    ele[5][23] != ele[8][23];
    ele[5][23] != ele[9][23];
    ele[5][24] != ele[10][24];
    ele[5][24] != ele[11][24];
    ele[5][24] != ele[12][24];
    ele[5][24] != ele[13][24];
    ele[5][24] != ele[14][24];
    ele[5][24] != ele[15][24];
    ele[5][24] != ele[16][24];
    ele[5][24] != ele[17][24];
    ele[5][24] != ele[18][24];
    ele[5][24] != ele[19][24];
    ele[5][24] != ele[20][24];
    ele[5][24] != ele[21][24];
    ele[5][24] != ele[22][24];
    ele[5][24] != ele[23][24];
    ele[5][24] != ele[24][24];
    ele[5][24] != ele[25][24];
    ele[5][24] != ele[26][24];
    ele[5][24] != ele[27][24];
    ele[5][24] != ele[28][24];
    ele[5][24] != ele[29][24];
    ele[5][24] != ele[30][24];
    ele[5][24] != ele[31][24];
    ele[5][24] != ele[32][24];
    ele[5][24] != ele[33][24];
    ele[5][24] != ele[34][24];
    ele[5][24] != ele[35][24];
    ele[5][24] != ele[5][25];
    ele[5][24] != ele[5][26];
    ele[5][24] != ele[5][27];
    ele[5][24] != ele[5][28];
    ele[5][24] != ele[5][29];
    ele[5][24] != ele[5][30];
    ele[5][24] != ele[5][31];
    ele[5][24] != ele[5][32];
    ele[5][24] != ele[5][33];
    ele[5][24] != ele[5][34];
    ele[5][24] != ele[5][35];
    ele[5][24] != ele[6][24];
    ele[5][24] != ele[7][24];
    ele[5][24] != ele[8][24];
    ele[5][24] != ele[9][24];
    ele[5][25] != ele[10][25];
    ele[5][25] != ele[11][25];
    ele[5][25] != ele[12][25];
    ele[5][25] != ele[13][25];
    ele[5][25] != ele[14][25];
    ele[5][25] != ele[15][25];
    ele[5][25] != ele[16][25];
    ele[5][25] != ele[17][25];
    ele[5][25] != ele[18][25];
    ele[5][25] != ele[19][25];
    ele[5][25] != ele[20][25];
    ele[5][25] != ele[21][25];
    ele[5][25] != ele[22][25];
    ele[5][25] != ele[23][25];
    ele[5][25] != ele[24][25];
    ele[5][25] != ele[25][25];
    ele[5][25] != ele[26][25];
    ele[5][25] != ele[27][25];
    ele[5][25] != ele[28][25];
    ele[5][25] != ele[29][25];
    ele[5][25] != ele[30][25];
    ele[5][25] != ele[31][25];
    ele[5][25] != ele[32][25];
    ele[5][25] != ele[33][25];
    ele[5][25] != ele[34][25];
    ele[5][25] != ele[35][25];
    ele[5][25] != ele[5][26];
    ele[5][25] != ele[5][27];
    ele[5][25] != ele[5][28];
    ele[5][25] != ele[5][29];
    ele[5][25] != ele[5][30];
    ele[5][25] != ele[5][31];
    ele[5][25] != ele[5][32];
    ele[5][25] != ele[5][33];
    ele[5][25] != ele[5][34];
    ele[5][25] != ele[5][35];
    ele[5][25] != ele[6][25];
    ele[5][25] != ele[7][25];
    ele[5][25] != ele[8][25];
    ele[5][25] != ele[9][25];
    ele[5][26] != ele[10][26];
    ele[5][26] != ele[11][26];
    ele[5][26] != ele[12][26];
    ele[5][26] != ele[13][26];
    ele[5][26] != ele[14][26];
    ele[5][26] != ele[15][26];
    ele[5][26] != ele[16][26];
    ele[5][26] != ele[17][26];
    ele[5][26] != ele[18][26];
    ele[5][26] != ele[19][26];
    ele[5][26] != ele[20][26];
    ele[5][26] != ele[21][26];
    ele[5][26] != ele[22][26];
    ele[5][26] != ele[23][26];
    ele[5][26] != ele[24][26];
    ele[5][26] != ele[25][26];
    ele[5][26] != ele[26][26];
    ele[5][26] != ele[27][26];
    ele[5][26] != ele[28][26];
    ele[5][26] != ele[29][26];
    ele[5][26] != ele[30][26];
    ele[5][26] != ele[31][26];
    ele[5][26] != ele[32][26];
    ele[5][26] != ele[33][26];
    ele[5][26] != ele[34][26];
    ele[5][26] != ele[35][26];
    ele[5][26] != ele[5][27];
    ele[5][26] != ele[5][28];
    ele[5][26] != ele[5][29];
    ele[5][26] != ele[5][30];
    ele[5][26] != ele[5][31];
    ele[5][26] != ele[5][32];
    ele[5][26] != ele[5][33];
    ele[5][26] != ele[5][34];
    ele[5][26] != ele[5][35];
    ele[5][26] != ele[6][26];
    ele[5][26] != ele[7][26];
    ele[5][26] != ele[8][26];
    ele[5][26] != ele[9][26];
    ele[5][27] != ele[10][27];
    ele[5][27] != ele[11][27];
    ele[5][27] != ele[12][27];
    ele[5][27] != ele[13][27];
    ele[5][27] != ele[14][27];
    ele[5][27] != ele[15][27];
    ele[5][27] != ele[16][27];
    ele[5][27] != ele[17][27];
    ele[5][27] != ele[18][27];
    ele[5][27] != ele[19][27];
    ele[5][27] != ele[20][27];
    ele[5][27] != ele[21][27];
    ele[5][27] != ele[22][27];
    ele[5][27] != ele[23][27];
    ele[5][27] != ele[24][27];
    ele[5][27] != ele[25][27];
    ele[5][27] != ele[26][27];
    ele[5][27] != ele[27][27];
    ele[5][27] != ele[28][27];
    ele[5][27] != ele[29][27];
    ele[5][27] != ele[30][27];
    ele[5][27] != ele[31][27];
    ele[5][27] != ele[32][27];
    ele[5][27] != ele[33][27];
    ele[5][27] != ele[34][27];
    ele[5][27] != ele[35][27];
    ele[5][27] != ele[5][28];
    ele[5][27] != ele[5][29];
    ele[5][27] != ele[5][30];
    ele[5][27] != ele[5][31];
    ele[5][27] != ele[5][32];
    ele[5][27] != ele[5][33];
    ele[5][27] != ele[5][34];
    ele[5][27] != ele[5][35];
    ele[5][27] != ele[6][27];
    ele[5][27] != ele[7][27];
    ele[5][27] != ele[8][27];
    ele[5][27] != ele[9][27];
    ele[5][28] != ele[10][28];
    ele[5][28] != ele[11][28];
    ele[5][28] != ele[12][28];
    ele[5][28] != ele[13][28];
    ele[5][28] != ele[14][28];
    ele[5][28] != ele[15][28];
    ele[5][28] != ele[16][28];
    ele[5][28] != ele[17][28];
    ele[5][28] != ele[18][28];
    ele[5][28] != ele[19][28];
    ele[5][28] != ele[20][28];
    ele[5][28] != ele[21][28];
    ele[5][28] != ele[22][28];
    ele[5][28] != ele[23][28];
    ele[5][28] != ele[24][28];
    ele[5][28] != ele[25][28];
    ele[5][28] != ele[26][28];
    ele[5][28] != ele[27][28];
    ele[5][28] != ele[28][28];
    ele[5][28] != ele[29][28];
    ele[5][28] != ele[30][28];
    ele[5][28] != ele[31][28];
    ele[5][28] != ele[32][28];
    ele[5][28] != ele[33][28];
    ele[5][28] != ele[34][28];
    ele[5][28] != ele[35][28];
    ele[5][28] != ele[5][29];
    ele[5][28] != ele[5][30];
    ele[5][28] != ele[5][31];
    ele[5][28] != ele[5][32];
    ele[5][28] != ele[5][33];
    ele[5][28] != ele[5][34];
    ele[5][28] != ele[5][35];
    ele[5][28] != ele[6][28];
    ele[5][28] != ele[7][28];
    ele[5][28] != ele[8][28];
    ele[5][28] != ele[9][28];
    ele[5][29] != ele[10][29];
    ele[5][29] != ele[11][29];
    ele[5][29] != ele[12][29];
    ele[5][29] != ele[13][29];
    ele[5][29] != ele[14][29];
    ele[5][29] != ele[15][29];
    ele[5][29] != ele[16][29];
    ele[5][29] != ele[17][29];
    ele[5][29] != ele[18][29];
    ele[5][29] != ele[19][29];
    ele[5][29] != ele[20][29];
    ele[5][29] != ele[21][29];
    ele[5][29] != ele[22][29];
    ele[5][29] != ele[23][29];
    ele[5][29] != ele[24][29];
    ele[5][29] != ele[25][29];
    ele[5][29] != ele[26][29];
    ele[5][29] != ele[27][29];
    ele[5][29] != ele[28][29];
    ele[5][29] != ele[29][29];
    ele[5][29] != ele[30][29];
    ele[5][29] != ele[31][29];
    ele[5][29] != ele[32][29];
    ele[5][29] != ele[33][29];
    ele[5][29] != ele[34][29];
    ele[5][29] != ele[35][29];
    ele[5][29] != ele[5][30];
    ele[5][29] != ele[5][31];
    ele[5][29] != ele[5][32];
    ele[5][29] != ele[5][33];
    ele[5][29] != ele[5][34];
    ele[5][29] != ele[5][35];
    ele[5][29] != ele[6][29];
    ele[5][29] != ele[7][29];
    ele[5][29] != ele[8][29];
    ele[5][29] != ele[9][29];
    ele[5][3] != ele[10][3];
    ele[5][3] != ele[11][3];
    ele[5][3] != ele[12][3];
    ele[5][3] != ele[13][3];
    ele[5][3] != ele[14][3];
    ele[5][3] != ele[15][3];
    ele[5][3] != ele[16][3];
    ele[5][3] != ele[17][3];
    ele[5][3] != ele[18][3];
    ele[5][3] != ele[19][3];
    ele[5][3] != ele[20][3];
    ele[5][3] != ele[21][3];
    ele[5][3] != ele[22][3];
    ele[5][3] != ele[23][3];
    ele[5][3] != ele[24][3];
    ele[5][3] != ele[25][3];
    ele[5][3] != ele[26][3];
    ele[5][3] != ele[27][3];
    ele[5][3] != ele[28][3];
    ele[5][3] != ele[29][3];
    ele[5][3] != ele[30][3];
    ele[5][3] != ele[31][3];
    ele[5][3] != ele[32][3];
    ele[5][3] != ele[33][3];
    ele[5][3] != ele[34][3];
    ele[5][3] != ele[35][3];
    ele[5][3] != ele[5][10];
    ele[5][3] != ele[5][11];
    ele[5][3] != ele[5][12];
    ele[5][3] != ele[5][13];
    ele[5][3] != ele[5][14];
    ele[5][3] != ele[5][15];
    ele[5][3] != ele[5][16];
    ele[5][3] != ele[5][17];
    ele[5][3] != ele[5][18];
    ele[5][3] != ele[5][19];
    ele[5][3] != ele[5][20];
    ele[5][3] != ele[5][21];
    ele[5][3] != ele[5][22];
    ele[5][3] != ele[5][23];
    ele[5][3] != ele[5][24];
    ele[5][3] != ele[5][25];
    ele[5][3] != ele[5][26];
    ele[5][3] != ele[5][27];
    ele[5][3] != ele[5][28];
    ele[5][3] != ele[5][29];
    ele[5][3] != ele[5][30];
    ele[5][3] != ele[5][31];
    ele[5][3] != ele[5][32];
    ele[5][3] != ele[5][33];
    ele[5][3] != ele[5][34];
    ele[5][3] != ele[5][35];
    ele[5][3] != ele[5][4];
    ele[5][3] != ele[5][5];
    ele[5][3] != ele[5][6];
    ele[5][3] != ele[5][7];
    ele[5][3] != ele[5][8];
    ele[5][3] != ele[5][9];
    ele[5][3] != ele[6][3];
    ele[5][3] != ele[7][3];
    ele[5][3] != ele[8][3];
    ele[5][3] != ele[9][3];
    ele[5][30] != ele[10][30];
    ele[5][30] != ele[11][30];
    ele[5][30] != ele[12][30];
    ele[5][30] != ele[13][30];
    ele[5][30] != ele[14][30];
    ele[5][30] != ele[15][30];
    ele[5][30] != ele[16][30];
    ele[5][30] != ele[17][30];
    ele[5][30] != ele[18][30];
    ele[5][30] != ele[19][30];
    ele[5][30] != ele[20][30];
    ele[5][30] != ele[21][30];
    ele[5][30] != ele[22][30];
    ele[5][30] != ele[23][30];
    ele[5][30] != ele[24][30];
    ele[5][30] != ele[25][30];
    ele[5][30] != ele[26][30];
    ele[5][30] != ele[27][30];
    ele[5][30] != ele[28][30];
    ele[5][30] != ele[29][30];
    ele[5][30] != ele[30][30];
    ele[5][30] != ele[31][30];
    ele[5][30] != ele[32][30];
    ele[5][30] != ele[33][30];
    ele[5][30] != ele[34][30];
    ele[5][30] != ele[35][30];
    ele[5][30] != ele[5][31];
    ele[5][30] != ele[5][32];
    ele[5][30] != ele[5][33];
    ele[5][30] != ele[5][34];
    ele[5][30] != ele[5][35];
    ele[5][30] != ele[6][30];
    ele[5][30] != ele[7][30];
    ele[5][30] != ele[8][30];
    ele[5][30] != ele[9][30];
    ele[5][31] != ele[10][31];
    ele[5][31] != ele[11][31];
    ele[5][31] != ele[12][31];
    ele[5][31] != ele[13][31];
    ele[5][31] != ele[14][31];
    ele[5][31] != ele[15][31];
    ele[5][31] != ele[16][31];
    ele[5][31] != ele[17][31];
    ele[5][31] != ele[18][31];
    ele[5][31] != ele[19][31];
    ele[5][31] != ele[20][31];
    ele[5][31] != ele[21][31];
    ele[5][31] != ele[22][31];
    ele[5][31] != ele[23][31];
    ele[5][31] != ele[24][31];
    ele[5][31] != ele[25][31];
    ele[5][31] != ele[26][31];
    ele[5][31] != ele[27][31];
    ele[5][31] != ele[28][31];
    ele[5][31] != ele[29][31];
    ele[5][31] != ele[30][31];
    ele[5][31] != ele[31][31];
    ele[5][31] != ele[32][31];
    ele[5][31] != ele[33][31];
    ele[5][31] != ele[34][31];
    ele[5][31] != ele[35][31];
    ele[5][31] != ele[5][32];
    ele[5][31] != ele[5][33];
    ele[5][31] != ele[5][34];
    ele[5][31] != ele[5][35];
    ele[5][31] != ele[6][31];
    ele[5][31] != ele[7][31];
    ele[5][31] != ele[8][31];
    ele[5][31] != ele[9][31];
    ele[5][32] != ele[10][32];
    ele[5][32] != ele[11][32];
    ele[5][32] != ele[12][32];
    ele[5][32] != ele[13][32];
    ele[5][32] != ele[14][32];
    ele[5][32] != ele[15][32];
    ele[5][32] != ele[16][32];
    ele[5][32] != ele[17][32];
    ele[5][32] != ele[18][32];
    ele[5][32] != ele[19][32];
    ele[5][32] != ele[20][32];
    ele[5][32] != ele[21][32];
    ele[5][32] != ele[22][32];
    ele[5][32] != ele[23][32];
    ele[5][32] != ele[24][32];
    ele[5][32] != ele[25][32];
    ele[5][32] != ele[26][32];
    ele[5][32] != ele[27][32];
    ele[5][32] != ele[28][32];
    ele[5][32] != ele[29][32];
    ele[5][32] != ele[30][32];
    ele[5][32] != ele[31][32];
    ele[5][32] != ele[32][32];
    ele[5][32] != ele[33][32];
    ele[5][32] != ele[34][32];
    ele[5][32] != ele[35][32];
    ele[5][32] != ele[5][33];
    ele[5][32] != ele[5][34];
    ele[5][32] != ele[5][35];
    ele[5][32] != ele[6][32];
    ele[5][32] != ele[7][32];
    ele[5][32] != ele[8][32];
    ele[5][32] != ele[9][32];
    ele[5][33] != ele[10][33];
    ele[5][33] != ele[11][33];
    ele[5][33] != ele[12][33];
    ele[5][33] != ele[13][33];
    ele[5][33] != ele[14][33];
    ele[5][33] != ele[15][33];
    ele[5][33] != ele[16][33];
    ele[5][33] != ele[17][33];
    ele[5][33] != ele[18][33];
    ele[5][33] != ele[19][33];
    ele[5][33] != ele[20][33];
    ele[5][33] != ele[21][33];
    ele[5][33] != ele[22][33];
    ele[5][33] != ele[23][33];
    ele[5][33] != ele[24][33];
    ele[5][33] != ele[25][33];
    ele[5][33] != ele[26][33];
    ele[5][33] != ele[27][33];
    ele[5][33] != ele[28][33];
    ele[5][33] != ele[29][33];
    ele[5][33] != ele[30][33];
    ele[5][33] != ele[31][33];
    ele[5][33] != ele[32][33];
    ele[5][33] != ele[33][33];
    ele[5][33] != ele[34][33];
    ele[5][33] != ele[35][33];
    ele[5][33] != ele[5][34];
    ele[5][33] != ele[5][35];
    ele[5][33] != ele[6][33];
    ele[5][33] != ele[7][33];
    ele[5][33] != ele[8][33];
    ele[5][33] != ele[9][33];
    ele[5][34] != ele[10][34];
    ele[5][34] != ele[11][34];
    ele[5][34] != ele[12][34];
    ele[5][34] != ele[13][34];
    ele[5][34] != ele[14][34];
    ele[5][34] != ele[15][34];
    ele[5][34] != ele[16][34];
    ele[5][34] != ele[17][34];
    ele[5][34] != ele[18][34];
    ele[5][34] != ele[19][34];
    ele[5][34] != ele[20][34];
    ele[5][34] != ele[21][34];
    ele[5][34] != ele[22][34];
    ele[5][34] != ele[23][34];
    ele[5][34] != ele[24][34];
    ele[5][34] != ele[25][34];
    ele[5][34] != ele[26][34];
    ele[5][34] != ele[27][34];
    ele[5][34] != ele[28][34];
    ele[5][34] != ele[29][34];
    ele[5][34] != ele[30][34];
    ele[5][34] != ele[31][34];
    ele[5][34] != ele[32][34];
    ele[5][34] != ele[33][34];
    ele[5][34] != ele[34][34];
    ele[5][34] != ele[35][34];
    ele[5][34] != ele[5][35];
    ele[5][34] != ele[6][34];
    ele[5][34] != ele[7][34];
    ele[5][34] != ele[8][34];
    ele[5][34] != ele[9][34];
    ele[5][35] != ele[10][35];
    ele[5][35] != ele[11][35];
    ele[5][35] != ele[12][35];
    ele[5][35] != ele[13][35];
    ele[5][35] != ele[14][35];
    ele[5][35] != ele[15][35];
    ele[5][35] != ele[16][35];
    ele[5][35] != ele[17][35];
    ele[5][35] != ele[18][35];
    ele[5][35] != ele[19][35];
    ele[5][35] != ele[20][35];
    ele[5][35] != ele[21][35];
    ele[5][35] != ele[22][35];
    ele[5][35] != ele[23][35];
    ele[5][35] != ele[24][35];
    ele[5][35] != ele[25][35];
    ele[5][35] != ele[26][35];
    ele[5][35] != ele[27][35];
    ele[5][35] != ele[28][35];
    ele[5][35] != ele[29][35];
    ele[5][35] != ele[30][35];
    ele[5][35] != ele[31][35];
    ele[5][35] != ele[32][35];
    ele[5][35] != ele[33][35];
    ele[5][35] != ele[34][35];
    ele[5][35] != ele[35][35];
    ele[5][35] != ele[6][35];
    ele[5][35] != ele[7][35];
    ele[5][35] != ele[8][35];
    ele[5][35] != ele[9][35];
    ele[5][4] != ele[10][4];
    ele[5][4] != ele[11][4];
    ele[5][4] != ele[12][4];
    ele[5][4] != ele[13][4];
    ele[5][4] != ele[14][4];
    ele[5][4] != ele[15][4];
    ele[5][4] != ele[16][4];
    ele[5][4] != ele[17][4];
    ele[5][4] != ele[18][4];
    ele[5][4] != ele[19][4];
    ele[5][4] != ele[20][4];
    ele[5][4] != ele[21][4];
    ele[5][4] != ele[22][4];
    ele[5][4] != ele[23][4];
    ele[5][4] != ele[24][4];
    ele[5][4] != ele[25][4];
    ele[5][4] != ele[26][4];
    ele[5][4] != ele[27][4];
    ele[5][4] != ele[28][4];
    ele[5][4] != ele[29][4];
    ele[5][4] != ele[30][4];
    ele[5][4] != ele[31][4];
    ele[5][4] != ele[32][4];
    ele[5][4] != ele[33][4];
    ele[5][4] != ele[34][4];
    ele[5][4] != ele[35][4];
    ele[5][4] != ele[5][10];
    ele[5][4] != ele[5][11];
    ele[5][4] != ele[5][12];
    ele[5][4] != ele[5][13];
    ele[5][4] != ele[5][14];
    ele[5][4] != ele[5][15];
    ele[5][4] != ele[5][16];
    ele[5][4] != ele[5][17];
    ele[5][4] != ele[5][18];
    ele[5][4] != ele[5][19];
    ele[5][4] != ele[5][20];
    ele[5][4] != ele[5][21];
    ele[5][4] != ele[5][22];
    ele[5][4] != ele[5][23];
    ele[5][4] != ele[5][24];
    ele[5][4] != ele[5][25];
    ele[5][4] != ele[5][26];
    ele[5][4] != ele[5][27];
    ele[5][4] != ele[5][28];
    ele[5][4] != ele[5][29];
    ele[5][4] != ele[5][30];
    ele[5][4] != ele[5][31];
    ele[5][4] != ele[5][32];
    ele[5][4] != ele[5][33];
    ele[5][4] != ele[5][34];
    ele[5][4] != ele[5][35];
    ele[5][4] != ele[5][5];
    ele[5][4] != ele[5][6];
    ele[5][4] != ele[5][7];
    ele[5][4] != ele[5][8];
    ele[5][4] != ele[5][9];
    ele[5][4] != ele[6][4];
    ele[5][4] != ele[7][4];
    ele[5][4] != ele[8][4];
    ele[5][4] != ele[9][4];
    ele[5][5] != ele[10][5];
    ele[5][5] != ele[11][5];
    ele[5][5] != ele[12][5];
    ele[5][5] != ele[13][5];
    ele[5][5] != ele[14][5];
    ele[5][5] != ele[15][5];
    ele[5][5] != ele[16][5];
    ele[5][5] != ele[17][5];
    ele[5][5] != ele[18][5];
    ele[5][5] != ele[19][5];
    ele[5][5] != ele[20][5];
    ele[5][5] != ele[21][5];
    ele[5][5] != ele[22][5];
    ele[5][5] != ele[23][5];
    ele[5][5] != ele[24][5];
    ele[5][5] != ele[25][5];
    ele[5][5] != ele[26][5];
    ele[5][5] != ele[27][5];
    ele[5][5] != ele[28][5];
    ele[5][5] != ele[29][5];
    ele[5][5] != ele[30][5];
    ele[5][5] != ele[31][5];
    ele[5][5] != ele[32][5];
    ele[5][5] != ele[33][5];
    ele[5][5] != ele[34][5];
    ele[5][5] != ele[35][5];
    ele[5][5] != ele[5][10];
    ele[5][5] != ele[5][11];
    ele[5][5] != ele[5][12];
    ele[5][5] != ele[5][13];
    ele[5][5] != ele[5][14];
    ele[5][5] != ele[5][15];
    ele[5][5] != ele[5][16];
    ele[5][5] != ele[5][17];
    ele[5][5] != ele[5][18];
    ele[5][5] != ele[5][19];
    ele[5][5] != ele[5][20];
    ele[5][5] != ele[5][21];
    ele[5][5] != ele[5][22];
    ele[5][5] != ele[5][23];
    ele[5][5] != ele[5][24];
    ele[5][5] != ele[5][25];
    ele[5][5] != ele[5][26];
    ele[5][5] != ele[5][27];
    ele[5][5] != ele[5][28];
    ele[5][5] != ele[5][29];
    ele[5][5] != ele[5][30];
    ele[5][5] != ele[5][31];
    ele[5][5] != ele[5][32];
    ele[5][5] != ele[5][33];
    ele[5][5] != ele[5][34];
    ele[5][5] != ele[5][35];
    ele[5][5] != ele[5][6];
    ele[5][5] != ele[5][7];
    ele[5][5] != ele[5][8];
    ele[5][5] != ele[5][9];
    ele[5][5] != ele[6][5];
    ele[5][5] != ele[7][5];
    ele[5][5] != ele[8][5];
    ele[5][5] != ele[9][5];
    ele[5][6] != ele[10][6];
    ele[5][6] != ele[11][6];
    ele[5][6] != ele[12][6];
    ele[5][6] != ele[13][6];
    ele[5][6] != ele[14][6];
    ele[5][6] != ele[15][6];
    ele[5][6] != ele[16][6];
    ele[5][6] != ele[17][6];
    ele[5][6] != ele[18][6];
    ele[5][6] != ele[19][6];
    ele[5][6] != ele[20][6];
    ele[5][6] != ele[21][6];
    ele[5][6] != ele[22][6];
    ele[5][6] != ele[23][6];
    ele[5][6] != ele[24][6];
    ele[5][6] != ele[25][6];
    ele[5][6] != ele[26][6];
    ele[5][6] != ele[27][6];
    ele[5][6] != ele[28][6];
    ele[5][6] != ele[29][6];
    ele[5][6] != ele[30][6];
    ele[5][6] != ele[31][6];
    ele[5][6] != ele[32][6];
    ele[5][6] != ele[33][6];
    ele[5][6] != ele[34][6];
    ele[5][6] != ele[35][6];
    ele[5][6] != ele[5][10];
    ele[5][6] != ele[5][11];
    ele[5][6] != ele[5][12];
    ele[5][6] != ele[5][13];
    ele[5][6] != ele[5][14];
    ele[5][6] != ele[5][15];
    ele[5][6] != ele[5][16];
    ele[5][6] != ele[5][17];
    ele[5][6] != ele[5][18];
    ele[5][6] != ele[5][19];
    ele[5][6] != ele[5][20];
    ele[5][6] != ele[5][21];
    ele[5][6] != ele[5][22];
    ele[5][6] != ele[5][23];
    ele[5][6] != ele[5][24];
    ele[5][6] != ele[5][25];
    ele[5][6] != ele[5][26];
    ele[5][6] != ele[5][27];
    ele[5][6] != ele[5][28];
    ele[5][6] != ele[5][29];
    ele[5][6] != ele[5][30];
    ele[5][6] != ele[5][31];
    ele[5][6] != ele[5][32];
    ele[5][6] != ele[5][33];
    ele[5][6] != ele[5][34];
    ele[5][6] != ele[5][35];
    ele[5][6] != ele[5][7];
    ele[5][6] != ele[5][8];
    ele[5][6] != ele[5][9];
    ele[5][6] != ele[6][6];
    ele[5][6] != ele[7][6];
    ele[5][6] != ele[8][6];
    ele[5][6] != ele[9][6];
    ele[5][7] != ele[10][7];
    ele[5][7] != ele[11][7];
    ele[5][7] != ele[12][7];
    ele[5][7] != ele[13][7];
    ele[5][7] != ele[14][7];
    ele[5][7] != ele[15][7];
    ele[5][7] != ele[16][7];
    ele[5][7] != ele[17][7];
    ele[5][7] != ele[18][7];
    ele[5][7] != ele[19][7];
    ele[5][7] != ele[20][7];
    ele[5][7] != ele[21][7];
    ele[5][7] != ele[22][7];
    ele[5][7] != ele[23][7];
    ele[5][7] != ele[24][7];
    ele[5][7] != ele[25][7];
    ele[5][7] != ele[26][7];
    ele[5][7] != ele[27][7];
    ele[5][7] != ele[28][7];
    ele[5][7] != ele[29][7];
    ele[5][7] != ele[30][7];
    ele[5][7] != ele[31][7];
    ele[5][7] != ele[32][7];
    ele[5][7] != ele[33][7];
    ele[5][7] != ele[34][7];
    ele[5][7] != ele[35][7];
    ele[5][7] != ele[5][10];
    ele[5][7] != ele[5][11];
    ele[5][7] != ele[5][12];
    ele[5][7] != ele[5][13];
    ele[5][7] != ele[5][14];
    ele[5][7] != ele[5][15];
    ele[5][7] != ele[5][16];
    ele[5][7] != ele[5][17];
    ele[5][7] != ele[5][18];
    ele[5][7] != ele[5][19];
    ele[5][7] != ele[5][20];
    ele[5][7] != ele[5][21];
    ele[5][7] != ele[5][22];
    ele[5][7] != ele[5][23];
    ele[5][7] != ele[5][24];
    ele[5][7] != ele[5][25];
    ele[5][7] != ele[5][26];
    ele[5][7] != ele[5][27];
    ele[5][7] != ele[5][28];
    ele[5][7] != ele[5][29];
    ele[5][7] != ele[5][30];
    ele[5][7] != ele[5][31];
    ele[5][7] != ele[5][32];
    ele[5][7] != ele[5][33];
    ele[5][7] != ele[5][34];
    ele[5][7] != ele[5][35];
    ele[5][7] != ele[5][8];
    ele[5][7] != ele[5][9];
    ele[5][7] != ele[6][7];
    ele[5][7] != ele[7][7];
    ele[5][7] != ele[8][7];
    ele[5][7] != ele[9][7];
    ele[5][8] != ele[10][8];
    ele[5][8] != ele[11][8];
    ele[5][8] != ele[12][8];
    ele[5][8] != ele[13][8];
    ele[5][8] != ele[14][8];
    ele[5][8] != ele[15][8];
    ele[5][8] != ele[16][8];
    ele[5][8] != ele[17][8];
    ele[5][8] != ele[18][8];
    ele[5][8] != ele[19][8];
    ele[5][8] != ele[20][8];
    ele[5][8] != ele[21][8];
    ele[5][8] != ele[22][8];
    ele[5][8] != ele[23][8];
    ele[5][8] != ele[24][8];
    ele[5][8] != ele[25][8];
    ele[5][8] != ele[26][8];
    ele[5][8] != ele[27][8];
    ele[5][8] != ele[28][8];
    ele[5][8] != ele[29][8];
    ele[5][8] != ele[30][8];
    ele[5][8] != ele[31][8];
    ele[5][8] != ele[32][8];
    ele[5][8] != ele[33][8];
    ele[5][8] != ele[34][8];
    ele[5][8] != ele[35][8];
    ele[5][8] != ele[5][10];
    ele[5][8] != ele[5][11];
    ele[5][8] != ele[5][12];
    ele[5][8] != ele[5][13];
    ele[5][8] != ele[5][14];
    ele[5][8] != ele[5][15];
    ele[5][8] != ele[5][16];
    ele[5][8] != ele[5][17];
    ele[5][8] != ele[5][18];
    ele[5][8] != ele[5][19];
    ele[5][8] != ele[5][20];
    ele[5][8] != ele[5][21];
    ele[5][8] != ele[5][22];
    ele[5][8] != ele[5][23];
    ele[5][8] != ele[5][24];
    ele[5][8] != ele[5][25];
    ele[5][8] != ele[5][26];
    ele[5][8] != ele[5][27];
    ele[5][8] != ele[5][28];
    ele[5][8] != ele[5][29];
    ele[5][8] != ele[5][30];
    ele[5][8] != ele[5][31];
    ele[5][8] != ele[5][32];
    ele[5][8] != ele[5][33];
    ele[5][8] != ele[5][34];
    ele[5][8] != ele[5][35];
    ele[5][8] != ele[5][9];
    ele[5][8] != ele[6][8];
    ele[5][8] != ele[7][8];
    ele[5][8] != ele[8][8];
    ele[5][8] != ele[9][8];
    ele[5][9] != ele[10][9];
    ele[5][9] != ele[11][9];
    ele[5][9] != ele[12][9];
    ele[5][9] != ele[13][9];
    ele[5][9] != ele[14][9];
    ele[5][9] != ele[15][9];
    ele[5][9] != ele[16][9];
    ele[5][9] != ele[17][9];
    ele[5][9] != ele[18][9];
    ele[5][9] != ele[19][9];
    ele[5][9] != ele[20][9];
    ele[5][9] != ele[21][9];
    ele[5][9] != ele[22][9];
    ele[5][9] != ele[23][9];
    ele[5][9] != ele[24][9];
    ele[5][9] != ele[25][9];
    ele[5][9] != ele[26][9];
    ele[5][9] != ele[27][9];
    ele[5][9] != ele[28][9];
    ele[5][9] != ele[29][9];
    ele[5][9] != ele[30][9];
    ele[5][9] != ele[31][9];
    ele[5][9] != ele[32][9];
    ele[5][9] != ele[33][9];
    ele[5][9] != ele[34][9];
    ele[5][9] != ele[35][9];
    ele[5][9] != ele[5][10];
    ele[5][9] != ele[5][11];
    ele[5][9] != ele[5][12];
    ele[5][9] != ele[5][13];
    ele[5][9] != ele[5][14];
    ele[5][9] != ele[5][15];
    ele[5][9] != ele[5][16];
    ele[5][9] != ele[5][17];
    ele[5][9] != ele[5][18];
    ele[5][9] != ele[5][19];
    ele[5][9] != ele[5][20];
    ele[5][9] != ele[5][21];
    ele[5][9] != ele[5][22];
    ele[5][9] != ele[5][23];
    ele[5][9] != ele[5][24];
    ele[5][9] != ele[5][25];
    ele[5][9] != ele[5][26];
    ele[5][9] != ele[5][27];
    ele[5][9] != ele[5][28];
    ele[5][9] != ele[5][29];
    ele[5][9] != ele[5][30];
    ele[5][9] != ele[5][31];
    ele[5][9] != ele[5][32];
    ele[5][9] != ele[5][33];
    ele[5][9] != ele[5][34];
    ele[5][9] != ele[5][35];
    ele[5][9] != ele[6][9];
    ele[5][9] != ele[7][9];
    ele[5][9] != ele[8][9];
    ele[5][9] != ele[9][9];
    ele[6][0] != ele[10][0];
    ele[6][0] != ele[10][1];
    ele[6][0] != ele[10][2];
    ele[6][0] != ele[10][3];
    ele[6][0] != ele[10][4];
    ele[6][0] != ele[10][5];
    ele[6][0] != ele[11][0];
    ele[6][0] != ele[11][1];
    ele[6][0] != ele[11][2];
    ele[6][0] != ele[11][3];
    ele[6][0] != ele[11][4];
    ele[6][0] != ele[11][5];
    ele[6][0] != ele[12][0];
    ele[6][0] != ele[13][0];
    ele[6][0] != ele[14][0];
    ele[6][0] != ele[15][0];
    ele[6][0] != ele[16][0];
    ele[6][0] != ele[17][0];
    ele[6][0] != ele[18][0];
    ele[6][0] != ele[19][0];
    ele[6][0] != ele[20][0];
    ele[6][0] != ele[21][0];
    ele[6][0] != ele[22][0];
    ele[6][0] != ele[23][0];
    ele[6][0] != ele[24][0];
    ele[6][0] != ele[25][0];
    ele[6][0] != ele[26][0];
    ele[6][0] != ele[27][0];
    ele[6][0] != ele[28][0];
    ele[6][0] != ele[29][0];
    ele[6][0] != ele[30][0];
    ele[6][0] != ele[31][0];
    ele[6][0] != ele[32][0];
    ele[6][0] != ele[33][0];
    ele[6][0] != ele[34][0];
    ele[6][0] != ele[35][0];
    ele[6][0] != ele[6][1];
    ele[6][0] != ele[6][10];
    ele[6][0] != ele[6][11];
    ele[6][0] != ele[6][12];
    ele[6][0] != ele[6][13];
    ele[6][0] != ele[6][14];
    ele[6][0] != ele[6][15];
    ele[6][0] != ele[6][16];
    ele[6][0] != ele[6][17];
    ele[6][0] != ele[6][18];
    ele[6][0] != ele[6][19];
    ele[6][0] != ele[6][2];
    ele[6][0] != ele[6][20];
    ele[6][0] != ele[6][21];
    ele[6][0] != ele[6][22];
    ele[6][0] != ele[6][23];
    ele[6][0] != ele[6][24];
    ele[6][0] != ele[6][25];
    ele[6][0] != ele[6][26];
    ele[6][0] != ele[6][27];
    ele[6][0] != ele[6][28];
    ele[6][0] != ele[6][29];
    ele[6][0] != ele[6][3];
    ele[6][0] != ele[6][30];
    ele[6][0] != ele[6][31];
    ele[6][0] != ele[6][32];
    ele[6][0] != ele[6][33];
    ele[6][0] != ele[6][34];
    ele[6][0] != ele[6][35];
    ele[6][0] != ele[6][4];
    ele[6][0] != ele[6][5];
    ele[6][0] != ele[6][6];
    ele[6][0] != ele[6][7];
    ele[6][0] != ele[6][8];
    ele[6][0] != ele[6][9];
    ele[6][0] != ele[7][0];
    ele[6][0] != ele[7][1];
    ele[6][0] != ele[7][2];
    ele[6][0] != ele[7][3];
    ele[6][0] != ele[7][4];
    ele[6][0] != ele[7][5];
    ele[6][0] != ele[8][0];
    ele[6][0] != ele[8][1];
    ele[6][0] != ele[8][2];
    ele[6][0] != ele[8][3];
    ele[6][0] != ele[8][4];
    ele[6][0] != ele[8][5];
    ele[6][0] != ele[9][0];
    ele[6][0] != ele[9][1];
    ele[6][0] != ele[9][2];
    ele[6][0] != ele[9][3];
    ele[6][0] != ele[9][4];
    ele[6][0] != ele[9][5];
    ele[6][1] != ele[10][0];
    ele[6][1] != ele[10][1];
    ele[6][1] != ele[10][2];
    ele[6][1] != ele[10][3];
    ele[6][1] != ele[10][4];
    ele[6][1] != ele[10][5];
    ele[6][1] != ele[11][0];
    ele[6][1] != ele[11][1];
    ele[6][1] != ele[11][2];
    ele[6][1] != ele[11][3];
    ele[6][1] != ele[11][4];
    ele[6][1] != ele[11][5];
    ele[6][1] != ele[12][1];
    ele[6][1] != ele[13][1];
    ele[6][1] != ele[14][1];
    ele[6][1] != ele[15][1];
    ele[6][1] != ele[16][1];
    ele[6][1] != ele[17][1];
    ele[6][1] != ele[18][1];
    ele[6][1] != ele[19][1];
    ele[6][1] != ele[20][1];
    ele[6][1] != ele[21][1];
    ele[6][1] != ele[22][1];
    ele[6][1] != ele[23][1];
    ele[6][1] != ele[24][1];
    ele[6][1] != ele[25][1];
    ele[6][1] != ele[26][1];
    ele[6][1] != ele[27][1];
    ele[6][1] != ele[28][1];
    ele[6][1] != ele[29][1];
    ele[6][1] != ele[30][1];
    ele[6][1] != ele[31][1];
    ele[6][1] != ele[32][1];
    ele[6][1] != ele[33][1];
    ele[6][1] != ele[34][1];
    ele[6][1] != ele[35][1];
    ele[6][1] != ele[6][10];
    ele[6][1] != ele[6][11];
    ele[6][1] != ele[6][12];
    ele[6][1] != ele[6][13];
    ele[6][1] != ele[6][14];
    ele[6][1] != ele[6][15];
    ele[6][1] != ele[6][16];
    ele[6][1] != ele[6][17];
    ele[6][1] != ele[6][18];
    ele[6][1] != ele[6][19];
    ele[6][1] != ele[6][2];
    ele[6][1] != ele[6][20];
    ele[6][1] != ele[6][21];
    ele[6][1] != ele[6][22];
    ele[6][1] != ele[6][23];
    ele[6][1] != ele[6][24];
    ele[6][1] != ele[6][25];
    ele[6][1] != ele[6][26];
    ele[6][1] != ele[6][27];
    ele[6][1] != ele[6][28];
    ele[6][1] != ele[6][29];
    ele[6][1] != ele[6][3];
    ele[6][1] != ele[6][30];
    ele[6][1] != ele[6][31];
    ele[6][1] != ele[6][32];
    ele[6][1] != ele[6][33];
    ele[6][1] != ele[6][34];
    ele[6][1] != ele[6][35];
    ele[6][1] != ele[6][4];
    ele[6][1] != ele[6][5];
    ele[6][1] != ele[6][6];
    ele[6][1] != ele[6][7];
    ele[6][1] != ele[6][8];
    ele[6][1] != ele[6][9];
    ele[6][1] != ele[7][0];
    ele[6][1] != ele[7][1];
    ele[6][1] != ele[7][2];
    ele[6][1] != ele[7][3];
    ele[6][1] != ele[7][4];
    ele[6][1] != ele[7][5];
    ele[6][1] != ele[8][0];
    ele[6][1] != ele[8][1];
    ele[6][1] != ele[8][2];
    ele[6][1] != ele[8][3];
    ele[6][1] != ele[8][4];
    ele[6][1] != ele[8][5];
    ele[6][1] != ele[9][0];
    ele[6][1] != ele[9][1];
    ele[6][1] != ele[9][2];
    ele[6][1] != ele[9][3];
    ele[6][1] != ele[9][4];
    ele[6][1] != ele[9][5];
    ele[6][10] != ele[10][10];
    ele[6][10] != ele[10][11];
    ele[6][10] != ele[10][6];
    ele[6][10] != ele[10][7];
    ele[6][10] != ele[10][8];
    ele[6][10] != ele[10][9];
    ele[6][10] != ele[11][10];
    ele[6][10] != ele[11][11];
    ele[6][10] != ele[11][6];
    ele[6][10] != ele[11][7];
    ele[6][10] != ele[11][8];
    ele[6][10] != ele[11][9];
    ele[6][10] != ele[12][10];
    ele[6][10] != ele[13][10];
    ele[6][10] != ele[14][10];
    ele[6][10] != ele[15][10];
    ele[6][10] != ele[16][10];
    ele[6][10] != ele[17][10];
    ele[6][10] != ele[18][10];
    ele[6][10] != ele[19][10];
    ele[6][10] != ele[20][10];
    ele[6][10] != ele[21][10];
    ele[6][10] != ele[22][10];
    ele[6][10] != ele[23][10];
    ele[6][10] != ele[24][10];
    ele[6][10] != ele[25][10];
    ele[6][10] != ele[26][10];
    ele[6][10] != ele[27][10];
    ele[6][10] != ele[28][10];
    ele[6][10] != ele[29][10];
    ele[6][10] != ele[30][10];
    ele[6][10] != ele[31][10];
    ele[6][10] != ele[32][10];
    ele[6][10] != ele[33][10];
    ele[6][10] != ele[34][10];
    ele[6][10] != ele[35][10];
    ele[6][10] != ele[6][11];
    ele[6][10] != ele[6][12];
    ele[6][10] != ele[6][13];
    ele[6][10] != ele[6][14];
    ele[6][10] != ele[6][15];
    ele[6][10] != ele[6][16];
    ele[6][10] != ele[6][17];
    ele[6][10] != ele[6][18];
    ele[6][10] != ele[6][19];
    ele[6][10] != ele[6][20];
    ele[6][10] != ele[6][21];
    ele[6][10] != ele[6][22];
    ele[6][10] != ele[6][23];
    ele[6][10] != ele[6][24];
    ele[6][10] != ele[6][25];
    ele[6][10] != ele[6][26];
    ele[6][10] != ele[6][27];
    ele[6][10] != ele[6][28];
    ele[6][10] != ele[6][29];
    ele[6][10] != ele[6][30];
    ele[6][10] != ele[6][31];
    ele[6][10] != ele[6][32];
    ele[6][10] != ele[6][33];
    ele[6][10] != ele[6][34];
    ele[6][10] != ele[6][35];
    ele[6][10] != ele[7][10];
    ele[6][10] != ele[7][11];
    ele[6][10] != ele[7][6];
    ele[6][10] != ele[7][7];
    ele[6][10] != ele[7][8];
    ele[6][10] != ele[7][9];
    ele[6][10] != ele[8][10];
    ele[6][10] != ele[8][11];
    ele[6][10] != ele[8][6];
    ele[6][10] != ele[8][7];
    ele[6][10] != ele[8][8];
    ele[6][10] != ele[8][9];
    ele[6][10] != ele[9][10];
    ele[6][10] != ele[9][11];
    ele[6][10] != ele[9][6];
    ele[6][10] != ele[9][7];
    ele[6][10] != ele[9][8];
    ele[6][10] != ele[9][9];
    ele[6][11] != ele[10][10];
    ele[6][11] != ele[10][11];
    ele[6][11] != ele[10][6];
    ele[6][11] != ele[10][7];
    ele[6][11] != ele[10][8];
    ele[6][11] != ele[10][9];
    ele[6][11] != ele[11][10];
    ele[6][11] != ele[11][11];
    ele[6][11] != ele[11][6];
    ele[6][11] != ele[11][7];
    ele[6][11] != ele[11][8];
    ele[6][11] != ele[11][9];
    ele[6][11] != ele[12][11];
    ele[6][11] != ele[13][11];
    ele[6][11] != ele[14][11];
    ele[6][11] != ele[15][11];
    ele[6][11] != ele[16][11];
    ele[6][11] != ele[17][11];
    ele[6][11] != ele[18][11];
    ele[6][11] != ele[19][11];
    ele[6][11] != ele[20][11];
    ele[6][11] != ele[21][11];
    ele[6][11] != ele[22][11];
    ele[6][11] != ele[23][11];
    ele[6][11] != ele[24][11];
    ele[6][11] != ele[25][11];
    ele[6][11] != ele[26][11];
    ele[6][11] != ele[27][11];
    ele[6][11] != ele[28][11];
    ele[6][11] != ele[29][11];
    ele[6][11] != ele[30][11];
    ele[6][11] != ele[31][11];
    ele[6][11] != ele[32][11];
    ele[6][11] != ele[33][11];
    ele[6][11] != ele[34][11];
    ele[6][11] != ele[35][11];
    ele[6][11] != ele[6][12];
    ele[6][11] != ele[6][13];
    ele[6][11] != ele[6][14];
    ele[6][11] != ele[6][15];
    ele[6][11] != ele[6][16];
    ele[6][11] != ele[6][17];
    ele[6][11] != ele[6][18];
    ele[6][11] != ele[6][19];
    ele[6][11] != ele[6][20];
    ele[6][11] != ele[6][21];
    ele[6][11] != ele[6][22];
    ele[6][11] != ele[6][23];
    ele[6][11] != ele[6][24];
    ele[6][11] != ele[6][25];
    ele[6][11] != ele[6][26];
    ele[6][11] != ele[6][27];
    ele[6][11] != ele[6][28];
    ele[6][11] != ele[6][29];
    ele[6][11] != ele[6][30];
    ele[6][11] != ele[6][31];
    ele[6][11] != ele[6][32];
    ele[6][11] != ele[6][33];
    ele[6][11] != ele[6][34];
    ele[6][11] != ele[6][35];
    ele[6][11] != ele[7][10];
    ele[6][11] != ele[7][11];
    ele[6][11] != ele[7][6];
    ele[6][11] != ele[7][7];
    ele[6][11] != ele[7][8];
    ele[6][11] != ele[7][9];
    ele[6][11] != ele[8][10];
    ele[6][11] != ele[8][11];
    ele[6][11] != ele[8][6];
    ele[6][11] != ele[8][7];
    ele[6][11] != ele[8][8];
    ele[6][11] != ele[8][9];
    ele[6][11] != ele[9][10];
    ele[6][11] != ele[9][11];
    ele[6][11] != ele[9][6];
    ele[6][11] != ele[9][7];
    ele[6][11] != ele[9][8];
    ele[6][11] != ele[9][9];
    ele[6][12] != ele[10][12];
    ele[6][12] != ele[10][13];
    ele[6][12] != ele[10][14];
    ele[6][12] != ele[10][15];
    ele[6][12] != ele[10][16];
    ele[6][12] != ele[10][17];
    ele[6][12] != ele[11][12];
    ele[6][12] != ele[11][13];
    ele[6][12] != ele[11][14];
    ele[6][12] != ele[11][15];
    ele[6][12] != ele[11][16];
    ele[6][12] != ele[11][17];
    ele[6][12] != ele[12][12];
    ele[6][12] != ele[13][12];
    ele[6][12] != ele[14][12];
    ele[6][12] != ele[15][12];
    ele[6][12] != ele[16][12];
    ele[6][12] != ele[17][12];
    ele[6][12] != ele[18][12];
    ele[6][12] != ele[19][12];
    ele[6][12] != ele[20][12];
    ele[6][12] != ele[21][12];
    ele[6][12] != ele[22][12];
    ele[6][12] != ele[23][12];
    ele[6][12] != ele[24][12];
    ele[6][12] != ele[25][12];
    ele[6][12] != ele[26][12];
    ele[6][12] != ele[27][12];
    ele[6][12] != ele[28][12];
    ele[6][12] != ele[29][12];
    ele[6][12] != ele[30][12];
    ele[6][12] != ele[31][12];
    ele[6][12] != ele[32][12];
    ele[6][12] != ele[33][12];
    ele[6][12] != ele[34][12];
    ele[6][12] != ele[35][12];
    ele[6][12] != ele[6][13];
    ele[6][12] != ele[6][14];
    ele[6][12] != ele[6][15];
    ele[6][12] != ele[6][16];
    ele[6][12] != ele[6][17];
    ele[6][12] != ele[6][18];
    ele[6][12] != ele[6][19];
    ele[6][12] != ele[6][20];
    ele[6][12] != ele[6][21];
    ele[6][12] != ele[6][22];
    ele[6][12] != ele[6][23];
    ele[6][12] != ele[6][24];
    ele[6][12] != ele[6][25];
    ele[6][12] != ele[6][26];
    ele[6][12] != ele[6][27];
    ele[6][12] != ele[6][28];
    ele[6][12] != ele[6][29];
    ele[6][12] != ele[6][30];
    ele[6][12] != ele[6][31];
    ele[6][12] != ele[6][32];
    ele[6][12] != ele[6][33];
    ele[6][12] != ele[6][34];
    ele[6][12] != ele[6][35];
    ele[6][12] != ele[7][12];
    ele[6][12] != ele[7][13];
    ele[6][12] != ele[7][14];
    ele[6][12] != ele[7][15];
    ele[6][12] != ele[7][16];
    ele[6][12] != ele[7][17];
    ele[6][12] != ele[8][12];
    ele[6][12] != ele[8][13];
    ele[6][12] != ele[8][14];
    ele[6][12] != ele[8][15];
    ele[6][12] != ele[8][16];
    ele[6][12] != ele[8][17];
    ele[6][12] != ele[9][12];
    ele[6][12] != ele[9][13];
    ele[6][12] != ele[9][14];
    ele[6][12] != ele[9][15];
    ele[6][12] != ele[9][16];
    ele[6][12] != ele[9][17];
    ele[6][13] != ele[10][12];
    ele[6][13] != ele[10][13];
    ele[6][13] != ele[10][14];
    ele[6][13] != ele[10][15];
    ele[6][13] != ele[10][16];
    ele[6][13] != ele[10][17];
    ele[6][13] != ele[11][12];
    ele[6][13] != ele[11][13];
    ele[6][13] != ele[11][14];
    ele[6][13] != ele[11][15];
    ele[6][13] != ele[11][16];
    ele[6][13] != ele[11][17];
    ele[6][13] != ele[12][13];
    ele[6][13] != ele[13][13];
    ele[6][13] != ele[14][13];
    ele[6][13] != ele[15][13];
    ele[6][13] != ele[16][13];
    ele[6][13] != ele[17][13];
    ele[6][13] != ele[18][13];
    ele[6][13] != ele[19][13];
    ele[6][13] != ele[20][13];
    ele[6][13] != ele[21][13];
    ele[6][13] != ele[22][13];
    ele[6][13] != ele[23][13];
    ele[6][13] != ele[24][13];
    ele[6][13] != ele[25][13];
    ele[6][13] != ele[26][13];
    ele[6][13] != ele[27][13];
    ele[6][13] != ele[28][13];
    ele[6][13] != ele[29][13];
    ele[6][13] != ele[30][13];
    ele[6][13] != ele[31][13];
    ele[6][13] != ele[32][13];
    ele[6][13] != ele[33][13];
    ele[6][13] != ele[34][13];
    ele[6][13] != ele[35][13];
    ele[6][13] != ele[6][14];
    ele[6][13] != ele[6][15];
    ele[6][13] != ele[6][16];
    ele[6][13] != ele[6][17];
    ele[6][13] != ele[6][18];
    ele[6][13] != ele[6][19];
    ele[6][13] != ele[6][20];
    ele[6][13] != ele[6][21];
    ele[6][13] != ele[6][22];
    ele[6][13] != ele[6][23];
    ele[6][13] != ele[6][24];
    ele[6][13] != ele[6][25];
    ele[6][13] != ele[6][26];
    ele[6][13] != ele[6][27];
    ele[6][13] != ele[6][28];
    ele[6][13] != ele[6][29];
    ele[6][13] != ele[6][30];
    ele[6][13] != ele[6][31];
    ele[6][13] != ele[6][32];
    ele[6][13] != ele[6][33];
    ele[6][13] != ele[6][34];
    ele[6][13] != ele[6][35];
    ele[6][13] != ele[7][12];
    ele[6][13] != ele[7][13];
    ele[6][13] != ele[7][14];
    ele[6][13] != ele[7][15];
    ele[6][13] != ele[7][16];
    ele[6][13] != ele[7][17];
    ele[6][13] != ele[8][12];
    ele[6][13] != ele[8][13];
    ele[6][13] != ele[8][14];
    ele[6][13] != ele[8][15];
    ele[6][13] != ele[8][16];
    ele[6][13] != ele[8][17];
    ele[6][13] != ele[9][12];
    ele[6][13] != ele[9][13];
    ele[6][13] != ele[9][14];
    ele[6][13] != ele[9][15];
    ele[6][13] != ele[9][16];
    ele[6][13] != ele[9][17];
    ele[6][14] != ele[10][12];
    ele[6][14] != ele[10][13];
    ele[6][14] != ele[10][14];
    ele[6][14] != ele[10][15];
    ele[6][14] != ele[10][16];
    ele[6][14] != ele[10][17];
    ele[6][14] != ele[11][12];
    ele[6][14] != ele[11][13];
    ele[6][14] != ele[11][14];
    ele[6][14] != ele[11][15];
    ele[6][14] != ele[11][16];
    ele[6][14] != ele[11][17];
    ele[6][14] != ele[12][14];
    ele[6][14] != ele[13][14];
    ele[6][14] != ele[14][14];
    ele[6][14] != ele[15][14];
    ele[6][14] != ele[16][14];
    ele[6][14] != ele[17][14];
    ele[6][14] != ele[18][14];
    ele[6][14] != ele[19][14];
    ele[6][14] != ele[20][14];
    ele[6][14] != ele[21][14];
    ele[6][14] != ele[22][14];
    ele[6][14] != ele[23][14];
    ele[6][14] != ele[24][14];
    ele[6][14] != ele[25][14];
    ele[6][14] != ele[26][14];
    ele[6][14] != ele[27][14];
    ele[6][14] != ele[28][14];
    ele[6][14] != ele[29][14];
    ele[6][14] != ele[30][14];
    ele[6][14] != ele[31][14];
    ele[6][14] != ele[32][14];
    ele[6][14] != ele[33][14];
    ele[6][14] != ele[34][14];
    ele[6][14] != ele[35][14];
    ele[6][14] != ele[6][15];
    ele[6][14] != ele[6][16];
    ele[6][14] != ele[6][17];
    ele[6][14] != ele[6][18];
    ele[6][14] != ele[6][19];
    ele[6][14] != ele[6][20];
    ele[6][14] != ele[6][21];
    ele[6][14] != ele[6][22];
    ele[6][14] != ele[6][23];
    ele[6][14] != ele[6][24];
    ele[6][14] != ele[6][25];
    ele[6][14] != ele[6][26];
    ele[6][14] != ele[6][27];
    ele[6][14] != ele[6][28];
    ele[6][14] != ele[6][29];
    ele[6][14] != ele[6][30];
    ele[6][14] != ele[6][31];
    ele[6][14] != ele[6][32];
    ele[6][14] != ele[6][33];
    ele[6][14] != ele[6][34];
    ele[6][14] != ele[6][35];
    ele[6][14] != ele[7][12];
    ele[6][14] != ele[7][13];
    ele[6][14] != ele[7][14];
    ele[6][14] != ele[7][15];
    ele[6][14] != ele[7][16];
    ele[6][14] != ele[7][17];
    ele[6][14] != ele[8][12];
    ele[6][14] != ele[8][13];
    ele[6][14] != ele[8][14];
    ele[6][14] != ele[8][15];
    ele[6][14] != ele[8][16];
    ele[6][14] != ele[8][17];
    ele[6][14] != ele[9][12];
    ele[6][14] != ele[9][13];
    ele[6][14] != ele[9][14];
    ele[6][14] != ele[9][15];
    ele[6][14] != ele[9][16];
    ele[6][14] != ele[9][17];
    ele[6][15] != ele[10][12];
    ele[6][15] != ele[10][13];
    ele[6][15] != ele[10][14];
    ele[6][15] != ele[10][15];
    ele[6][15] != ele[10][16];
    ele[6][15] != ele[10][17];
    ele[6][15] != ele[11][12];
    ele[6][15] != ele[11][13];
    ele[6][15] != ele[11][14];
    ele[6][15] != ele[11][15];
    ele[6][15] != ele[11][16];
    ele[6][15] != ele[11][17];
    ele[6][15] != ele[12][15];
    ele[6][15] != ele[13][15];
    ele[6][15] != ele[14][15];
    ele[6][15] != ele[15][15];
    ele[6][15] != ele[16][15];
    ele[6][15] != ele[17][15];
    ele[6][15] != ele[18][15];
    ele[6][15] != ele[19][15];
    ele[6][15] != ele[20][15];
    ele[6][15] != ele[21][15];
    ele[6][15] != ele[22][15];
    ele[6][15] != ele[23][15];
    ele[6][15] != ele[24][15];
    ele[6][15] != ele[25][15];
    ele[6][15] != ele[26][15];
    ele[6][15] != ele[27][15];
    ele[6][15] != ele[28][15];
    ele[6][15] != ele[29][15];
    ele[6][15] != ele[30][15];
    ele[6][15] != ele[31][15];
    ele[6][15] != ele[32][15];
    ele[6][15] != ele[33][15];
    ele[6][15] != ele[34][15];
    ele[6][15] != ele[35][15];
    ele[6][15] != ele[6][16];
    ele[6][15] != ele[6][17];
    ele[6][15] != ele[6][18];
    ele[6][15] != ele[6][19];
    ele[6][15] != ele[6][20];
    ele[6][15] != ele[6][21];
    ele[6][15] != ele[6][22];
    ele[6][15] != ele[6][23];
    ele[6][15] != ele[6][24];
    ele[6][15] != ele[6][25];
    ele[6][15] != ele[6][26];
    ele[6][15] != ele[6][27];
    ele[6][15] != ele[6][28];
    ele[6][15] != ele[6][29];
    ele[6][15] != ele[6][30];
    ele[6][15] != ele[6][31];
    ele[6][15] != ele[6][32];
    ele[6][15] != ele[6][33];
    ele[6][15] != ele[6][34];
    ele[6][15] != ele[6][35];
    ele[6][15] != ele[7][12];
    ele[6][15] != ele[7][13];
    ele[6][15] != ele[7][14];
    ele[6][15] != ele[7][15];
    ele[6][15] != ele[7][16];
    ele[6][15] != ele[7][17];
    ele[6][15] != ele[8][12];
    ele[6][15] != ele[8][13];
    ele[6][15] != ele[8][14];
    ele[6][15] != ele[8][15];
    ele[6][15] != ele[8][16];
    ele[6][15] != ele[8][17];
    ele[6][15] != ele[9][12];
    ele[6][15] != ele[9][13];
    ele[6][15] != ele[9][14];
    ele[6][15] != ele[9][15];
    ele[6][15] != ele[9][16];
    ele[6][15] != ele[9][17];
    ele[6][16] != ele[10][12];
    ele[6][16] != ele[10][13];
    ele[6][16] != ele[10][14];
    ele[6][16] != ele[10][15];
    ele[6][16] != ele[10][16];
    ele[6][16] != ele[10][17];
    ele[6][16] != ele[11][12];
    ele[6][16] != ele[11][13];
    ele[6][16] != ele[11][14];
    ele[6][16] != ele[11][15];
    ele[6][16] != ele[11][16];
    ele[6][16] != ele[11][17];
    ele[6][16] != ele[12][16];
    ele[6][16] != ele[13][16];
    ele[6][16] != ele[14][16];
    ele[6][16] != ele[15][16];
    ele[6][16] != ele[16][16];
    ele[6][16] != ele[17][16];
    ele[6][16] != ele[18][16];
    ele[6][16] != ele[19][16];
    ele[6][16] != ele[20][16];
    ele[6][16] != ele[21][16];
    ele[6][16] != ele[22][16];
    ele[6][16] != ele[23][16];
    ele[6][16] != ele[24][16];
    ele[6][16] != ele[25][16];
    ele[6][16] != ele[26][16];
    ele[6][16] != ele[27][16];
    ele[6][16] != ele[28][16];
    ele[6][16] != ele[29][16];
    ele[6][16] != ele[30][16];
    ele[6][16] != ele[31][16];
    ele[6][16] != ele[32][16];
    ele[6][16] != ele[33][16];
    ele[6][16] != ele[34][16];
    ele[6][16] != ele[35][16];
    ele[6][16] != ele[6][17];
    ele[6][16] != ele[6][18];
    ele[6][16] != ele[6][19];
    ele[6][16] != ele[6][20];
    ele[6][16] != ele[6][21];
    ele[6][16] != ele[6][22];
    ele[6][16] != ele[6][23];
    ele[6][16] != ele[6][24];
    ele[6][16] != ele[6][25];
    ele[6][16] != ele[6][26];
    ele[6][16] != ele[6][27];
    ele[6][16] != ele[6][28];
    ele[6][16] != ele[6][29];
    ele[6][16] != ele[6][30];
    ele[6][16] != ele[6][31];
    ele[6][16] != ele[6][32];
    ele[6][16] != ele[6][33];
    ele[6][16] != ele[6][34];
    ele[6][16] != ele[6][35];
    ele[6][16] != ele[7][12];
    ele[6][16] != ele[7][13];
    ele[6][16] != ele[7][14];
    ele[6][16] != ele[7][15];
    ele[6][16] != ele[7][16];
    ele[6][16] != ele[7][17];
    ele[6][16] != ele[8][12];
    ele[6][16] != ele[8][13];
    ele[6][16] != ele[8][14];
    ele[6][16] != ele[8][15];
    ele[6][16] != ele[8][16];
    ele[6][16] != ele[8][17];
    ele[6][16] != ele[9][12];
    ele[6][16] != ele[9][13];
    ele[6][16] != ele[9][14];
    ele[6][16] != ele[9][15];
    ele[6][16] != ele[9][16];
    ele[6][16] != ele[9][17];
    ele[6][17] != ele[10][12];
    ele[6][17] != ele[10][13];
    ele[6][17] != ele[10][14];
    ele[6][17] != ele[10][15];
    ele[6][17] != ele[10][16];
    ele[6][17] != ele[10][17];
    ele[6][17] != ele[11][12];
    ele[6][17] != ele[11][13];
    ele[6][17] != ele[11][14];
    ele[6][17] != ele[11][15];
    ele[6][17] != ele[11][16];
    ele[6][17] != ele[11][17];
    ele[6][17] != ele[12][17];
    ele[6][17] != ele[13][17];
    ele[6][17] != ele[14][17];
    ele[6][17] != ele[15][17];
    ele[6][17] != ele[16][17];
    ele[6][17] != ele[17][17];
    ele[6][17] != ele[18][17];
    ele[6][17] != ele[19][17];
    ele[6][17] != ele[20][17];
    ele[6][17] != ele[21][17];
    ele[6][17] != ele[22][17];
    ele[6][17] != ele[23][17];
    ele[6][17] != ele[24][17];
    ele[6][17] != ele[25][17];
    ele[6][17] != ele[26][17];
    ele[6][17] != ele[27][17];
    ele[6][17] != ele[28][17];
    ele[6][17] != ele[29][17];
    ele[6][17] != ele[30][17];
    ele[6][17] != ele[31][17];
    ele[6][17] != ele[32][17];
    ele[6][17] != ele[33][17];
    ele[6][17] != ele[34][17];
    ele[6][17] != ele[35][17];
    ele[6][17] != ele[6][18];
    ele[6][17] != ele[6][19];
    ele[6][17] != ele[6][20];
    ele[6][17] != ele[6][21];
    ele[6][17] != ele[6][22];
    ele[6][17] != ele[6][23];
    ele[6][17] != ele[6][24];
    ele[6][17] != ele[6][25];
    ele[6][17] != ele[6][26];
    ele[6][17] != ele[6][27];
    ele[6][17] != ele[6][28];
    ele[6][17] != ele[6][29];
    ele[6][17] != ele[6][30];
    ele[6][17] != ele[6][31];
    ele[6][17] != ele[6][32];
    ele[6][17] != ele[6][33];
    ele[6][17] != ele[6][34];
    ele[6][17] != ele[6][35];
    ele[6][17] != ele[7][12];
    ele[6][17] != ele[7][13];
    ele[6][17] != ele[7][14];
    ele[6][17] != ele[7][15];
    ele[6][17] != ele[7][16];
    ele[6][17] != ele[7][17];
    ele[6][17] != ele[8][12];
    ele[6][17] != ele[8][13];
    ele[6][17] != ele[8][14];
    ele[6][17] != ele[8][15];
    ele[6][17] != ele[8][16];
    ele[6][17] != ele[8][17];
    ele[6][17] != ele[9][12];
    ele[6][17] != ele[9][13];
    ele[6][17] != ele[9][14];
    ele[6][17] != ele[9][15];
    ele[6][17] != ele[9][16];
    ele[6][17] != ele[9][17];
    ele[6][18] != ele[10][18];
    ele[6][18] != ele[10][19];
    ele[6][18] != ele[10][20];
    ele[6][18] != ele[10][21];
    ele[6][18] != ele[10][22];
    ele[6][18] != ele[10][23];
    ele[6][18] != ele[11][18];
    ele[6][18] != ele[11][19];
    ele[6][18] != ele[11][20];
    ele[6][18] != ele[11][21];
    ele[6][18] != ele[11][22];
    ele[6][18] != ele[11][23];
    ele[6][18] != ele[12][18];
    ele[6][18] != ele[13][18];
    ele[6][18] != ele[14][18];
    ele[6][18] != ele[15][18];
    ele[6][18] != ele[16][18];
    ele[6][18] != ele[17][18];
    ele[6][18] != ele[18][18];
    ele[6][18] != ele[19][18];
    ele[6][18] != ele[20][18];
    ele[6][18] != ele[21][18];
    ele[6][18] != ele[22][18];
    ele[6][18] != ele[23][18];
    ele[6][18] != ele[24][18];
    ele[6][18] != ele[25][18];
    ele[6][18] != ele[26][18];
    ele[6][18] != ele[27][18];
    ele[6][18] != ele[28][18];
    ele[6][18] != ele[29][18];
    ele[6][18] != ele[30][18];
    ele[6][18] != ele[31][18];
    ele[6][18] != ele[32][18];
    ele[6][18] != ele[33][18];
    ele[6][18] != ele[34][18];
    ele[6][18] != ele[35][18];
    ele[6][18] != ele[6][19];
    ele[6][18] != ele[6][20];
    ele[6][18] != ele[6][21];
    ele[6][18] != ele[6][22];
    ele[6][18] != ele[6][23];
    ele[6][18] != ele[6][24];
    ele[6][18] != ele[6][25];
    ele[6][18] != ele[6][26];
    ele[6][18] != ele[6][27];
    ele[6][18] != ele[6][28];
    ele[6][18] != ele[6][29];
    ele[6][18] != ele[6][30];
    ele[6][18] != ele[6][31];
    ele[6][18] != ele[6][32];
    ele[6][18] != ele[6][33];
    ele[6][18] != ele[6][34];
    ele[6][18] != ele[6][35];
    ele[6][18] != ele[7][18];
    ele[6][18] != ele[7][19];
    ele[6][18] != ele[7][20];
    ele[6][18] != ele[7][21];
    ele[6][18] != ele[7][22];
    ele[6][18] != ele[7][23];
    ele[6][18] != ele[8][18];
    ele[6][18] != ele[8][19];
    ele[6][18] != ele[8][20];
    ele[6][18] != ele[8][21];
    ele[6][18] != ele[8][22];
    ele[6][18] != ele[8][23];
    ele[6][18] != ele[9][18];
    ele[6][18] != ele[9][19];
    ele[6][18] != ele[9][20];
    ele[6][18] != ele[9][21];
    ele[6][18] != ele[9][22];
    ele[6][18] != ele[9][23];
    ele[6][19] != ele[10][18];
    ele[6][19] != ele[10][19];
    ele[6][19] != ele[10][20];
    ele[6][19] != ele[10][21];
    ele[6][19] != ele[10][22];
    ele[6][19] != ele[10][23];
    ele[6][19] != ele[11][18];
    ele[6][19] != ele[11][19];
    ele[6][19] != ele[11][20];
    ele[6][19] != ele[11][21];
    ele[6][19] != ele[11][22];
    ele[6][19] != ele[11][23];
    ele[6][19] != ele[12][19];
    ele[6][19] != ele[13][19];
    ele[6][19] != ele[14][19];
    ele[6][19] != ele[15][19];
    ele[6][19] != ele[16][19];
    ele[6][19] != ele[17][19];
    ele[6][19] != ele[18][19];
    ele[6][19] != ele[19][19];
    ele[6][19] != ele[20][19];
    ele[6][19] != ele[21][19];
    ele[6][19] != ele[22][19];
    ele[6][19] != ele[23][19];
    ele[6][19] != ele[24][19];
    ele[6][19] != ele[25][19];
    ele[6][19] != ele[26][19];
    ele[6][19] != ele[27][19];
    ele[6][19] != ele[28][19];
    ele[6][19] != ele[29][19];
    ele[6][19] != ele[30][19];
    ele[6][19] != ele[31][19];
    ele[6][19] != ele[32][19];
    ele[6][19] != ele[33][19];
    ele[6][19] != ele[34][19];
    ele[6][19] != ele[35][19];
    ele[6][19] != ele[6][20];
    ele[6][19] != ele[6][21];
    ele[6][19] != ele[6][22];
    ele[6][19] != ele[6][23];
    ele[6][19] != ele[6][24];
    ele[6][19] != ele[6][25];
    ele[6][19] != ele[6][26];
    ele[6][19] != ele[6][27];
    ele[6][19] != ele[6][28];
    ele[6][19] != ele[6][29];
    ele[6][19] != ele[6][30];
    ele[6][19] != ele[6][31];
    ele[6][19] != ele[6][32];
    ele[6][19] != ele[6][33];
    ele[6][19] != ele[6][34];
    ele[6][19] != ele[6][35];
    ele[6][19] != ele[7][18];
    ele[6][19] != ele[7][19];
    ele[6][19] != ele[7][20];
    ele[6][19] != ele[7][21];
    ele[6][19] != ele[7][22];
    ele[6][19] != ele[7][23];
    ele[6][19] != ele[8][18];
    ele[6][19] != ele[8][19];
    ele[6][19] != ele[8][20];
    ele[6][19] != ele[8][21];
    ele[6][19] != ele[8][22];
    ele[6][19] != ele[8][23];
    ele[6][19] != ele[9][18];
    ele[6][19] != ele[9][19];
    ele[6][19] != ele[9][20];
    ele[6][19] != ele[9][21];
    ele[6][19] != ele[9][22];
    ele[6][19] != ele[9][23];
    ele[6][2] != ele[10][0];
    ele[6][2] != ele[10][1];
    ele[6][2] != ele[10][2];
    ele[6][2] != ele[10][3];
    ele[6][2] != ele[10][4];
    ele[6][2] != ele[10][5];
    ele[6][2] != ele[11][0];
    ele[6][2] != ele[11][1];
    ele[6][2] != ele[11][2];
    ele[6][2] != ele[11][3];
    ele[6][2] != ele[11][4];
    ele[6][2] != ele[11][5];
    ele[6][2] != ele[12][2];
    ele[6][2] != ele[13][2];
    ele[6][2] != ele[14][2];
    ele[6][2] != ele[15][2];
    ele[6][2] != ele[16][2];
    ele[6][2] != ele[17][2];
    ele[6][2] != ele[18][2];
    ele[6][2] != ele[19][2];
    ele[6][2] != ele[20][2];
    ele[6][2] != ele[21][2];
    ele[6][2] != ele[22][2];
    ele[6][2] != ele[23][2];
    ele[6][2] != ele[24][2];
    ele[6][2] != ele[25][2];
    ele[6][2] != ele[26][2];
    ele[6][2] != ele[27][2];
    ele[6][2] != ele[28][2];
    ele[6][2] != ele[29][2];
    ele[6][2] != ele[30][2];
    ele[6][2] != ele[31][2];
    ele[6][2] != ele[32][2];
    ele[6][2] != ele[33][2];
    ele[6][2] != ele[34][2];
    ele[6][2] != ele[35][2];
    ele[6][2] != ele[6][10];
    ele[6][2] != ele[6][11];
    ele[6][2] != ele[6][12];
    ele[6][2] != ele[6][13];
    ele[6][2] != ele[6][14];
    ele[6][2] != ele[6][15];
    ele[6][2] != ele[6][16];
    ele[6][2] != ele[6][17];
    ele[6][2] != ele[6][18];
    ele[6][2] != ele[6][19];
    ele[6][2] != ele[6][20];
    ele[6][2] != ele[6][21];
    ele[6][2] != ele[6][22];
    ele[6][2] != ele[6][23];
    ele[6][2] != ele[6][24];
    ele[6][2] != ele[6][25];
    ele[6][2] != ele[6][26];
    ele[6][2] != ele[6][27];
    ele[6][2] != ele[6][28];
    ele[6][2] != ele[6][29];
    ele[6][2] != ele[6][3];
    ele[6][2] != ele[6][30];
    ele[6][2] != ele[6][31];
    ele[6][2] != ele[6][32];
    ele[6][2] != ele[6][33];
    ele[6][2] != ele[6][34];
    ele[6][2] != ele[6][35];
    ele[6][2] != ele[6][4];
    ele[6][2] != ele[6][5];
    ele[6][2] != ele[6][6];
    ele[6][2] != ele[6][7];
    ele[6][2] != ele[6][8];
    ele[6][2] != ele[6][9];
    ele[6][2] != ele[7][0];
    ele[6][2] != ele[7][1];
    ele[6][2] != ele[7][2];
    ele[6][2] != ele[7][3];
    ele[6][2] != ele[7][4];
    ele[6][2] != ele[7][5];
    ele[6][2] != ele[8][0];
    ele[6][2] != ele[8][1];
    ele[6][2] != ele[8][2];
    ele[6][2] != ele[8][3];
    ele[6][2] != ele[8][4];
    ele[6][2] != ele[8][5];
    ele[6][2] != ele[9][0];
    ele[6][2] != ele[9][1];
    ele[6][2] != ele[9][2];
    ele[6][2] != ele[9][3];
    ele[6][2] != ele[9][4];
    ele[6][2] != ele[9][5];
    ele[6][20] != ele[10][18];
    ele[6][20] != ele[10][19];
    ele[6][20] != ele[10][20];
    ele[6][20] != ele[10][21];
    ele[6][20] != ele[10][22];
    ele[6][20] != ele[10][23];
    ele[6][20] != ele[11][18];
    ele[6][20] != ele[11][19];
    ele[6][20] != ele[11][20];
    ele[6][20] != ele[11][21];
    ele[6][20] != ele[11][22];
    ele[6][20] != ele[11][23];
    ele[6][20] != ele[12][20];
    ele[6][20] != ele[13][20];
    ele[6][20] != ele[14][20];
    ele[6][20] != ele[15][20];
    ele[6][20] != ele[16][20];
    ele[6][20] != ele[17][20];
    ele[6][20] != ele[18][20];
    ele[6][20] != ele[19][20];
    ele[6][20] != ele[20][20];
    ele[6][20] != ele[21][20];
    ele[6][20] != ele[22][20];
    ele[6][20] != ele[23][20];
    ele[6][20] != ele[24][20];
    ele[6][20] != ele[25][20];
    ele[6][20] != ele[26][20];
    ele[6][20] != ele[27][20];
    ele[6][20] != ele[28][20];
    ele[6][20] != ele[29][20];
    ele[6][20] != ele[30][20];
    ele[6][20] != ele[31][20];
    ele[6][20] != ele[32][20];
    ele[6][20] != ele[33][20];
    ele[6][20] != ele[34][20];
    ele[6][20] != ele[35][20];
    ele[6][20] != ele[6][21];
    ele[6][20] != ele[6][22];
    ele[6][20] != ele[6][23];
    ele[6][20] != ele[6][24];
    ele[6][20] != ele[6][25];
    ele[6][20] != ele[6][26];
    ele[6][20] != ele[6][27];
    ele[6][20] != ele[6][28];
    ele[6][20] != ele[6][29];
    ele[6][20] != ele[6][30];
    ele[6][20] != ele[6][31];
    ele[6][20] != ele[6][32];
    ele[6][20] != ele[6][33];
    ele[6][20] != ele[6][34];
    ele[6][20] != ele[6][35];
    ele[6][20] != ele[7][18];
    ele[6][20] != ele[7][19];
    ele[6][20] != ele[7][20];
    ele[6][20] != ele[7][21];
    ele[6][20] != ele[7][22];
    ele[6][20] != ele[7][23];
    ele[6][20] != ele[8][18];
    ele[6][20] != ele[8][19];
    ele[6][20] != ele[8][20];
    ele[6][20] != ele[8][21];
    ele[6][20] != ele[8][22];
    ele[6][20] != ele[8][23];
    ele[6][20] != ele[9][18];
    ele[6][20] != ele[9][19];
    ele[6][20] != ele[9][20];
    ele[6][20] != ele[9][21];
    ele[6][20] != ele[9][22];
    ele[6][20] != ele[9][23];
    ele[6][21] != ele[10][18];
    ele[6][21] != ele[10][19];
    ele[6][21] != ele[10][20];
    ele[6][21] != ele[10][21];
    ele[6][21] != ele[10][22];
    ele[6][21] != ele[10][23];
    ele[6][21] != ele[11][18];
    ele[6][21] != ele[11][19];
    ele[6][21] != ele[11][20];
    ele[6][21] != ele[11][21];
    ele[6][21] != ele[11][22];
    ele[6][21] != ele[11][23];
    ele[6][21] != ele[12][21];
    ele[6][21] != ele[13][21];
    ele[6][21] != ele[14][21];
    ele[6][21] != ele[15][21];
    ele[6][21] != ele[16][21];
    ele[6][21] != ele[17][21];
    ele[6][21] != ele[18][21];
    ele[6][21] != ele[19][21];
    ele[6][21] != ele[20][21];
    ele[6][21] != ele[21][21];
    ele[6][21] != ele[22][21];
    ele[6][21] != ele[23][21];
    ele[6][21] != ele[24][21];
    ele[6][21] != ele[25][21];
    ele[6][21] != ele[26][21];
    ele[6][21] != ele[27][21];
    ele[6][21] != ele[28][21];
    ele[6][21] != ele[29][21];
    ele[6][21] != ele[30][21];
    ele[6][21] != ele[31][21];
    ele[6][21] != ele[32][21];
    ele[6][21] != ele[33][21];
    ele[6][21] != ele[34][21];
    ele[6][21] != ele[35][21];
    ele[6][21] != ele[6][22];
    ele[6][21] != ele[6][23];
    ele[6][21] != ele[6][24];
    ele[6][21] != ele[6][25];
    ele[6][21] != ele[6][26];
    ele[6][21] != ele[6][27];
    ele[6][21] != ele[6][28];
    ele[6][21] != ele[6][29];
    ele[6][21] != ele[6][30];
    ele[6][21] != ele[6][31];
    ele[6][21] != ele[6][32];
    ele[6][21] != ele[6][33];
    ele[6][21] != ele[6][34];
    ele[6][21] != ele[6][35];
    ele[6][21] != ele[7][18];
    ele[6][21] != ele[7][19];
    ele[6][21] != ele[7][20];
    ele[6][21] != ele[7][21];
    ele[6][21] != ele[7][22];
    ele[6][21] != ele[7][23];
    ele[6][21] != ele[8][18];
    ele[6][21] != ele[8][19];
    ele[6][21] != ele[8][20];
    ele[6][21] != ele[8][21];
    ele[6][21] != ele[8][22];
    ele[6][21] != ele[8][23];
    ele[6][21] != ele[9][18];
    ele[6][21] != ele[9][19];
    ele[6][21] != ele[9][20];
    ele[6][21] != ele[9][21];
    ele[6][21] != ele[9][22];
    ele[6][21] != ele[9][23];
    ele[6][22] != ele[10][18];
    ele[6][22] != ele[10][19];
    ele[6][22] != ele[10][20];
    ele[6][22] != ele[10][21];
    ele[6][22] != ele[10][22];
    ele[6][22] != ele[10][23];
    ele[6][22] != ele[11][18];
    ele[6][22] != ele[11][19];
    ele[6][22] != ele[11][20];
    ele[6][22] != ele[11][21];
    ele[6][22] != ele[11][22];
    ele[6][22] != ele[11][23];
    ele[6][22] != ele[12][22];
    ele[6][22] != ele[13][22];
    ele[6][22] != ele[14][22];
    ele[6][22] != ele[15][22];
    ele[6][22] != ele[16][22];
    ele[6][22] != ele[17][22];
    ele[6][22] != ele[18][22];
    ele[6][22] != ele[19][22];
    ele[6][22] != ele[20][22];
    ele[6][22] != ele[21][22];
    ele[6][22] != ele[22][22];
    ele[6][22] != ele[23][22];
    ele[6][22] != ele[24][22];
    ele[6][22] != ele[25][22];
    ele[6][22] != ele[26][22];
    ele[6][22] != ele[27][22];
    ele[6][22] != ele[28][22];
    ele[6][22] != ele[29][22];
    ele[6][22] != ele[30][22];
    ele[6][22] != ele[31][22];
    ele[6][22] != ele[32][22];
    ele[6][22] != ele[33][22];
    ele[6][22] != ele[34][22];
    ele[6][22] != ele[35][22];
    ele[6][22] != ele[6][23];
    ele[6][22] != ele[6][24];
    ele[6][22] != ele[6][25];
    ele[6][22] != ele[6][26];
    ele[6][22] != ele[6][27];
    ele[6][22] != ele[6][28];
    ele[6][22] != ele[6][29];
    ele[6][22] != ele[6][30];
    ele[6][22] != ele[6][31];
    ele[6][22] != ele[6][32];
    ele[6][22] != ele[6][33];
    ele[6][22] != ele[6][34];
    ele[6][22] != ele[6][35];
    ele[6][22] != ele[7][18];
    ele[6][22] != ele[7][19];
    ele[6][22] != ele[7][20];
    ele[6][22] != ele[7][21];
    ele[6][22] != ele[7][22];
    ele[6][22] != ele[7][23];
    ele[6][22] != ele[8][18];
    ele[6][22] != ele[8][19];
    ele[6][22] != ele[8][20];
    ele[6][22] != ele[8][21];
    ele[6][22] != ele[8][22];
    ele[6][22] != ele[8][23];
    ele[6][22] != ele[9][18];
    ele[6][22] != ele[9][19];
    ele[6][22] != ele[9][20];
    ele[6][22] != ele[9][21];
    ele[6][22] != ele[9][22];
    ele[6][22] != ele[9][23];
    ele[6][23] != ele[10][18];
    ele[6][23] != ele[10][19];
    ele[6][23] != ele[10][20];
    ele[6][23] != ele[10][21];
    ele[6][23] != ele[10][22];
    ele[6][23] != ele[10][23];
    ele[6][23] != ele[11][18];
    ele[6][23] != ele[11][19];
    ele[6][23] != ele[11][20];
    ele[6][23] != ele[11][21];
    ele[6][23] != ele[11][22];
    ele[6][23] != ele[11][23];
    ele[6][23] != ele[12][23];
    ele[6][23] != ele[13][23];
    ele[6][23] != ele[14][23];
    ele[6][23] != ele[15][23];
    ele[6][23] != ele[16][23];
    ele[6][23] != ele[17][23];
    ele[6][23] != ele[18][23];
    ele[6][23] != ele[19][23];
    ele[6][23] != ele[20][23];
    ele[6][23] != ele[21][23];
    ele[6][23] != ele[22][23];
    ele[6][23] != ele[23][23];
    ele[6][23] != ele[24][23];
    ele[6][23] != ele[25][23];
    ele[6][23] != ele[26][23];
    ele[6][23] != ele[27][23];
    ele[6][23] != ele[28][23];
    ele[6][23] != ele[29][23];
    ele[6][23] != ele[30][23];
    ele[6][23] != ele[31][23];
    ele[6][23] != ele[32][23];
    ele[6][23] != ele[33][23];
    ele[6][23] != ele[34][23];
    ele[6][23] != ele[35][23];
    ele[6][23] != ele[6][24];
    ele[6][23] != ele[6][25];
    ele[6][23] != ele[6][26];
    ele[6][23] != ele[6][27];
    ele[6][23] != ele[6][28];
    ele[6][23] != ele[6][29];
    ele[6][23] != ele[6][30];
    ele[6][23] != ele[6][31];
    ele[6][23] != ele[6][32];
    ele[6][23] != ele[6][33];
    ele[6][23] != ele[6][34];
    ele[6][23] != ele[6][35];
    ele[6][23] != ele[7][18];
    ele[6][23] != ele[7][19];
    ele[6][23] != ele[7][20];
    ele[6][23] != ele[7][21];
    ele[6][23] != ele[7][22];
    ele[6][23] != ele[7][23];
    ele[6][23] != ele[8][18];
    ele[6][23] != ele[8][19];
    ele[6][23] != ele[8][20];
    ele[6][23] != ele[8][21];
    ele[6][23] != ele[8][22];
    ele[6][23] != ele[8][23];
    ele[6][23] != ele[9][18];
    ele[6][23] != ele[9][19];
    ele[6][23] != ele[9][20];
    ele[6][23] != ele[9][21];
    ele[6][23] != ele[9][22];
    ele[6][23] != ele[9][23];
    ele[6][24] != ele[10][24];
    ele[6][24] != ele[10][25];
    ele[6][24] != ele[10][26];
    ele[6][24] != ele[10][27];
    ele[6][24] != ele[10][28];
    ele[6][24] != ele[10][29];
    ele[6][24] != ele[11][24];
    ele[6][24] != ele[11][25];
    ele[6][24] != ele[11][26];
    ele[6][24] != ele[11][27];
    ele[6][24] != ele[11][28];
    ele[6][24] != ele[11][29];
    ele[6][24] != ele[12][24];
    ele[6][24] != ele[13][24];
    ele[6][24] != ele[14][24];
    ele[6][24] != ele[15][24];
    ele[6][24] != ele[16][24];
    ele[6][24] != ele[17][24];
    ele[6][24] != ele[18][24];
    ele[6][24] != ele[19][24];
    ele[6][24] != ele[20][24];
    ele[6][24] != ele[21][24];
    ele[6][24] != ele[22][24];
    ele[6][24] != ele[23][24];
    ele[6][24] != ele[24][24];
    ele[6][24] != ele[25][24];
    ele[6][24] != ele[26][24];
    ele[6][24] != ele[27][24];
    ele[6][24] != ele[28][24];
    ele[6][24] != ele[29][24];
    ele[6][24] != ele[30][24];
    ele[6][24] != ele[31][24];
    ele[6][24] != ele[32][24];
    ele[6][24] != ele[33][24];
    ele[6][24] != ele[34][24];
    ele[6][24] != ele[35][24];
    ele[6][24] != ele[6][25];
    ele[6][24] != ele[6][26];
    ele[6][24] != ele[6][27];
    ele[6][24] != ele[6][28];
    ele[6][24] != ele[6][29];
    ele[6][24] != ele[6][30];
    ele[6][24] != ele[6][31];
    ele[6][24] != ele[6][32];
    ele[6][24] != ele[6][33];
    ele[6][24] != ele[6][34];
    ele[6][24] != ele[6][35];
    ele[6][24] != ele[7][24];
    ele[6][24] != ele[7][25];
    ele[6][24] != ele[7][26];
    ele[6][24] != ele[7][27];
    ele[6][24] != ele[7][28];
    ele[6][24] != ele[7][29];
    ele[6][24] != ele[8][24];
    ele[6][24] != ele[8][25];
    ele[6][24] != ele[8][26];
    ele[6][24] != ele[8][27];
    ele[6][24] != ele[8][28];
    ele[6][24] != ele[8][29];
    ele[6][24] != ele[9][24];
    ele[6][24] != ele[9][25];
    ele[6][24] != ele[9][26];
    ele[6][24] != ele[9][27];
    ele[6][24] != ele[9][28];
    ele[6][24] != ele[9][29];
    ele[6][25] != ele[10][24];
    ele[6][25] != ele[10][25];
    ele[6][25] != ele[10][26];
    ele[6][25] != ele[10][27];
    ele[6][25] != ele[10][28];
    ele[6][25] != ele[10][29];
    ele[6][25] != ele[11][24];
    ele[6][25] != ele[11][25];
    ele[6][25] != ele[11][26];
    ele[6][25] != ele[11][27];
    ele[6][25] != ele[11][28];
    ele[6][25] != ele[11][29];
    ele[6][25] != ele[12][25];
    ele[6][25] != ele[13][25];
    ele[6][25] != ele[14][25];
    ele[6][25] != ele[15][25];
    ele[6][25] != ele[16][25];
    ele[6][25] != ele[17][25];
    ele[6][25] != ele[18][25];
    ele[6][25] != ele[19][25];
    ele[6][25] != ele[20][25];
    ele[6][25] != ele[21][25];
    ele[6][25] != ele[22][25];
    ele[6][25] != ele[23][25];
    ele[6][25] != ele[24][25];
    ele[6][25] != ele[25][25];
    ele[6][25] != ele[26][25];
    ele[6][25] != ele[27][25];
    ele[6][25] != ele[28][25];
    ele[6][25] != ele[29][25];
    ele[6][25] != ele[30][25];
    ele[6][25] != ele[31][25];
    ele[6][25] != ele[32][25];
    ele[6][25] != ele[33][25];
    ele[6][25] != ele[34][25];
    ele[6][25] != ele[35][25];
    ele[6][25] != ele[6][26];
    ele[6][25] != ele[6][27];
    ele[6][25] != ele[6][28];
    ele[6][25] != ele[6][29];
    ele[6][25] != ele[6][30];
    ele[6][25] != ele[6][31];
    ele[6][25] != ele[6][32];
    ele[6][25] != ele[6][33];
    ele[6][25] != ele[6][34];
    ele[6][25] != ele[6][35];
    ele[6][25] != ele[7][24];
    ele[6][25] != ele[7][25];
    ele[6][25] != ele[7][26];
    ele[6][25] != ele[7][27];
    ele[6][25] != ele[7][28];
    ele[6][25] != ele[7][29];
    ele[6][25] != ele[8][24];
    ele[6][25] != ele[8][25];
    ele[6][25] != ele[8][26];
    ele[6][25] != ele[8][27];
    ele[6][25] != ele[8][28];
    ele[6][25] != ele[8][29];
    ele[6][25] != ele[9][24];
    ele[6][25] != ele[9][25];
    ele[6][25] != ele[9][26];
    ele[6][25] != ele[9][27];
    ele[6][25] != ele[9][28];
    ele[6][25] != ele[9][29];
    ele[6][26] != ele[10][24];
    ele[6][26] != ele[10][25];
    ele[6][26] != ele[10][26];
    ele[6][26] != ele[10][27];
    ele[6][26] != ele[10][28];
    ele[6][26] != ele[10][29];
    ele[6][26] != ele[11][24];
    ele[6][26] != ele[11][25];
    ele[6][26] != ele[11][26];
    ele[6][26] != ele[11][27];
    ele[6][26] != ele[11][28];
    ele[6][26] != ele[11][29];
    ele[6][26] != ele[12][26];
    ele[6][26] != ele[13][26];
    ele[6][26] != ele[14][26];
    ele[6][26] != ele[15][26];
    ele[6][26] != ele[16][26];
    ele[6][26] != ele[17][26];
    ele[6][26] != ele[18][26];
    ele[6][26] != ele[19][26];
    ele[6][26] != ele[20][26];
    ele[6][26] != ele[21][26];
    ele[6][26] != ele[22][26];
    ele[6][26] != ele[23][26];
    ele[6][26] != ele[24][26];
    ele[6][26] != ele[25][26];
    ele[6][26] != ele[26][26];
    ele[6][26] != ele[27][26];
    ele[6][26] != ele[28][26];
    ele[6][26] != ele[29][26];
    ele[6][26] != ele[30][26];
    ele[6][26] != ele[31][26];
    ele[6][26] != ele[32][26];
    ele[6][26] != ele[33][26];
    ele[6][26] != ele[34][26];
    ele[6][26] != ele[35][26];
    ele[6][26] != ele[6][27];
    ele[6][26] != ele[6][28];
    ele[6][26] != ele[6][29];
    ele[6][26] != ele[6][30];
    ele[6][26] != ele[6][31];
    ele[6][26] != ele[6][32];
    ele[6][26] != ele[6][33];
    ele[6][26] != ele[6][34];
    ele[6][26] != ele[6][35];
    ele[6][26] != ele[7][24];
    ele[6][26] != ele[7][25];
    ele[6][26] != ele[7][26];
    ele[6][26] != ele[7][27];
    ele[6][26] != ele[7][28];
    ele[6][26] != ele[7][29];
    ele[6][26] != ele[8][24];
    ele[6][26] != ele[8][25];
    ele[6][26] != ele[8][26];
    ele[6][26] != ele[8][27];
    ele[6][26] != ele[8][28];
    ele[6][26] != ele[8][29];
    ele[6][26] != ele[9][24];
    ele[6][26] != ele[9][25];
    ele[6][26] != ele[9][26];
    ele[6][26] != ele[9][27];
    ele[6][26] != ele[9][28];
    ele[6][26] != ele[9][29];
    ele[6][27] != ele[10][24];
    ele[6][27] != ele[10][25];
    ele[6][27] != ele[10][26];
    ele[6][27] != ele[10][27];
    ele[6][27] != ele[10][28];
    ele[6][27] != ele[10][29];
    ele[6][27] != ele[11][24];
    ele[6][27] != ele[11][25];
    ele[6][27] != ele[11][26];
    ele[6][27] != ele[11][27];
    ele[6][27] != ele[11][28];
    ele[6][27] != ele[11][29];
    ele[6][27] != ele[12][27];
    ele[6][27] != ele[13][27];
    ele[6][27] != ele[14][27];
    ele[6][27] != ele[15][27];
    ele[6][27] != ele[16][27];
    ele[6][27] != ele[17][27];
    ele[6][27] != ele[18][27];
    ele[6][27] != ele[19][27];
    ele[6][27] != ele[20][27];
    ele[6][27] != ele[21][27];
    ele[6][27] != ele[22][27];
    ele[6][27] != ele[23][27];
    ele[6][27] != ele[24][27];
    ele[6][27] != ele[25][27];
    ele[6][27] != ele[26][27];
    ele[6][27] != ele[27][27];
    ele[6][27] != ele[28][27];
    ele[6][27] != ele[29][27];
    ele[6][27] != ele[30][27];
    ele[6][27] != ele[31][27];
    ele[6][27] != ele[32][27];
    ele[6][27] != ele[33][27];
    ele[6][27] != ele[34][27];
    ele[6][27] != ele[35][27];
    ele[6][27] != ele[6][28];
    ele[6][27] != ele[6][29];
    ele[6][27] != ele[6][30];
    ele[6][27] != ele[6][31];
    ele[6][27] != ele[6][32];
    ele[6][27] != ele[6][33];
    ele[6][27] != ele[6][34];
    ele[6][27] != ele[6][35];
    ele[6][27] != ele[7][24];
    ele[6][27] != ele[7][25];
    ele[6][27] != ele[7][26];
    ele[6][27] != ele[7][27];
    ele[6][27] != ele[7][28];
    ele[6][27] != ele[7][29];
    ele[6][27] != ele[8][24];
    ele[6][27] != ele[8][25];
    ele[6][27] != ele[8][26];
    ele[6][27] != ele[8][27];
    ele[6][27] != ele[8][28];
    ele[6][27] != ele[8][29];
    ele[6][27] != ele[9][24];
    ele[6][27] != ele[9][25];
    ele[6][27] != ele[9][26];
    ele[6][27] != ele[9][27];
    ele[6][27] != ele[9][28];
    ele[6][27] != ele[9][29];
    ele[6][28] != ele[10][24];
    ele[6][28] != ele[10][25];
    ele[6][28] != ele[10][26];
    ele[6][28] != ele[10][27];
    ele[6][28] != ele[10][28];
    ele[6][28] != ele[10][29];
    ele[6][28] != ele[11][24];
    ele[6][28] != ele[11][25];
    ele[6][28] != ele[11][26];
    ele[6][28] != ele[11][27];
    ele[6][28] != ele[11][28];
    ele[6][28] != ele[11][29];
    ele[6][28] != ele[12][28];
    ele[6][28] != ele[13][28];
    ele[6][28] != ele[14][28];
    ele[6][28] != ele[15][28];
    ele[6][28] != ele[16][28];
    ele[6][28] != ele[17][28];
    ele[6][28] != ele[18][28];
    ele[6][28] != ele[19][28];
    ele[6][28] != ele[20][28];
    ele[6][28] != ele[21][28];
    ele[6][28] != ele[22][28];
    ele[6][28] != ele[23][28];
    ele[6][28] != ele[24][28];
    ele[6][28] != ele[25][28];
    ele[6][28] != ele[26][28];
    ele[6][28] != ele[27][28];
    ele[6][28] != ele[28][28];
    ele[6][28] != ele[29][28];
    ele[6][28] != ele[30][28];
    ele[6][28] != ele[31][28];
    ele[6][28] != ele[32][28];
    ele[6][28] != ele[33][28];
    ele[6][28] != ele[34][28];
    ele[6][28] != ele[35][28];
    ele[6][28] != ele[6][29];
    ele[6][28] != ele[6][30];
    ele[6][28] != ele[6][31];
    ele[6][28] != ele[6][32];
    ele[6][28] != ele[6][33];
    ele[6][28] != ele[6][34];
    ele[6][28] != ele[6][35];
    ele[6][28] != ele[7][24];
    ele[6][28] != ele[7][25];
    ele[6][28] != ele[7][26];
    ele[6][28] != ele[7][27];
    ele[6][28] != ele[7][28];
    ele[6][28] != ele[7][29];
    ele[6][28] != ele[8][24];
    ele[6][28] != ele[8][25];
    ele[6][28] != ele[8][26];
    ele[6][28] != ele[8][27];
    ele[6][28] != ele[8][28];
    ele[6][28] != ele[8][29];
    ele[6][28] != ele[9][24];
    ele[6][28] != ele[9][25];
    ele[6][28] != ele[9][26];
    ele[6][28] != ele[9][27];
    ele[6][28] != ele[9][28];
    ele[6][28] != ele[9][29];
    ele[6][29] != ele[10][24];
    ele[6][29] != ele[10][25];
    ele[6][29] != ele[10][26];
    ele[6][29] != ele[10][27];
    ele[6][29] != ele[10][28];
    ele[6][29] != ele[10][29];
    ele[6][29] != ele[11][24];
    ele[6][29] != ele[11][25];
    ele[6][29] != ele[11][26];
    ele[6][29] != ele[11][27];
    ele[6][29] != ele[11][28];
    ele[6][29] != ele[11][29];
    ele[6][29] != ele[12][29];
    ele[6][29] != ele[13][29];
    ele[6][29] != ele[14][29];
    ele[6][29] != ele[15][29];
    ele[6][29] != ele[16][29];
    ele[6][29] != ele[17][29];
    ele[6][29] != ele[18][29];
    ele[6][29] != ele[19][29];
    ele[6][29] != ele[20][29];
    ele[6][29] != ele[21][29];
    ele[6][29] != ele[22][29];
    ele[6][29] != ele[23][29];
    ele[6][29] != ele[24][29];
    ele[6][29] != ele[25][29];
    ele[6][29] != ele[26][29];
    ele[6][29] != ele[27][29];
    ele[6][29] != ele[28][29];
    ele[6][29] != ele[29][29];
    ele[6][29] != ele[30][29];
    ele[6][29] != ele[31][29];
    ele[6][29] != ele[32][29];
    ele[6][29] != ele[33][29];
    ele[6][29] != ele[34][29];
    ele[6][29] != ele[35][29];
    ele[6][29] != ele[6][30];
    ele[6][29] != ele[6][31];
    ele[6][29] != ele[6][32];
    ele[6][29] != ele[6][33];
    ele[6][29] != ele[6][34];
    ele[6][29] != ele[6][35];
    ele[6][29] != ele[7][24];
    ele[6][29] != ele[7][25];
    ele[6][29] != ele[7][26];
    ele[6][29] != ele[7][27];
    ele[6][29] != ele[7][28];
    ele[6][29] != ele[7][29];
    ele[6][29] != ele[8][24];
    ele[6][29] != ele[8][25];
    ele[6][29] != ele[8][26];
    ele[6][29] != ele[8][27];
    ele[6][29] != ele[8][28];
    ele[6][29] != ele[8][29];
    ele[6][29] != ele[9][24];
    ele[6][29] != ele[9][25];
    ele[6][29] != ele[9][26];
    ele[6][29] != ele[9][27];
    ele[6][29] != ele[9][28];
    ele[6][29] != ele[9][29];
    ele[6][3] != ele[10][0];
    ele[6][3] != ele[10][1];
    ele[6][3] != ele[10][2];
    ele[6][3] != ele[10][3];
    ele[6][3] != ele[10][4];
    ele[6][3] != ele[10][5];
    ele[6][3] != ele[11][0];
    ele[6][3] != ele[11][1];
    ele[6][3] != ele[11][2];
    ele[6][3] != ele[11][3];
    ele[6][3] != ele[11][4];
    ele[6][3] != ele[11][5];
    ele[6][3] != ele[12][3];
    ele[6][3] != ele[13][3];
    ele[6][3] != ele[14][3];
    ele[6][3] != ele[15][3];
    ele[6][3] != ele[16][3];
    ele[6][3] != ele[17][3];
    ele[6][3] != ele[18][3];
    ele[6][3] != ele[19][3];
    ele[6][3] != ele[20][3];
    ele[6][3] != ele[21][3];
    ele[6][3] != ele[22][3];
    ele[6][3] != ele[23][3];
    ele[6][3] != ele[24][3];
    ele[6][3] != ele[25][3];
    ele[6][3] != ele[26][3];
    ele[6][3] != ele[27][3];
    ele[6][3] != ele[28][3];
    ele[6][3] != ele[29][3];
    ele[6][3] != ele[30][3];
    ele[6][3] != ele[31][3];
    ele[6][3] != ele[32][3];
    ele[6][3] != ele[33][3];
    ele[6][3] != ele[34][3];
    ele[6][3] != ele[35][3];
    ele[6][3] != ele[6][10];
    ele[6][3] != ele[6][11];
    ele[6][3] != ele[6][12];
    ele[6][3] != ele[6][13];
    ele[6][3] != ele[6][14];
    ele[6][3] != ele[6][15];
    ele[6][3] != ele[6][16];
    ele[6][3] != ele[6][17];
    ele[6][3] != ele[6][18];
    ele[6][3] != ele[6][19];
    ele[6][3] != ele[6][20];
    ele[6][3] != ele[6][21];
    ele[6][3] != ele[6][22];
    ele[6][3] != ele[6][23];
    ele[6][3] != ele[6][24];
    ele[6][3] != ele[6][25];
    ele[6][3] != ele[6][26];
    ele[6][3] != ele[6][27];
    ele[6][3] != ele[6][28];
    ele[6][3] != ele[6][29];
    ele[6][3] != ele[6][30];
    ele[6][3] != ele[6][31];
    ele[6][3] != ele[6][32];
    ele[6][3] != ele[6][33];
    ele[6][3] != ele[6][34];
    ele[6][3] != ele[6][35];
    ele[6][3] != ele[6][4];
    ele[6][3] != ele[6][5];
    ele[6][3] != ele[6][6];
    ele[6][3] != ele[6][7];
    ele[6][3] != ele[6][8];
    ele[6][3] != ele[6][9];
    ele[6][3] != ele[7][0];
    ele[6][3] != ele[7][1];
    ele[6][3] != ele[7][2];
    ele[6][3] != ele[7][3];
    ele[6][3] != ele[7][4];
    ele[6][3] != ele[7][5];
    ele[6][3] != ele[8][0];
    ele[6][3] != ele[8][1];
    ele[6][3] != ele[8][2];
    ele[6][3] != ele[8][3];
    ele[6][3] != ele[8][4];
    ele[6][3] != ele[8][5];
    ele[6][3] != ele[9][0];
    ele[6][3] != ele[9][1];
    ele[6][3] != ele[9][2];
    ele[6][3] != ele[9][3];
    ele[6][3] != ele[9][4];
    ele[6][3] != ele[9][5];
    ele[6][30] != ele[10][30];
    ele[6][30] != ele[10][31];
    ele[6][30] != ele[10][32];
    ele[6][30] != ele[10][33];
    ele[6][30] != ele[10][34];
    ele[6][30] != ele[10][35];
    ele[6][30] != ele[11][30];
    ele[6][30] != ele[11][31];
    ele[6][30] != ele[11][32];
    ele[6][30] != ele[11][33];
    ele[6][30] != ele[11][34];
    ele[6][30] != ele[11][35];
    ele[6][30] != ele[12][30];
    ele[6][30] != ele[13][30];
    ele[6][30] != ele[14][30];
    ele[6][30] != ele[15][30];
    ele[6][30] != ele[16][30];
    ele[6][30] != ele[17][30];
    ele[6][30] != ele[18][30];
    ele[6][30] != ele[19][30];
    ele[6][30] != ele[20][30];
    ele[6][30] != ele[21][30];
    ele[6][30] != ele[22][30];
    ele[6][30] != ele[23][30];
    ele[6][30] != ele[24][30];
    ele[6][30] != ele[25][30];
    ele[6][30] != ele[26][30];
    ele[6][30] != ele[27][30];
    ele[6][30] != ele[28][30];
    ele[6][30] != ele[29][30];
    ele[6][30] != ele[30][30];
    ele[6][30] != ele[31][30];
    ele[6][30] != ele[32][30];
    ele[6][30] != ele[33][30];
    ele[6][30] != ele[34][30];
    ele[6][30] != ele[35][30];
    ele[6][30] != ele[6][31];
    ele[6][30] != ele[6][32];
    ele[6][30] != ele[6][33];
    ele[6][30] != ele[6][34];
    ele[6][30] != ele[6][35];
    ele[6][30] != ele[7][30];
    ele[6][30] != ele[7][31];
    ele[6][30] != ele[7][32];
    ele[6][30] != ele[7][33];
    ele[6][30] != ele[7][34];
    ele[6][30] != ele[7][35];
    ele[6][30] != ele[8][30];
    ele[6][30] != ele[8][31];
    ele[6][30] != ele[8][32];
    ele[6][30] != ele[8][33];
    ele[6][30] != ele[8][34];
    ele[6][30] != ele[8][35];
    ele[6][30] != ele[9][30];
    ele[6][30] != ele[9][31];
    ele[6][30] != ele[9][32];
    ele[6][30] != ele[9][33];
    ele[6][30] != ele[9][34];
    ele[6][30] != ele[9][35];
    ele[6][31] != ele[10][30];
    ele[6][31] != ele[10][31];
    ele[6][31] != ele[10][32];
    ele[6][31] != ele[10][33];
    ele[6][31] != ele[10][34];
    ele[6][31] != ele[10][35];
    ele[6][31] != ele[11][30];
    ele[6][31] != ele[11][31];
    ele[6][31] != ele[11][32];
    ele[6][31] != ele[11][33];
    ele[6][31] != ele[11][34];
    ele[6][31] != ele[11][35];
    ele[6][31] != ele[12][31];
    ele[6][31] != ele[13][31];
    ele[6][31] != ele[14][31];
    ele[6][31] != ele[15][31];
    ele[6][31] != ele[16][31];
    ele[6][31] != ele[17][31];
    ele[6][31] != ele[18][31];
    ele[6][31] != ele[19][31];
    ele[6][31] != ele[20][31];
    ele[6][31] != ele[21][31];
    ele[6][31] != ele[22][31];
    ele[6][31] != ele[23][31];
    ele[6][31] != ele[24][31];
    ele[6][31] != ele[25][31];
    ele[6][31] != ele[26][31];
    ele[6][31] != ele[27][31];
    ele[6][31] != ele[28][31];
    ele[6][31] != ele[29][31];
    ele[6][31] != ele[30][31];
    ele[6][31] != ele[31][31];
    ele[6][31] != ele[32][31];
    ele[6][31] != ele[33][31];
    ele[6][31] != ele[34][31];
    ele[6][31] != ele[35][31];
    ele[6][31] != ele[6][32];
    ele[6][31] != ele[6][33];
    ele[6][31] != ele[6][34];
    ele[6][31] != ele[6][35];
    ele[6][31] != ele[7][30];
    ele[6][31] != ele[7][31];
    ele[6][31] != ele[7][32];
    ele[6][31] != ele[7][33];
    ele[6][31] != ele[7][34];
    ele[6][31] != ele[7][35];
    ele[6][31] != ele[8][30];
    ele[6][31] != ele[8][31];
    ele[6][31] != ele[8][32];
    ele[6][31] != ele[8][33];
    ele[6][31] != ele[8][34];
    ele[6][31] != ele[8][35];
    ele[6][31] != ele[9][30];
    ele[6][31] != ele[9][31];
    ele[6][31] != ele[9][32];
    ele[6][31] != ele[9][33];
    ele[6][31] != ele[9][34];
    ele[6][31] != ele[9][35];
    ele[6][32] != ele[10][30];
    ele[6][32] != ele[10][31];
    ele[6][32] != ele[10][32];
    ele[6][32] != ele[10][33];
    ele[6][32] != ele[10][34];
    ele[6][32] != ele[10][35];
    ele[6][32] != ele[11][30];
    ele[6][32] != ele[11][31];
    ele[6][32] != ele[11][32];
    ele[6][32] != ele[11][33];
    ele[6][32] != ele[11][34];
    ele[6][32] != ele[11][35];
    ele[6][32] != ele[12][32];
    ele[6][32] != ele[13][32];
    ele[6][32] != ele[14][32];
    ele[6][32] != ele[15][32];
    ele[6][32] != ele[16][32];
    ele[6][32] != ele[17][32];
    ele[6][32] != ele[18][32];
    ele[6][32] != ele[19][32];
    ele[6][32] != ele[20][32];
    ele[6][32] != ele[21][32];
    ele[6][32] != ele[22][32];
    ele[6][32] != ele[23][32];
    ele[6][32] != ele[24][32];
    ele[6][32] != ele[25][32];
    ele[6][32] != ele[26][32];
    ele[6][32] != ele[27][32];
    ele[6][32] != ele[28][32];
    ele[6][32] != ele[29][32];
    ele[6][32] != ele[30][32];
    ele[6][32] != ele[31][32];
    ele[6][32] != ele[32][32];
    ele[6][32] != ele[33][32];
    ele[6][32] != ele[34][32];
    ele[6][32] != ele[35][32];
    ele[6][32] != ele[6][33];
    ele[6][32] != ele[6][34];
    ele[6][32] != ele[6][35];
    ele[6][32] != ele[7][30];
    ele[6][32] != ele[7][31];
    ele[6][32] != ele[7][32];
    ele[6][32] != ele[7][33];
    ele[6][32] != ele[7][34];
    ele[6][32] != ele[7][35];
    ele[6][32] != ele[8][30];
    ele[6][32] != ele[8][31];
    ele[6][32] != ele[8][32];
    ele[6][32] != ele[8][33];
    ele[6][32] != ele[8][34];
    ele[6][32] != ele[8][35];
    ele[6][32] != ele[9][30];
    ele[6][32] != ele[9][31];
    ele[6][32] != ele[9][32];
    ele[6][32] != ele[9][33];
    ele[6][32] != ele[9][34];
    ele[6][32] != ele[9][35];
    ele[6][33] != ele[10][30];
    ele[6][33] != ele[10][31];
    ele[6][33] != ele[10][32];
    ele[6][33] != ele[10][33];
    ele[6][33] != ele[10][34];
    ele[6][33] != ele[10][35];
    ele[6][33] != ele[11][30];
    ele[6][33] != ele[11][31];
    ele[6][33] != ele[11][32];
    ele[6][33] != ele[11][33];
    ele[6][33] != ele[11][34];
    ele[6][33] != ele[11][35];
    ele[6][33] != ele[12][33];
    ele[6][33] != ele[13][33];
    ele[6][33] != ele[14][33];
    ele[6][33] != ele[15][33];
    ele[6][33] != ele[16][33];
    ele[6][33] != ele[17][33];
    ele[6][33] != ele[18][33];
    ele[6][33] != ele[19][33];
    ele[6][33] != ele[20][33];
    ele[6][33] != ele[21][33];
    ele[6][33] != ele[22][33];
    ele[6][33] != ele[23][33];
    ele[6][33] != ele[24][33];
    ele[6][33] != ele[25][33];
    ele[6][33] != ele[26][33];
    ele[6][33] != ele[27][33];
    ele[6][33] != ele[28][33];
    ele[6][33] != ele[29][33];
    ele[6][33] != ele[30][33];
    ele[6][33] != ele[31][33];
    ele[6][33] != ele[32][33];
    ele[6][33] != ele[33][33];
    ele[6][33] != ele[34][33];
    ele[6][33] != ele[35][33];
    ele[6][33] != ele[6][34];
    ele[6][33] != ele[6][35];
    ele[6][33] != ele[7][30];
    ele[6][33] != ele[7][31];
    ele[6][33] != ele[7][32];
    ele[6][33] != ele[7][33];
    ele[6][33] != ele[7][34];
    ele[6][33] != ele[7][35];
    ele[6][33] != ele[8][30];
    ele[6][33] != ele[8][31];
    ele[6][33] != ele[8][32];
    ele[6][33] != ele[8][33];
    ele[6][33] != ele[8][34];
    ele[6][33] != ele[8][35];
    ele[6][33] != ele[9][30];
    ele[6][33] != ele[9][31];
    ele[6][33] != ele[9][32];
    ele[6][33] != ele[9][33];
    ele[6][33] != ele[9][34];
    ele[6][33] != ele[9][35];
    ele[6][34] != ele[10][30];
    ele[6][34] != ele[10][31];
    ele[6][34] != ele[10][32];
    ele[6][34] != ele[10][33];
    ele[6][34] != ele[10][34];
    ele[6][34] != ele[10][35];
    ele[6][34] != ele[11][30];
    ele[6][34] != ele[11][31];
    ele[6][34] != ele[11][32];
    ele[6][34] != ele[11][33];
    ele[6][34] != ele[11][34];
    ele[6][34] != ele[11][35];
    ele[6][34] != ele[12][34];
    ele[6][34] != ele[13][34];
    ele[6][34] != ele[14][34];
    ele[6][34] != ele[15][34];
    ele[6][34] != ele[16][34];
    ele[6][34] != ele[17][34];
    ele[6][34] != ele[18][34];
    ele[6][34] != ele[19][34];
    ele[6][34] != ele[20][34];
    ele[6][34] != ele[21][34];
    ele[6][34] != ele[22][34];
    ele[6][34] != ele[23][34];
    ele[6][34] != ele[24][34];
    ele[6][34] != ele[25][34];
    ele[6][34] != ele[26][34];
    ele[6][34] != ele[27][34];
    ele[6][34] != ele[28][34];
    ele[6][34] != ele[29][34];
    ele[6][34] != ele[30][34];
    ele[6][34] != ele[31][34];
    ele[6][34] != ele[32][34];
    ele[6][34] != ele[33][34];
    ele[6][34] != ele[34][34];
    ele[6][34] != ele[35][34];
    ele[6][34] != ele[6][35];
    ele[6][34] != ele[7][30];
    ele[6][34] != ele[7][31];
    ele[6][34] != ele[7][32];
    ele[6][34] != ele[7][33];
    ele[6][34] != ele[7][34];
    ele[6][34] != ele[7][35];
    ele[6][34] != ele[8][30];
    ele[6][34] != ele[8][31];
    ele[6][34] != ele[8][32];
    ele[6][34] != ele[8][33];
    ele[6][34] != ele[8][34];
    ele[6][34] != ele[8][35];
    ele[6][34] != ele[9][30];
    ele[6][34] != ele[9][31];
    ele[6][34] != ele[9][32];
    ele[6][34] != ele[9][33];
    ele[6][34] != ele[9][34];
    ele[6][34] != ele[9][35];
    ele[6][35] != ele[10][30];
    ele[6][35] != ele[10][31];
    ele[6][35] != ele[10][32];
    ele[6][35] != ele[10][33];
    ele[6][35] != ele[10][34];
    ele[6][35] != ele[10][35];
    ele[6][35] != ele[11][30];
    ele[6][35] != ele[11][31];
    ele[6][35] != ele[11][32];
    ele[6][35] != ele[11][33];
    ele[6][35] != ele[11][34];
    ele[6][35] != ele[11][35];
    ele[6][35] != ele[12][35];
    ele[6][35] != ele[13][35];
    ele[6][35] != ele[14][35];
    ele[6][35] != ele[15][35];
    ele[6][35] != ele[16][35];
    ele[6][35] != ele[17][35];
    ele[6][35] != ele[18][35];
    ele[6][35] != ele[19][35];
    ele[6][35] != ele[20][35];
    ele[6][35] != ele[21][35];
    ele[6][35] != ele[22][35];
    ele[6][35] != ele[23][35];
    ele[6][35] != ele[24][35];
    ele[6][35] != ele[25][35];
    ele[6][35] != ele[26][35];
    ele[6][35] != ele[27][35];
    ele[6][35] != ele[28][35];
    ele[6][35] != ele[29][35];
    ele[6][35] != ele[30][35];
    ele[6][35] != ele[31][35];
    ele[6][35] != ele[32][35];
    ele[6][35] != ele[33][35];
    ele[6][35] != ele[34][35];
    ele[6][35] != ele[35][35];
    ele[6][35] != ele[7][30];
    ele[6][35] != ele[7][31];
    ele[6][35] != ele[7][32];
    ele[6][35] != ele[7][33];
    ele[6][35] != ele[7][34];
    ele[6][35] != ele[7][35];
    ele[6][35] != ele[8][30];
    ele[6][35] != ele[8][31];
    ele[6][35] != ele[8][32];
    ele[6][35] != ele[8][33];
    ele[6][35] != ele[8][34];
    ele[6][35] != ele[8][35];
    ele[6][35] != ele[9][30];
    ele[6][35] != ele[9][31];
    ele[6][35] != ele[9][32];
    ele[6][35] != ele[9][33];
    ele[6][35] != ele[9][34];
    ele[6][35] != ele[9][35];
    ele[6][4] != ele[10][0];
    ele[6][4] != ele[10][1];
    ele[6][4] != ele[10][2];
    ele[6][4] != ele[10][3];
    ele[6][4] != ele[10][4];
    ele[6][4] != ele[10][5];
    ele[6][4] != ele[11][0];
    ele[6][4] != ele[11][1];
    ele[6][4] != ele[11][2];
    ele[6][4] != ele[11][3];
    ele[6][4] != ele[11][4];
    ele[6][4] != ele[11][5];
    ele[6][4] != ele[12][4];
    ele[6][4] != ele[13][4];
    ele[6][4] != ele[14][4];
    ele[6][4] != ele[15][4];
    ele[6][4] != ele[16][4];
    ele[6][4] != ele[17][4];
    ele[6][4] != ele[18][4];
    ele[6][4] != ele[19][4];
    ele[6][4] != ele[20][4];
    ele[6][4] != ele[21][4];
    ele[6][4] != ele[22][4];
    ele[6][4] != ele[23][4];
    ele[6][4] != ele[24][4];
    ele[6][4] != ele[25][4];
    ele[6][4] != ele[26][4];
    ele[6][4] != ele[27][4];
    ele[6][4] != ele[28][4];
    ele[6][4] != ele[29][4];
    ele[6][4] != ele[30][4];
    ele[6][4] != ele[31][4];
    ele[6][4] != ele[32][4];
    ele[6][4] != ele[33][4];
    ele[6][4] != ele[34][4];
    ele[6][4] != ele[35][4];
    ele[6][4] != ele[6][10];
    ele[6][4] != ele[6][11];
    ele[6][4] != ele[6][12];
    ele[6][4] != ele[6][13];
    ele[6][4] != ele[6][14];
    ele[6][4] != ele[6][15];
    ele[6][4] != ele[6][16];
    ele[6][4] != ele[6][17];
    ele[6][4] != ele[6][18];
    ele[6][4] != ele[6][19];
    ele[6][4] != ele[6][20];
    ele[6][4] != ele[6][21];
    ele[6][4] != ele[6][22];
    ele[6][4] != ele[6][23];
    ele[6][4] != ele[6][24];
    ele[6][4] != ele[6][25];
    ele[6][4] != ele[6][26];
    ele[6][4] != ele[6][27];
    ele[6][4] != ele[6][28];
    ele[6][4] != ele[6][29];
    ele[6][4] != ele[6][30];
    ele[6][4] != ele[6][31];
    ele[6][4] != ele[6][32];
    ele[6][4] != ele[6][33];
    ele[6][4] != ele[6][34];
    ele[6][4] != ele[6][35];
    ele[6][4] != ele[6][5];
    ele[6][4] != ele[6][6];
    ele[6][4] != ele[6][7];
    ele[6][4] != ele[6][8];
    ele[6][4] != ele[6][9];
    ele[6][4] != ele[7][0];
    ele[6][4] != ele[7][1];
    ele[6][4] != ele[7][2];
    ele[6][4] != ele[7][3];
    ele[6][4] != ele[7][4];
    ele[6][4] != ele[7][5];
    ele[6][4] != ele[8][0];
    ele[6][4] != ele[8][1];
    ele[6][4] != ele[8][2];
    ele[6][4] != ele[8][3];
    ele[6][4] != ele[8][4];
    ele[6][4] != ele[8][5];
    ele[6][4] != ele[9][0];
    ele[6][4] != ele[9][1];
    ele[6][4] != ele[9][2];
    ele[6][4] != ele[9][3];
    ele[6][4] != ele[9][4];
    ele[6][4] != ele[9][5];
    ele[6][5] != ele[10][0];
    ele[6][5] != ele[10][1];
    ele[6][5] != ele[10][2];
    ele[6][5] != ele[10][3];
    ele[6][5] != ele[10][4];
    ele[6][5] != ele[10][5];
    ele[6][5] != ele[11][0];
    ele[6][5] != ele[11][1];
    ele[6][5] != ele[11][2];
    ele[6][5] != ele[11][3];
    ele[6][5] != ele[11][4];
    ele[6][5] != ele[11][5];
    ele[6][5] != ele[12][5];
    ele[6][5] != ele[13][5];
    ele[6][5] != ele[14][5];
    ele[6][5] != ele[15][5];
    ele[6][5] != ele[16][5];
    ele[6][5] != ele[17][5];
    ele[6][5] != ele[18][5];
    ele[6][5] != ele[19][5];
    ele[6][5] != ele[20][5];
    ele[6][5] != ele[21][5];
    ele[6][5] != ele[22][5];
    ele[6][5] != ele[23][5];
    ele[6][5] != ele[24][5];
    ele[6][5] != ele[25][5];
    ele[6][5] != ele[26][5];
    ele[6][5] != ele[27][5];
    ele[6][5] != ele[28][5];
    ele[6][5] != ele[29][5];
    ele[6][5] != ele[30][5];
    ele[6][5] != ele[31][5];
    ele[6][5] != ele[32][5];
    ele[6][5] != ele[33][5];
    ele[6][5] != ele[34][5];
    ele[6][5] != ele[35][5];
    ele[6][5] != ele[6][10];
    ele[6][5] != ele[6][11];
    ele[6][5] != ele[6][12];
    ele[6][5] != ele[6][13];
    ele[6][5] != ele[6][14];
    ele[6][5] != ele[6][15];
    ele[6][5] != ele[6][16];
    ele[6][5] != ele[6][17];
    ele[6][5] != ele[6][18];
    ele[6][5] != ele[6][19];
    ele[6][5] != ele[6][20];
    ele[6][5] != ele[6][21];
    ele[6][5] != ele[6][22];
    ele[6][5] != ele[6][23];
    ele[6][5] != ele[6][24];
    ele[6][5] != ele[6][25];
    ele[6][5] != ele[6][26];
    ele[6][5] != ele[6][27];
    ele[6][5] != ele[6][28];
    ele[6][5] != ele[6][29];
    ele[6][5] != ele[6][30];
    ele[6][5] != ele[6][31];
    ele[6][5] != ele[6][32];
    ele[6][5] != ele[6][33];
    ele[6][5] != ele[6][34];
    ele[6][5] != ele[6][35];
    ele[6][5] != ele[6][6];
    ele[6][5] != ele[6][7];
    ele[6][5] != ele[6][8];
    ele[6][5] != ele[6][9];
    ele[6][5] != ele[7][0];
    ele[6][5] != ele[7][1];
    ele[6][5] != ele[7][2];
    ele[6][5] != ele[7][3];
    ele[6][5] != ele[7][4];
    ele[6][5] != ele[7][5];
    ele[6][5] != ele[8][0];
    ele[6][5] != ele[8][1];
    ele[6][5] != ele[8][2];
    ele[6][5] != ele[8][3];
    ele[6][5] != ele[8][4];
    ele[6][5] != ele[8][5];
    ele[6][5] != ele[9][0];
    ele[6][5] != ele[9][1];
    ele[6][5] != ele[9][2];
    ele[6][5] != ele[9][3];
    ele[6][5] != ele[9][4];
    ele[6][5] != ele[9][5];
    ele[6][6] != ele[10][10];
    ele[6][6] != ele[10][11];
    ele[6][6] != ele[10][6];
    ele[6][6] != ele[10][7];
    ele[6][6] != ele[10][8];
    ele[6][6] != ele[10][9];
    ele[6][6] != ele[11][10];
    ele[6][6] != ele[11][11];
    ele[6][6] != ele[11][6];
    ele[6][6] != ele[11][7];
    ele[6][6] != ele[11][8];
    ele[6][6] != ele[11][9];
    ele[6][6] != ele[12][6];
    ele[6][6] != ele[13][6];
    ele[6][6] != ele[14][6];
    ele[6][6] != ele[15][6];
    ele[6][6] != ele[16][6];
    ele[6][6] != ele[17][6];
    ele[6][6] != ele[18][6];
    ele[6][6] != ele[19][6];
    ele[6][6] != ele[20][6];
    ele[6][6] != ele[21][6];
    ele[6][6] != ele[22][6];
    ele[6][6] != ele[23][6];
    ele[6][6] != ele[24][6];
    ele[6][6] != ele[25][6];
    ele[6][6] != ele[26][6];
    ele[6][6] != ele[27][6];
    ele[6][6] != ele[28][6];
    ele[6][6] != ele[29][6];
    ele[6][6] != ele[30][6];
    ele[6][6] != ele[31][6];
    ele[6][6] != ele[32][6];
    ele[6][6] != ele[33][6];
    ele[6][6] != ele[34][6];
    ele[6][6] != ele[35][6];
    ele[6][6] != ele[6][10];
    ele[6][6] != ele[6][11];
    ele[6][6] != ele[6][12];
    ele[6][6] != ele[6][13];
    ele[6][6] != ele[6][14];
    ele[6][6] != ele[6][15];
    ele[6][6] != ele[6][16];
    ele[6][6] != ele[6][17];
    ele[6][6] != ele[6][18];
    ele[6][6] != ele[6][19];
    ele[6][6] != ele[6][20];
    ele[6][6] != ele[6][21];
    ele[6][6] != ele[6][22];
    ele[6][6] != ele[6][23];
    ele[6][6] != ele[6][24];
    ele[6][6] != ele[6][25];
    ele[6][6] != ele[6][26];
    ele[6][6] != ele[6][27];
    ele[6][6] != ele[6][28];
    ele[6][6] != ele[6][29];
    ele[6][6] != ele[6][30];
    ele[6][6] != ele[6][31];
    ele[6][6] != ele[6][32];
    ele[6][6] != ele[6][33];
    ele[6][6] != ele[6][34];
    ele[6][6] != ele[6][35];
    ele[6][6] != ele[6][7];
    ele[6][6] != ele[6][8];
    ele[6][6] != ele[6][9];
    ele[6][6] != ele[7][10];
    ele[6][6] != ele[7][11];
    ele[6][6] != ele[7][6];
    ele[6][6] != ele[7][7];
    ele[6][6] != ele[7][8];
    ele[6][6] != ele[7][9];
    ele[6][6] != ele[8][10];
    ele[6][6] != ele[8][11];
    ele[6][6] != ele[8][6];
    ele[6][6] != ele[8][7];
    ele[6][6] != ele[8][8];
    ele[6][6] != ele[8][9];
    ele[6][6] != ele[9][10];
    ele[6][6] != ele[9][11];
    ele[6][6] != ele[9][6];
    ele[6][6] != ele[9][7];
    ele[6][6] != ele[9][8];
    ele[6][6] != ele[9][9];
    ele[6][7] != ele[10][10];
    ele[6][7] != ele[10][11];
    ele[6][7] != ele[10][6];
    ele[6][7] != ele[10][7];
    ele[6][7] != ele[10][8];
    ele[6][7] != ele[10][9];
    ele[6][7] != ele[11][10];
    ele[6][7] != ele[11][11];
    ele[6][7] != ele[11][6];
    ele[6][7] != ele[11][7];
    ele[6][7] != ele[11][8];
    ele[6][7] != ele[11][9];
    ele[6][7] != ele[12][7];
    ele[6][7] != ele[13][7];
    ele[6][7] != ele[14][7];
    ele[6][7] != ele[15][7];
    ele[6][7] != ele[16][7];
    ele[6][7] != ele[17][7];
    ele[6][7] != ele[18][7];
    ele[6][7] != ele[19][7];
    ele[6][7] != ele[20][7];
    ele[6][7] != ele[21][7];
    ele[6][7] != ele[22][7];
    ele[6][7] != ele[23][7];
    ele[6][7] != ele[24][7];
    ele[6][7] != ele[25][7];
    ele[6][7] != ele[26][7];
    ele[6][7] != ele[27][7];
    ele[6][7] != ele[28][7];
    ele[6][7] != ele[29][7];
    ele[6][7] != ele[30][7];
    ele[6][7] != ele[31][7];
    ele[6][7] != ele[32][7];
    ele[6][7] != ele[33][7];
    ele[6][7] != ele[34][7];
    ele[6][7] != ele[35][7];
    ele[6][7] != ele[6][10];
    ele[6][7] != ele[6][11];
    ele[6][7] != ele[6][12];
    ele[6][7] != ele[6][13];
    ele[6][7] != ele[6][14];
    ele[6][7] != ele[6][15];
    ele[6][7] != ele[6][16];
    ele[6][7] != ele[6][17];
    ele[6][7] != ele[6][18];
    ele[6][7] != ele[6][19];
    ele[6][7] != ele[6][20];
    ele[6][7] != ele[6][21];
    ele[6][7] != ele[6][22];
    ele[6][7] != ele[6][23];
    ele[6][7] != ele[6][24];
    ele[6][7] != ele[6][25];
    ele[6][7] != ele[6][26];
    ele[6][7] != ele[6][27];
    ele[6][7] != ele[6][28];
    ele[6][7] != ele[6][29];
    ele[6][7] != ele[6][30];
    ele[6][7] != ele[6][31];
    ele[6][7] != ele[6][32];
    ele[6][7] != ele[6][33];
    ele[6][7] != ele[6][34];
    ele[6][7] != ele[6][35];
    ele[6][7] != ele[6][8];
    ele[6][7] != ele[6][9];
    ele[6][7] != ele[7][10];
    ele[6][7] != ele[7][11];
    ele[6][7] != ele[7][6];
    ele[6][7] != ele[7][7];
    ele[6][7] != ele[7][8];
    ele[6][7] != ele[7][9];
    ele[6][7] != ele[8][10];
    ele[6][7] != ele[8][11];
    ele[6][7] != ele[8][6];
    ele[6][7] != ele[8][7];
    ele[6][7] != ele[8][8];
    ele[6][7] != ele[8][9];
    ele[6][7] != ele[9][10];
    ele[6][7] != ele[9][11];
    ele[6][7] != ele[9][6];
    ele[6][7] != ele[9][7];
    ele[6][7] != ele[9][8];
    ele[6][7] != ele[9][9];
    ele[6][8] != ele[10][10];
    ele[6][8] != ele[10][11];
    ele[6][8] != ele[10][6];
    ele[6][8] != ele[10][7];
    ele[6][8] != ele[10][8];
    ele[6][8] != ele[10][9];
    ele[6][8] != ele[11][10];
    ele[6][8] != ele[11][11];
    ele[6][8] != ele[11][6];
    ele[6][8] != ele[11][7];
    ele[6][8] != ele[11][8];
    ele[6][8] != ele[11][9];
    ele[6][8] != ele[12][8];
    ele[6][8] != ele[13][8];
    ele[6][8] != ele[14][8];
    ele[6][8] != ele[15][8];
    ele[6][8] != ele[16][8];
    ele[6][8] != ele[17][8];
    ele[6][8] != ele[18][8];
    ele[6][8] != ele[19][8];
    ele[6][8] != ele[20][8];
    ele[6][8] != ele[21][8];
    ele[6][8] != ele[22][8];
    ele[6][8] != ele[23][8];
    ele[6][8] != ele[24][8];
    ele[6][8] != ele[25][8];
    ele[6][8] != ele[26][8];
    ele[6][8] != ele[27][8];
    ele[6][8] != ele[28][8];
    ele[6][8] != ele[29][8];
    ele[6][8] != ele[30][8];
    ele[6][8] != ele[31][8];
    ele[6][8] != ele[32][8];
    ele[6][8] != ele[33][8];
    ele[6][8] != ele[34][8];
    ele[6][8] != ele[35][8];
    ele[6][8] != ele[6][10];
    ele[6][8] != ele[6][11];
    ele[6][8] != ele[6][12];
    ele[6][8] != ele[6][13];
    ele[6][8] != ele[6][14];
    ele[6][8] != ele[6][15];
    ele[6][8] != ele[6][16];
    ele[6][8] != ele[6][17];
    ele[6][8] != ele[6][18];
    ele[6][8] != ele[6][19];
    ele[6][8] != ele[6][20];
    ele[6][8] != ele[6][21];
    ele[6][8] != ele[6][22];
    ele[6][8] != ele[6][23];
    ele[6][8] != ele[6][24];
    ele[6][8] != ele[6][25];
    ele[6][8] != ele[6][26];
    ele[6][8] != ele[6][27];
    ele[6][8] != ele[6][28];
    ele[6][8] != ele[6][29];
    ele[6][8] != ele[6][30];
    ele[6][8] != ele[6][31];
    ele[6][8] != ele[6][32];
    ele[6][8] != ele[6][33];
    ele[6][8] != ele[6][34];
    ele[6][8] != ele[6][35];
    ele[6][8] != ele[6][9];
    ele[6][8] != ele[7][10];
    ele[6][8] != ele[7][11];
    ele[6][8] != ele[7][6];
    ele[6][8] != ele[7][7];
    ele[6][8] != ele[7][8];
    ele[6][8] != ele[7][9];
    ele[6][8] != ele[8][10];
    ele[6][8] != ele[8][11];
    ele[6][8] != ele[8][6];
    ele[6][8] != ele[8][7];
    ele[6][8] != ele[8][8];
    ele[6][8] != ele[8][9];
    ele[6][8] != ele[9][10];
    ele[6][8] != ele[9][11];
    ele[6][8] != ele[9][6];
    ele[6][8] != ele[9][7];
    ele[6][8] != ele[9][8];
    ele[6][8] != ele[9][9];
    ele[6][9] != ele[10][10];
    ele[6][9] != ele[10][11];
    ele[6][9] != ele[10][6];
    ele[6][9] != ele[10][7];
    ele[6][9] != ele[10][8];
    ele[6][9] != ele[10][9];
    ele[6][9] != ele[11][10];
    ele[6][9] != ele[11][11];
    ele[6][9] != ele[11][6];
    ele[6][9] != ele[11][7];
    ele[6][9] != ele[11][8];
    ele[6][9] != ele[11][9];
    ele[6][9] != ele[12][9];
    ele[6][9] != ele[13][9];
    ele[6][9] != ele[14][9];
    ele[6][9] != ele[15][9];
    ele[6][9] != ele[16][9];
    ele[6][9] != ele[17][9];
    ele[6][9] != ele[18][9];
    ele[6][9] != ele[19][9];
    ele[6][9] != ele[20][9];
    ele[6][9] != ele[21][9];
    ele[6][9] != ele[22][9];
    ele[6][9] != ele[23][9];
    ele[6][9] != ele[24][9];
    ele[6][9] != ele[25][9];
    ele[6][9] != ele[26][9];
    ele[6][9] != ele[27][9];
    ele[6][9] != ele[28][9];
    ele[6][9] != ele[29][9];
    ele[6][9] != ele[30][9];
    ele[6][9] != ele[31][9];
    ele[6][9] != ele[32][9];
    ele[6][9] != ele[33][9];
    ele[6][9] != ele[34][9];
    ele[6][9] != ele[35][9];
    ele[6][9] != ele[6][10];
    ele[6][9] != ele[6][11];
    ele[6][9] != ele[6][12];
    ele[6][9] != ele[6][13];
    ele[6][9] != ele[6][14];
    ele[6][9] != ele[6][15];
    ele[6][9] != ele[6][16];
    ele[6][9] != ele[6][17];
    ele[6][9] != ele[6][18];
    ele[6][9] != ele[6][19];
    ele[6][9] != ele[6][20];
    ele[6][9] != ele[6][21];
    ele[6][9] != ele[6][22];
    ele[6][9] != ele[6][23];
    ele[6][9] != ele[6][24];
    ele[6][9] != ele[6][25];
    ele[6][9] != ele[6][26];
    ele[6][9] != ele[6][27];
    ele[6][9] != ele[6][28];
    ele[6][9] != ele[6][29];
    ele[6][9] != ele[6][30];
    ele[6][9] != ele[6][31];
    ele[6][9] != ele[6][32];
    ele[6][9] != ele[6][33];
    ele[6][9] != ele[6][34];
    ele[6][9] != ele[6][35];
    ele[6][9] != ele[7][10];
    ele[6][9] != ele[7][11];
    ele[6][9] != ele[7][6];
    ele[6][9] != ele[7][7];
    ele[6][9] != ele[7][8];
    ele[6][9] != ele[7][9];
    ele[6][9] != ele[8][10];
    ele[6][9] != ele[8][11];
    ele[6][9] != ele[8][6];
    ele[6][9] != ele[8][7];
    ele[6][9] != ele[8][8];
    ele[6][9] != ele[8][9];
    ele[6][9] != ele[9][10];
    ele[6][9] != ele[9][11];
    ele[6][9] != ele[9][6];
    ele[6][9] != ele[9][7];
    ele[6][9] != ele[9][8];
    ele[6][9] != ele[9][9];
    ele[7][0] != ele[10][0];
    ele[7][0] != ele[10][1];
    ele[7][0] != ele[10][2];
    ele[7][0] != ele[10][3];
    ele[7][0] != ele[10][4];
    ele[7][0] != ele[10][5];
    ele[7][0] != ele[11][0];
    ele[7][0] != ele[11][1];
    ele[7][0] != ele[11][2];
    ele[7][0] != ele[11][3];
    ele[7][0] != ele[11][4];
    ele[7][0] != ele[11][5];
    ele[7][0] != ele[12][0];
    ele[7][0] != ele[13][0];
    ele[7][0] != ele[14][0];
    ele[7][0] != ele[15][0];
    ele[7][0] != ele[16][0];
    ele[7][0] != ele[17][0];
    ele[7][0] != ele[18][0];
    ele[7][0] != ele[19][0];
    ele[7][0] != ele[20][0];
    ele[7][0] != ele[21][0];
    ele[7][0] != ele[22][0];
    ele[7][0] != ele[23][0];
    ele[7][0] != ele[24][0];
    ele[7][0] != ele[25][0];
    ele[7][0] != ele[26][0];
    ele[7][0] != ele[27][0];
    ele[7][0] != ele[28][0];
    ele[7][0] != ele[29][0];
    ele[7][0] != ele[30][0];
    ele[7][0] != ele[31][0];
    ele[7][0] != ele[32][0];
    ele[7][0] != ele[33][0];
    ele[7][0] != ele[34][0];
    ele[7][0] != ele[35][0];
    ele[7][0] != ele[7][1];
    ele[7][0] != ele[7][10];
    ele[7][0] != ele[7][11];
    ele[7][0] != ele[7][12];
    ele[7][0] != ele[7][13];
    ele[7][0] != ele[7][14];
    ele[7][0] != ele[7][15];
    ele[7][0] != ele[7][16];
    ele[7][0] != ele[7][17];
    ele[7][0] != ele[7][18];
    ele[7][0] != ele[7][19];
    ele[7][0] != ele[7][2];
    ele[7][0] != ele[7][20];
    ele[7][0] != ele[7][21];
    ele[7][0] != ele[7][22];
    ele[7][0] != ele[7][23];
    ele[7][0] != ele[7][24];
    ele[7][0] != ele[7][25];
    ele[7][0] != ele[7][26];
    ele[7][0] != ele[7][27];
    ele[7][0] != ele[7][28];
    ele[7][0] != ele[7][29];
    ele[7][0] != ele[7][3];
    ele[7][0] != ele[7][30];
    ele[7][0] != ele[7][31];
    ele[7][0] != ele[7][32];
    ele[7][0] != ele[7][33];
    ele[7][0] != ele[7][34];
    ele[7][0] != ele[7][35];
    ele[7][0] != ele[7][4];
    ele[7][0] != ele[7][5];
    ele[7][0] != ele[7][6];
    ele[7][0] != ele[7][7];
    ele[7][0] != ele[7][8];
    ele[7][0] != ele[7][9];
    ele[7][0] != ele[8][0];
    ele[7][0] != ele[8][1];
    ele[7][0] != ele[8][2];
    ele[7][0] != ele[8][3];
    ele[7][0] != ele[8][4];
    ele[7][0] != ele[8][5];
    ele[7][0] != ele[9][0];
    ele[7][0] != ele[9][1];
    ele[7][0] != ele[9][2];
    ele[7][0] != ele[9][3];
    ele[7][0] != ele[9][4];
    ele[7][0] != ele[9][5];
    ele[7][1] != ele[10][0];
    ele[7][1] != ele[10][1];
    ele[7][1] != ele[10][2];
    ele[7][1] != ele[10][3];
    ele[7][1] != ele[10][4];
    ele[7][1] != ele[10][5];
    ele[7][1] != ele[11][0];
    ele[7][1] != ele[11][1];
    ele[7][1] != ele[11][2];
    ele[7][1] != ele[11][3];
    ele[7][1] != ele[11][4];
    ele[7][1] != ele[11][5];
    ele[7][1] != ele[12][1];
    ele[7][1] != ele[13][1];
    ele[7][1] != ele[14][1];
    ele[7][1] != ele[15][1];
    ele[7][1] != ele[16][1];
    ele[7][1] != ele[17][1];
    ele[7][1] != ele[18][1];
    ele[7][1] != ele[19][1];
    ele[7][1] != ele[20][1];
    ele[7][1] != ele[21][1];
    ele[7][1] != ele[22][1];
    ele[7][1] != ele[23][1];
    ele[7][1] != ele[24][1];
    ele[7][1] != ele[25][1];
    ele[7][1] != ele[26][1];
    ele[7][1] != ele[27][1];
    ele[7][1] != ele[28][1];
    ele[7][1] != ele[29][1];
    ele[7][1] != ele[30][1];
    ele[7][1] != ele[31][1];
    ele[7][1] != ele[32][1];
    ele[7][1] != ele[33][1];
    ele[7][1] != ele[34][1];
    ele[7][1] != ele[35][1];
    ele[7][1] != ele[7][10];
    ele[7][1] != ele[7][11];
    ele[7][1] != ele[7][12];
    ele[7][1] != ele[7][13];
    ele[7][1] != ele[7][14];
    ele[7][1] != ele[7][15];
    ele[7][1] != ele[7][16];
    ele[7][1] != ele[7][17];
    ele[7][1] != ele[7][18];
    ele[7][1] != ele[7][19];
    ele[7][1] != ele[7][2];
    ele[7][1] != ele[7][20];
    ele[7][1] != ele[7][21];
    ele[7][1] != ele[7][22];
    ele[7][1] != ele[7][23];
    ele[7][1] != ele[7][24];
    ele[7][1] != ele[7][25];
    ele[7][1] != ele[7][26];
    ele[7][1] != ele[7][27];
    ele[7][1] != ele[7][28];
    ele[7][1] != ele[7][29];
    ele[7][1] != ele[7][3];
    ele[7][1] != ele[7][30];
    ele[7][1] != ele[7][31];
    ele[7][1] != ele[7][32];
    ele[7][1] != ele[7][33];
    ele[7][1] != ele[7][34];
    ele[7][1] != ele[7][35];
    ele[7][1] != ele[7][4];
    ele[7][1] != ele[7][5];
    ele[7][1] != ele[7][6];
    ele[7][1] != ele[7][7];
    ele[7][1] != ele[7][8];
    ele[7][1] != ele[7][9];
    ele[7][1] != ele[8][0];
    ele[7][1] != ele[8][1];
    ele[7][1] != ele[8][2];
    ele[7][1] != ele[8][3];
    ele[7][1] != ele[8][4];
    ele[7][1] != ele[8][5];
    ele[7][1] != ele[9][0];
    ele[7][1] != ele[9][1];
    ele[7][1] != ele[9][2];
    ele[7][1] != ele[9][3];
    ele[7][1] != ele[9][4];
    ele[7][1] != ele[9][5];
    ele[7][10] != ele[10][10];
    ele[7][10] != ele[10][11];
    ele[7][10] != ele[10][6];
    ele[7][10] != ele[10][7];
    ele[7][10] != ele[10][8];
    ele[7][10] != ele[10][9];
    ele[7][10] != ele[11][10];
    ele[7][10] != ele[11][11];
    ele[7][10] != ele[11][6];
    ele[7][10] != ele[11][7];
    ele[7][10] != ele[11][8];
    ele[7][10] != ele[11][9];
    ele[7][10] != ele[12][10];
    ele[7][10] != ele[13][10];
    ele[7][10] != ele[14][10];
    ele[7][10] != ele[15][10];
    ele[7][10] != ele[16][10];
    ele[7][10] != ele[17][10];
    ele[7][10] != ele[18][10];
    ele[7][10] != ele[19][10];
    ele[7][10] != ele[20][10];
    ele[7][10] != ele[21][10];
    ele[7][10] != ele[22][10];
    ele[7][10] != ele[23][10];
    ele[7][10] != ele[24][10];
    ele[7][10] != ele[25][10];
    ele[7][10] != ele[26][10];
    ele[7][10] != ele[27][10];
    ele[7][10] != ele[28][10];
    ele[7][10] != ele[29][10];
    ele[7][10] != ele[30][10];
    ele[7][10] != ele[31][10];
    ele[7][10] != ele[32][10];
    ele[7][10] != ele[33][10];
    ele[7][10] != ele[34][10];
    ele[7][10] != ele[35][10];
    ele[7][10] != ele[7][11];
    ele[7][10] != ele[7][12];
    ele[7][10] != ele[7][13];
    ele[7][10] != ele[7][14];
    ele[7][10] != ele[7][15];
    ele[7][10] != ele[7][16];
    ele[7][10] != ele[7][17];
    ele[7][10] != ele[7][18];
    ele[7][10] != ele[7][19];
    ele[7][10] != ele[7][20];
    ele[7][10] != ele[7][21];
    ele[7][10] != ele[7][22];
    ele[7][10] != ele[7][23];
    ele[7][10] != ele[7][24];
    ele[7][10] != ele[7][25];
    ele[7][10] != ele[7][26];
    ele[7][10] != ele[7][27];
    ele[7][10] != ele[7][28];
    ele[7][10] != ele[7][29];
    ele[7][10] != ele[7][30];
    ele[7][10] != ele[7][31];
    ele[7][10] != ele[7][32];
    ele[7][10] != ele[7][33];
    ele[7][10] != ele[7][34];
    ele[7][10] != ele[7][35];
    ele[7][10] != ele[8][10];
    ele[7][10] != ele[8][11];
    ele[7][10] != ele[8][6];
    ele[7][10] != ele[8][7];
    ele[7][10] != ele[8][8];
    ele[7][10] != ele[8][9];
    ele[7][10] != ele[9][10];
    ele[7][10] != ele[9][11];
    ele[7][10] != ele[9][6];
    ele[7][10] != ele[9][7];
    ele[7][10] != ele[9][8];
    ele[7][10] != ele[9][9];
    ele[7][11] != ele[10][10];
    ele[7][11] != ele[10][11];
    ele[7][11] != ele[10][6];
    ele[7][11] != ele[10][7];
    ele[7][11] != ele[10][8];
    ele[7][11] != ele[10][9];
    ele[7][11] != ele[11][10];
    ele[7][11] != ele[11][11];
    ele[7][11] != ele[11][6];
    ele[7][11] != ele[11][7];
    ele[7][11] != ele[11][8];
    ele[7][11] != ele[11][9];
    ele[7][11] != ele[12][11];
    ele[7][11] != ele[13][11];
    ele[7][11] != ele[14][11];
    ele[7][11] != ele[15][11];
    ele[7][11] != ele[16][11];
    ele[7][11] != ele[17][11];
    ele[7][11] != ele[18][11];
    ele[7][11] != ele[19][11];
    ele[7][11] != ele[20][11];
    ele[7][11] != ele[21][11];
    ele[7][11] != ele[22][11];
    ele[7][11] != ele[23][11];
    ele[7][11] != ele[24][11];
    ele[7][11] != ele[25][11];
    ele[7][11] != ele[26][11];
    ele[7][11] != ele[27][11];
    ele[7][11] != ele[28][11];
    ele[7][11] != ele[29][11];
    ele[7][11] != ele[30][11];
    ele[7][11] != ele[31][11];
    ele[7][11] != ele[32][11];
    ele[7][11] != ele[33][11];
    ele[7][11] != ele[34][11];
    ele[7][11] != ele[35][11];
    ele[7][11] != ele[7][12];
    ele[7][11] != ele[7][13];
    ele[7][11] != ele[7][14];
    ele[7][11] != ele[7][15];
    ele[7][11] != ele[7][16];
    ele[7][11] != ele[7][17];
    ele[7][11] != ele[7][18];
    ele[7][11] != ele[7][19];
    ele[7][11] != ele[7][20];
    ele[7][11] != ele[7][21];
    ele[7][11] != ele[7][22];
    ele[7][11] != ele[7][23];
    ele[7][11] != ele[7][24];
    ele[7][11] != ele[7][25];
    ele[7][11] != ele[7][26];
    ele[7][11] != ele[7][27];
    ele[7][11] != ele[7][28];
    ele[7][11] != ele[7][29];
    ele[7][11] != ele[7][30];
    ele[7][11] != ele[7][31];
    ele[7][11] != ele[7][32];
    ele[7][11] != ele[7][33];
    ele[7][11] != ele[7][34];
    ele[7][11] != ele[7][35];
    ele[7][11] != ele[8][10];
    ele[7][11] != ele[8][11];
    ele[7][11] != ele[8][6];
    ele[7][11] != ele[8][7];
    ele[7][11] != ele[8][8];
    ele[7][11] != ele[8][9];
    ele[7][11] != ele[9][10];
    ele[7][11] != ele[9][11];
    ele[7][11] != ele[9][6];
    ele[7][11] != ele[9][7];
    ele[7][11] != ele[9][8];
    ele[7][11] != ele[9][9];
    ele[7][12] != ele[10][12];
    ele[7][12] != ele[10][13];
    ele[7][12] != ele[10][14];
    ele[7][12] != ele[10][15];
    ele[7][12] != ele[10][16];
    ele[7][12] != ele[10][17];
    ele[7][12] != ele[11][12];
    ele[7][12] != ele[11][13];
    ele[7][12] != ele[11][14];
    ele[7][12] != ele[11][15];
    ele[7][12] != ele[11][16];
    ele[7][12] != ele[11][17];
    ele[7][12] != ele[12][12];
    ele[7][12] != ele[13][12];
    ele[7][12] != ele[14][12];
    ele[7][12] != ele[15][12];
    ele[7][12] != ele[16][12];
    ele[7][12] != ele[17][12];
    ele[7][12] != ele[18][12];
    ele[7][12] != ele[19][12];
    ele[7][12] != ele[20][12];
    ele[7][12] != ele[21][12];
    ele[7][12] != ele[22][12];
    ele[7][12] != ele[23][12];
    ele[7][12] != ele[24][12];
    ele[7][12] != ele[25][12];
    ele[7][12] != ele[26][12];
    ele[7][12] != ele[27][12];
    ele[7][12] != ele[28][12];
    ele[7][12] != ele[29][12];
    ele[7][12] != ele[30][12];
    ele[7][12] != ele[31][12];
    ele[7][12] != ele[32][12];
    ele[7][12] != ele[33][12];
    ele[7][12] != ele[34][12];
    ele[7][12] != ele[35][12];
    ele[7][12] != ele[7][13];
    ele[7][12] != ele[7][14];
    ele[7][12] != ele[7][15];
    ele[7][12] != ele[7][16];
    ele[7][12] != ele[7][17];
    ele[7][12] != ele[7][18];
    ele[7][12] != ele[7][19];
    ele[7][12] != ele[7][20];
    ele[7][12] != ele[7][21];
    ele[7][12] != ele[7][22];
    ele[7][12] != ele[7][23];
    ele[7][12] != ele[7][24];
    ele[7][12] != ele[7][25];
    ele[7][12] != ele[7][26];
    ele[7][12] != ele[7][27];
    ele[7][12] != ele[7][28];
    ele[7][12] != ele[7][29];
    ele[7][12] != ele[7][30];
    ele[7][12] != ele[7][31];
    ele[7][12] != ele[7][32];
    ele[7][12] != ele[7][33];
    ele[7][12] != ele[7][34];
    ele[7][12] != ele[7][35];
    ele[7][12] != ele[8][12];
    ele[7][12] != ele[8][13];
    ele[7][12] != ele[8][14];
    ele[7][12] != ele[8][15];
    ele[7][12] != ele[8][16];
    ele[7][12] != ele[8][17];
    ele[7][12] != ele[9][12];
    ele[7][12] != ele[9][13];
    ele[7][12] != ele[9][14];
    ele[7][12] != ele[9][15];
    ele[7][12] != ele[9][16];
    ele[7][12] != ele[9][17];
    ele[7][13] != ele[10][12];
    ele[7][13] != ele[10][13];
    ele[7][13] != ele[10][14];
    ele[7][13] != ele[10][15];
    ele[7][13] != ele[10][16];
    ele[7][13] != ele[10][17];
    ele[7][13] != ele[11][12];
    ele[7][13] != ele[11][13];
    ele[7][13] != ele[11][14];
    ele[7][13] != ele[11][15];
    ele[7][13] != ele[11][16];
    ele[7][13] != ele[11][17];
    ele[7][13] != ele[12][13];
    ele[7][13] != ele[13][13];
    ele[7][13] != ele[14][13];
    ele[7][13] != ele[15][13];
    ele[7][13] != ele[16][13];
    ele[7][13] != ele[17][13];
    ele[7][13] != ele[18][13];
    ele[7][13] != ele[19][13];
    ele[7][13] != ele[20][13];
    ele[7][13] != ele[21][13];
    ele[7][13] != ele[22][13];
    ele[7][13] != ele[23][13];
    ele[7][13] != ele[24][13];
    ele[7][13] != ele[25][13];
    ele[7][13] != ele[26][13];
    ele[7][13] != ele[27][13];
    ele[7][13] != ele[28][13];
    ele[7][13] != ele[29][13];
    ele[7][13] != ele[30][13];
    ele[7][13] != ele[31][13];
    ele[7][13] != ele[32][13];
    ele[7][13] != ele[33][13];
    ele[7][13] != ele[34][13];
    ele[7][13] != ele[35][13];
    ele[7][13] != ele[7][14];
    ele[7][13] != ele[7][15];
    ele[7][13] != ele[7][16];
    ele[7][13] != ele[7][17];
    ele[7][13] != ele[7][18];
    ele[7][13] != ele[7][19];
    ele[7][13] != ele[7][20];
    ele[7][13] != ele[7][21];
    ele[7][13] != ele[7][22];
    ele[7][13] != ele[7][23];
    ele[7][13] != ele[7][24];
    ele[7][13] != ele[7][25];
    ele[7][13] != ele[7][26];
    ele[7][13] != ele[7][27];
    ele[7][13] != ele[7][28];
    ele[7][13] != ele[7][29];
    ele[7][13] != ele[7][30];
    ele[7][13] != ele[7][31];
    ele[7][13] != ele[7][32];
    ele[7][13] != ele[7][33];
    ele[7][13] != ele[7][34];
    ele[7][13] != ele[7][35];
    ele[7][13] != ele[8][12];
    ele[7][13] != ele[8][13];
    ele[7][13] != ele[8][14];
    ele[7][13] != ele[8][15];
    ele[7][13] != ele[8][16];
    ele[7][13] != ele[8][17];
    ele[7][13] != ele[9][12];
    ele[7][13] != ele[9][13];
    ele[7][13] != ele[9][14];
    ele[7][13] != ele[9][15];
    ele[7][13] != ele[9][16];
    ele[7][13] != ele[9][17];
    ele[7][14] != ele[10][12];
    ele[7][14] != ele[10][13];
    ele[7][14] != ele[10][14];
    ele[7][14] != ele[10][15];
    ele[7][14] != ele[10][16];
    ele[7][14] != ele[10][17];
    ele[7][14] != ele[11][12];
    ele[7][14] != ele[11][13];
    ele[7][14] != ele[11][14];
    ele[7][14] != ele[11][15];
    ele[7][14] != ele[11][16];
    ele[7][14] != ele[11][17];
    ele[7][14] != ele[12][14];
    ele[7][14] != ele[13][14];
    ele[7][14] != ele[14][14];
    ele[7][14] != ele[15][14];
    ele[7][14] != ele[16][14];
    ele[7][14] != ele[17][14];
    ele[7][14] != ele[18][14];
    ele[7][14] != ele[19][14];
    ele[7][14] != ele[20][14];
    ele[7][14] != ele[21][14];
    ele[7][14] != ele[22][14];
    ele[7][14] != ele[23][14];
    ele[7][14] != ele[24][14];
    ele[7][14] != ele[25][14];
    ele[7][14] != ele[26][14];
    ele[7][14] != ele[27][14];
    ele[7][14] != ele[28][14];
    ele[7][14] != ele[29][14];
    ele[7][14] != ele[30][14];
    ele[7][14] != ele[31][14];
    ele[7][14] != ele[32][14];
    ele[7][14] != ele[33][14];
    ele[7][14] != ele[34][14];
    ele[7][14] != ele[35][14];
    ele[7][14] != ele[7][15];
    ele[7][14] != ele[7][16];
    ele[7][14] != ele[7][17];
    ele[7][14] != ele[7][18];
    ele[7][14] != ele[7][19];
    ele[7][14] != ele[7][20];
    ele[7][14] != ele[7][21];
    ele[7][14] != ele[7][22];
    ele[7][14] != ele[7][23];
    ele[7][14] != ele[7][24];
    ele[7][14] != ele[7][25];
    ele[7][14] != ele[7][26];
    ele[7][14] != ele[7][27];
    ele[7][14] != ele[7][28];
    ele[7][14] != ele[7][29];
    ele[7][14] != ele[7][30];
    ele[7][14] != ele[7][31];
    ele[7][14] != ele[7][32];
    ele[7][14] != ele[7][33];
    ele[7][14] != ele[7][34];
    ele[7][14] != ele[7][35];
    ele[7][14] != ele[8][12];
    ele[7][14] != ele[8][13];
    ele[7][14] != ele[8][14];
    ele[7][14] != ele[8][15];
    ele[7][14] != ele[8][16];
    ele[7][14] != ele[8][17];
    ele[7][14] != ele[9][12];
    ele[7][14] != ele[9][13];
    ele[7][14] != ele[9][14];
    ele[7][14] != ele[9][15];
    ele[7][14] != ele[9][16];
    ele[7][14] != ele[9][17];
    ele[7][15] != ele[10][12];
    ele[7][15] != ele[10][13];
    ele[7][15] != ele[10][14];
    ele[7][15] != ele[10][15];
    ele[7][15] != ele[10][16];
    ele[7][15] != ele[10][17];
    ele[7][15] != ele[11][12];
    ele[7][15] != ele[11][13];
    ele[7][15] != ele[11][14];
    ele[7][15] != ele[11][15];
    ele[7][15] != ele[11][16];
    ele[7][15] != ele[11][17];
    ele[7][15] != ele[12][15];
    ele[7][15] != ele[13][15];
    ele[7][15] != ele[14][15];
    ele[7][15] != ele[15][15];
    ele[7][15] != ele[16][15];
    ele[7][15] != ele[17][15];
    ele[7][15] != ele[18][15];
    ele[7][15] != ele[19][15];
    ele[7][15] != ele[20][15];
    ele[7][15] != ele[21][15];
    ele[7][15] != ele[22][15];
    ele[7][15] != ele[23][15];
    ele[7][15] != ele[24][15];
    ele[7][15] != ele[25][15];
    ele[7][15] != ele[26][15];
    ele[7][15] != ele[27][15];
    ele[7][15] != ele[28][15];
    ele[7][15] != ele[29][15];
    ele[7][15] != ele[30][15];
    ele[7][15] != ele[31][15];
    ele[7][15] != ele[32][15];
    ele[7][15] != ele[33][15];
    ele[7][15] != ele[34][15];
    ele[7][15] != ele[35][15];
    ele[7][15] != ele[7][16];
    ele[7][15] != ele[7][17];
    ele[7][15] != ele[7][18];
    ele[7][15] != ele[7][19];
    ele[7][15] != ele[7][20];
    ele[7][15] != ele[7][21];
    ele[7][15] != ele[7][22];
    ele[7][15] != ele[7][23];
    ele[7][15] != ele[7][24];
    ele[7][15] != ele[7][25];
    ele[7][15] != ele[7][26];
    ele[7][15] != ele[7][27];
    ele[7][15] != ele[7][28];
    ele[7][15] != ele[7][29];
    ele[7][15] != ele[7][30];
    ele[7][15] != ele[7][31];
    ele[7][15] != ele[7][32];
    ele[7][15] != ele[7][33];
    ele[7][15] != ele[7][34];
    ele[7][15] != ele[7][35];
    ele[7][15] != ele[8][12];
    ele[7][15] != ele[8][13];
    ele[7][15] != ele[8][14];
    ele[7][15] != ele[8][15];
    ele[7][15] != ele[8][16];
    ele[7][15] != ele[8][17];
    ele[7][15] != ele[9][12];
    ele[7][15] != ele[9][13];
    ele[7][15] != ele[9][14];
    ele[7][15] != ele[9][15];
    ele[7][15] != ele[9][16];
    ele[7][15] != ele[9][17];
    ele[7][16] != ele[10][12];
    ele[7][16] != ele[10][13];
    ele[7][16] != ele[10][14];
    ele[7][16] != ele[10][15];
    ele[7][16] != ele[10][16];
    ele[7][16] != ele[10][17];
    ele[7][16] != ele[11][12];
    ele[7][16] != ele[11][13];
    ele[7][16] != ele[11][14];
    ele[7][16] != ele[11][15];
    ele[7][16] != ele[11][16];
    ele[7][16] != ele[11][17];
    ele[7][16] != ele[12][16];
    ele[7][16] != ele[13][16];
    ele[7][16] != ele[14][16];
    ele[7][16] != ele[15][16];
    ele[7][16] != ele[16][16];
    ele[7][16] != ele[17][16];
    ele[7][16] != ele[18][16];
    ele[7][16] != ele[19][16];
    ele[7][16] != ele[20][16];
    ele[7][16] != ele[21][16];
    ele[7][16] != ele[22][16];
    ele[7][16] != ele[23][16];
    ele[7][16] != ele[24][16];
    ele[7][16] != ele[25][16];
    ele[7][16] != ele[26][16];
    ele[7][16] != ele[27][16];
    ele[7][16] != ele[28][16];
    ele[7][16] != ele[29][16];
    ele[7][16] != ele[30][16];
    ele[7][16] != ele[31][16];
    ele[7][16] != ele[32][16];
    ele[7][16] != ele[33][16];
    ele[7][16] != ele[34][16];
    ele[7][16] != ele[35][16];
    ele[7][16] != ele[7][17];
    ele[7][16] != ele[7][18];
    ele[7][16] != ele[7][19];
    ele[7][16] != ele[7][20];
    ele[7][16] != ele[7][21];
    ele[7][16] != ele[7][22];
    ele[7][16] != ele[7][23];
    ele[7][16] != ele[7][24];
    ele[7][16] != ele[7][25];
    ele[7][16] != ele[7][26];
    ele[7][16] != ele[7][27];
    ele[7][16] != ele[7][28];
    ele[7][16] != ele[7][29];
    ele[7][16] != ele[7][30];
    ele[7][16] != ele[7][31];
    ele[7][16] != ele[7][32];
    ele[7][16] != ele[7][33];
    ele[7][16] != ele[7][34];
    ele[7][16] != ele[7][35];
    ele[7][16] != ele[8][12];
    ele[7][16] != ele[8][13];
    ele[7][16] != ele[8][14];
    ele[7][16] != ele[8][15];
    ele[7][16] != ele[8][16];
    ele[7][16] != ele[8][17];
    ele[7][16] != ele[9][12];
    ele[7][16] != ele[9][13];
    ele[7][16] != ele[9][14];
    ele[7][16] != ele[9][15];
    ele[7][16] != ele[9][16];
    ele[7][16] != ele[9][17];
    ele[7][17] != ele[10][12];
    ele[7][17] != ele[10][13];
    ele[7][17] != ele[10][14];
    ele[7][17] != ele[10][15];
    ele[7][17] != ele[10][16];
    ele[7][17] != ele[10][17];
    ele[7][17] != ele[11][12];
    ele[7][17] != ele[11][13];
    ele[7][17] != ele[11][14];
    ele[7][17] != ele[11][15];
    ele[7][17] != ele[11][16];
    ele[7][17] != ele[11][17];
    ele[7][17] != ele[12][17];
    ele[7][17] != ele[13][17];
    ele[7][17] != ele[14][17];
    ele[7][17] != ele[15][17];
    ele[7][17] != ele[16][17];
    ele[7][17] != ele[17][17];
    ele[7][17] != ele[18][17];
    ele[7][17] != ele[19][17];
    ele[7][17] != ele[20][17];
    ele[7][17] != ele[21][17];
    ele[7][17] != ele[22][17];
    ele[7][17] != ele[23][17];
    ele[7][17] != ele[24][17];
    ele[7][17] != ele[25][17];
    ele[7][17] != ele[26][17];
    ele[7][17] != ele[27][17];
    ele[7][17] != ele[28][17];
    ele[7][17] != ele[29][17];
    ele[7][17] != ele[30][17];
    ele[7][17] != ele[31][17];
    ele[7][17] != ele[32][17];
    ele[7][17] != ele[33][17];
    ele[7][17] != ele[34][17];
    ele[7][17] != ele[35][17];
    ele[7][17] != ele[7][18];
    ele[7][17] != ele[7][19];
    ele[7][17] != ele[7][20];
    ele[7][17] != ele[7][21];
    ele[7][17] != ele[7][22];
    ele[7][17] != ele[7][23];
    ele[7][17] != ele[7][24];
    ele[7][17] != ele[7][25];
    ele[7][17] != ele[7][26];
    ele[7][17] != ele[7][27];
    ele[7][17] != ele[7][28];
    ele[7][17] != ele[7][29];
    ele[7][17] != ele[7][30];
    ele[7][17] != ele[7][31];
    ele[7][17] != ele[7][32];
    ele[7][17] != ele[7][33];
    ele[7][17] != ele[7][34];
    ele[7][17] != ele[7][35];
    ele[7][17] != ele[8][12];
    ele[7][17] != ele[8][13];
    ele[7][17] != ele[8][14];
    ele[7][17] != ele[8][15];
    ele[7][17] != ele[8][16];
    ele[7][17] != ele[8][17];
    ele[7][17] != ele[9][12];
    ele[7][17] != ele[9][13];
    ele[7][17] != ele[9][14];
    ele[7][17] != ele[9][15];
    ele[7][17] != ele[9][16];
    ele[7][17] != ele[9][17];
    ele[7][18] != ele[10][18];
    ele[7][18] != ele[10][19];
    ele[7][18] != ele[10][20];
    ele[7][18] != ele[10][21];
    ele[7][18] != ele[10][22];
    ele[7][18] != ele[10][23];
    ele[7][18] != ele[11][18];
    ele[7][18] != ele[11][19];
    ele[7][18] != ele[11][20];
    ele[7][18] != ele[11][21];
    ele[7][18] != ele[11][22];
    ele[7][18] != ele[11][23];
    ele[7][18] != ele[12][18];
    ele[7][18] != ele[13][18];
    ele[7][18] != ele[14][18];
    ele[7][18] != ele[15][18];
    ele[7][18] != ele[16][18];
    ele[7][18] != ele[17][18];
    ele[7][18] != ele[18][18];
    ele[7][18] != ele[19][18];
    ele[7][18] != ele[20][18];
    ele[7][18] != ele[21][18];
    ele[7][18] != ele[22][18];
    ele[7][18] != ele[23][18];
    ele[7][18] != ele[24][18];
    ele[7][18] != ele[25][18];
    ele[7][18] != ele[26][18];
    ele[7][18] != ele[27][18];
    ele[7][18] != ele[28][18];
    ele[7][18] != ele[29][18];
    ele[7][18] != ele[30][18];
    ele[7][18] != ele[31][18];
    ele[7][18] != ele[32][18];
    ele[7][18] != ele[33][18];
    ele[7][18] != ele[34][18];
    ele[7][18] != ele[35][18];
    ele[7][18] != ele[7][19];
    ele[7][18] != ele[7][20];
    ele[7][18] != ele[7][21];
    ele[7][18] != ele[7][22];
    ele[7][18] != ele[7][23];
    ele[7][18] != ele[7][24];
    ele[7][18] != ele[7][25];
    ele[7][18] != ele[7][26];
    ele[7][18] != ele[7][27];
    ele[7][18] != ele[7][28];
    ele[7][18] != ele[7][29];
    ele[7][18] != ele[7][30];
    ele[7][18] != ele[7][31];
    ele[7][18] != ele[7][32];
    ele[7][18] != ele[7][33];
    ele[7][18] != ele[7][34];
    ele[7][18] != ele[7][35];
    ele[7][18] != ele[8][18];
    ele[7][18] != ele[8][19];
    ele[7][18] != ele[8][20];
    ele[7][18] != ele[8][21];
    ele[7][18] != ele[8][22];
    ele[7][18] != ele[8][23];
    ele[7][18] != ele[9][18];
    ele[7][18] != ele[9][19];
    ele[7][18] != ele[9][20];
    ele[7][18] != ele[9][21];
    ele[7][18] != ele[9][22];
    ele[7][18] != ele[9][23];
    ele[7][19] != ele[10][18];
    ele[7][19] != ele[10][19];
    ele[7][19] != ele[10][20];
    ele[7][19] != ele[10][21];
    ele[7][19] != ele[10][22];
    ele[7][19] != ele[10][23];
    ele[7][19] != ele[11][18];
    ele[7][19] != ele[11][19];
    ele[7][19] != ele[11][20];
    ele[7][19] != ele[11][21];
    ele[7][19] != ele[11][22];
    ele[7][19] != ele[11][23];
    ele[7][19] != ele[12][19];
    ele[7][19] != ele[13][19];
    ele[7][19] != ele[14][19];
    ele[7][19] != ele[15][19];
    ele[7][19] != ele[16][19];
    ele[7][19] != ele[17][19];
    ele[7][19] != ele[18][19];
    ele[7][19] != ele[19][19];
    ele[7][19] != ele[20][19];
    ele[7][19] != ele[21][19];
    ele[7][19] != ele[22][19];
    ele[7][19] != ele[23][19];
    ele[7][19] != ele[24][19];
    ele[7][19] != ele[25][19];
    ele[7][19] != ele[26][19];
    ele[7][19] != ele[27][19];
    ele[7][19] != ele[28][19];
    ele[7][19] != ele[29][19];
    ele[7][19] != ele[30][19];
    ele[7][19] != ele[31][19];
    ele[7][19] != ele[32][19];
    ele[7][19] != ele[33][19];
    ele[7][19] != ele[34][19];
    ele[7][19] != ele[35][19];
    ele[7][19] != ele[7][20];
    ele[7][19] != ele[7][21];
    ele[7][19] != ele[7][22];
    ele[7][19] != ele[7][23];
    ele[7][19] != ele[7][24];
    ele[7][19] != ele[7][25];
    ele[7][19] != ele[7][26];
    ele[7][19] != ele[7][27];
    ele[7][19] != ele[7][28];
    ele[7][19] != ele[7][29];
    ele[7][19] != ele[7][30];
    ele[7][19] != ele[7][31];
    ele[7][19] != ele[7][32];
    ele[7][19] != ele[7][33];
    ele[7][19] != ele[7][34];
    ele[7][19] != ele[7][35];
    ele[7][19] != ele[8][18];
    ele[7][19] != ele[8][19];
    ele[7][19] != ele[8][20];
    ele[7][19] != ele[8][21];
    ele[7][19] != ele[8][22];
    ele[7][19] != ele[8][23];
    ele[7][19] != ele[9][18];
    ele[7][19] != ele[9][19];
    ele[7][19] != ele[9][20];
    ele[7][19] != ele[9][21];
    ele[7][19] != ele[9][22];
    ele[7][19] != ele[9][23];
    ele[7][2] != ele[10][0];
    ele[7][2] != ele[10][1];
    ele[7][2] != ele[10][2];
    ele[7][2] != ele[10][3];
    ele[7][2] != ele[10][4];
    ele[7][2] != ele[10][5];
    ele[7][2] != ele[11][0];
    ele[7][2] != ele[11][1];
    ele[7][2] != ele[11][2];
    ele[7][2] != ele[11][3];
    ele[7][2] != ele[11][4];
    ele[7][2] != ele[11][5];
    ele[7][2] != ele[12][2];
    ele[7][2] != ele[13][2];
    ele[7][2] != ele[14][2];
    ele[7][2] != ele[15][2];
    ele[7][2] != ele[16][2];
    ele[7][2] != ele[17][2];
    ele[7][2] != ele[18][2];
    ele[7][2] != ele[19][2];
    ele[7][2] != ele[20][2];
    ele[7][2] != ele[21][2];
    ele[7][2] != ele[22][2];
    ele[7][2] != ele[23][2];
    ele[7][2] != ele[24][2];
    ele[7][2] != ele[25][2];
    ele[7][2] != ele[26][2];
    ele[7][2] != ele[27][2];
    ele[7][2] != ele[28][2];
    ele[7][2] != ele[29][2];
    ele[7][2] != ele[30][2];
    ele[7][2] != ele[31][2];
    ele[7][2] != ele[32][2];
    ele[7][2] != ele[33][2];
    ele[7][2] != ele[34][2];
    ele[7][2] != ele[35][2];
    ele[7][2] != ele[7][10];
    ele[7][2] != ele[7][11];
    ele[7][2] != ele[7][12];
    ele[7][2] != ele[7][13];
    ele[7][2] != ele[7][14];
    ele[7][2] != ele[7][15];
    ele[7][2] != ele[7][16];
    ele[7][2] != ele[7][17];
    ele[7][2] != ele[7][18];
    ele[7][2] != ele[7][19];
    ele[7][2] != ele[7][20];
    ele[7][2] != ele[7][21];
    ele[7][2] != ele[7][22];
    ele[7][2] != ele[7][23];
    ele[7][2] != ele[7][24];
    ele[7][2] != ele[7][25];
    ele[7][2] != ele[7][26];
    ele[7][2] != ele[7][27];
    ele[7][2] != ele[7][28];
    ele[7][2] != ele[7][29];
    ele[7][2] != ele[7][3];
    ele[7][2] != ele[7][30];
    ele[7][2] != ele[7][31];
    ele[7][2] != ele[7][32];
    ele[7][2] != ele[7][33];
    ele[7][2] != ele[7][34];
    ele[7][2] != ele[7][35];
    ele[7][2] != ele[7][4];
    ele[7][2] != ele[7][5];
    ele[7][2] != ele[7][6];
    ele[7][2] != ele[7][7];
    ele[7][2] != ele[7][8];
    ele[7][2] != ele[7][9];
    ele[7][2] != ele[8][0];
    ele[7][2] != ele[8][1];
    ele[7][2] != ele[8][2];
    ele[7][2] != ele[8][3];
    ele[7][2] != ele[8][4];
    ele[7][2] != ele[8][5];
    ele[7][2] != ele[9][0];
    ele[7][2] != ele[9][1];
    ele[7][2] != ele[9][2];
    ele[7][2] != ele[9][3];
    ele[7][2] != ele[9][4];
    ele[7][2] != ele[9][5];
    ele[7][20] != ele[10][18];
    ele[7][20] != ele[10][19];
    ele[7][20] != ele[10][20];
    ele[7][20] != ele[10][21];
    ele[7][20] != ele[10][22];
    ele[7][20] != ele[10][23];
    ele[7][20] != ele[11][18];
    ele[7][20] != ele[11][19];
    ele[7][20] != ele[11][20];
    ele[7][20] != ele[11][21];
    ele[7][20] != ele[11][22];
    ele[7][20] != ele[11][23];
    ele[7][20] != ele[12][20];
    ele[7][20] != ele[13][20];
    ele[7][20] != ele[14][20];
    ele[7][20] != ele[15][20];
    ele[7][20] != ele[16][20];
    ele[7][20] != ele[17][20];
    ele[7][20] != ele[18][20];
    ele[7][20] != ele[19][20];
    ele[7][20] != ele[20][20];
    ele[7][20] != ele[21][20];
    ele[7][20] != ele[22][20];
    ele[7][20] != ele[23][20];
    ele[7][20] != ele[24][20];
    ele[7][20] != ele[25][20];
    ele[7][20] != ele[26][20];
    ele[7][20] != ele[27][20];
    ele[7][20] != ele[28][20];
    ele[7][20] != ele[29][20];
    ele[7][20] != ele[30][20];
    ele[7][20] != ele[31][20];
    ele[7][20] != ele[32][20];
    ele[7][20] != ele[33][20];
    ele[7][20] != ele[34][20];
    ele[7][20] != ele[35][20];
    ele[7][20] != ele[7][21];
    ele[7][20] != ele[7][22];
    ele[7][20] != ele[7][23];
    ele[7][20] != ele[7][24];
    ele[7][20] != ele[7][25];
    ele[7][20] != ele[7][26];
    ele[7][20] != ele[7][27];
    ele[7][20] != ele[7][28];
    ele[7][20] != ele[7][29];
    ele[7][20] != ele[7][30];
    ele[7][20] != ele[7][31];
    ele[7][20] != ele[7][32];
    ele[7][20] != ele[7][33];
    ele[7][20] != ele[7][34];
    ele[7][20] != ele[7][35];
    ele[7][20] != ele[8][18];
    ele[7][20] != ele[8][19];
    ele[7][20] != ele[8][20];
    ele[7][20] != ele[8][21];
    ele[7][20] != ele[8][22];
    ele[7][20] != ele[8][23];
    ele[7][20] != ele[9][18];
    ele[7][20] != ele[9][19];
    ele[7][20] != ele[9][20];
    ele[7][20] != ele[9][21];
    ele[7][20] != ele[9][22];
    ele[7][20] != ele[9][23];
    ele[7][21] != ele[10][18];
    ele[7][21] != ele[10][19];
    ele[7][21] != ele[10][20];
    ele[7][21] != ele[10][21];
    ele[7][21] != ele[10][22];
    ele[7][21] != ele[10][23];
    ele[7][21] != ele[11][18];
    ele[7][21] != ele[11][19];
    ele[7][21] != ele[11][20];
    ele[7][21] != ele[11][21];
    ele[7][21] != ele[11][22];
    ele[7][21] != ele[11][23];
    ele[7][21] != ele[12][21];
    ele[7][21] != ele[13][21];
    ele[7][21] != ele[14][21];
    ele[7][21] != ele[15][21];
    ele[7][21] != ele[16][21];
    ele[7][21] != ele[17][21];
    ele[7][21] != ele[18][21];
    ele[7][21] != ele[19][21];
    ele[7][21] != ele[20][21];
    ele[7][21] != ele[21][21];
    ele[7][21] != ele[22][21];
    ele[7][21] != ele[23][21];
    ele[7][21] != ele[24][21];
    ele[7][21] != ele[25][21];
    ele[7][21] != ele[26][21];
    ele[7][21] != ele[27][21];
    ele[7][21] != ele[28][21];
    ele[7][21] != ele[29][21];
    ele[7][21] != ele[30][21];
    ele[7][21] != ele[31][21];
    ele[7][21] != ele[32][21];
    ele[7][21] != ele[33][21];
    ele[7][21] != ele[34][21];
    ele[7][21] != ele[35][21];
    ele[7][21] != ele[7][22];
    ele[7][21] != ele[7][23];
    ele[7][21] != ele[7][24];
    ele[7][21] != ele[7][25];
    ele[7][21] != ele[7][26];
    ele[7][21] != ele[7][27];
    ele[7][21] != ele[7][28];
    ele[7][21] != ele[7][29];
    ele[7][21] != ele[7][30];
    ele[7][21] != ele[7][31];
    ele[7][21] != ele[7][32];
    ele[7][21] != ele[7][33];
    ele[7][21] != ele[7][34];
    ele[7][21] != ele[7][35];
    ele[7][21] != ele[8][18];
    ele[7][21] != ele[8][19];
    ele[7][21] != ele[8][20];
    ele[7][21] != ele[8][21];
    ele[7][21] != ele[8][22];
    ele[7][21] != ele[8][23];
    ele[7][21] != ele[9][18];
    ele[7][21] != ele[9][19];
    ele[7][21] != ele[9][20];
    ele[7][21] != ele[9][21];
    ele[7][21] != ele[9][22];
    ele[7][21] != ele[9][23];
    ele[7][22] != ele[10][18];
    ele[7][22] != ele[10][19];
    ele[7][22] != ele[10][20];
    ele[7][22] != ele[10][21];
    ele[7][22] != ele[10][22];
    ele[7][22] != ele[10][23];
    ele[7][22] != ele[11][18];
    ele[7][22] != ele[11][19];
    ele[7][22] != ele[11][20];
    ele[7][22] != ele[11][21];
    ele[7][22] != ele[11][22];
    ele[7][22] != ele[11][23];
    ele[7][22] != ele[12][22];
    ele[7][22] != ele[13][22];
    ele[7][22] != ele[14][22];
    ele[7][22] != ele[15][22];
    ele[7][22] != ele[16][22];
    ele[7][22] != ele[17][22];
    ele[7][22] != ele[18][22];
    ele[7][22] != ele[19][22];
    ele[7][22] != ele[20][22];
    ele[7][22] != ele[21][22];
    ele[7][22] != ele[22][22];
    ele[7][22] != ele[23][22];
    ele[7][22] != ele[24][22];
    ele[7][22] != ele[25][22];
    ele[7][22] != ele[26][22];
    ele[7][22] != ele[27][22];
    ele[7][22] != ele[28][22];
    ele[7][22] != ele[29][22];
    ele[7][22] != ele[30][22];
    ele[7][22] != ele[31][22];
    ele[7][22] != ele[32][22];
    ele[7][22] != ele[33][22];
    ele[7][22] != ele[34][22];
    ele[7][22] != ele[35][22];
    ele[7][22] != ele[7][23];
    ele[7][22] != ele[7][24];
    ele[7][22] != ele[7][25];
    ele[7][22] != ele[7][26];
    ele[7][22] != ele[7][27];
    ele[7][22] != ele[7][28];
    ele[7][22] != ele[7][29];
    ele[7][22] != ele[7][30];
    ele[7][22] != ele[7][31];
    ele[7][22] != ele[7][32];
    ele[7][22] != ele[7][33];
    ele[7][22] != ele[7][34];
    ele[7][22] != ele[7][35];
    ele[7][22] != ele[8][18];
    ele[7][22] != ele[8][19];
    ele[7][22] != ele[8][20];
    ele[7][22] != ele[8][21];
    ele[7][22] != ele[8][22];
    ele[7][22] != ele[8][23];
    ele[7][22] != ele[9][18];
    ele[7][22] != ele[9][19];
    ele[7][22] != ele[9][20];
    ele[7][22] != ele[9][21];
    ele[7][22] != ele[9][22];
    ele[7][22] != ele[9][23];
    ele[7][23] != ele[10][18];
    ele[7][23] != ele[10][19];
    ele[7][23] != ele[10][20];
    ele[7][23] != ele[10][21];
    ele[7][23] != ele[10][22];
    ele[7][23] != ele[10][23];
    ele[7][23] != ele[11][18];
    ele[7][23] != ele[11][19];
    ele[7][23] != ele[11][20];
    ele[7][23] != ele[11][21];
    ele[7][23] != ele[11][22];
    ele[7][23] != ele[11][23];
    ele[7][23] != ele[12][23];
    ele[7][23] != ele[13][23];
    ele[7][23] != ele[14][23];
    ele[7][23] != ele[15][23];
    ele[7][23] != ele[16][23];
    ele[7][23] != ele[17][23];
    ele[7][23] != ele[18][23];
    ele[7][23] != ele[19][23];
    ele[7][23] != ele[20][23];
    ele[7][23] != ele[21][23];
    ele[7][23] != ele[22][23];
    ele[7][23] != ele[23][23];
    ele[7][23] != ele[24][23];
    ele[7][23] != ele[25][23];
    ele[7][23] != ele[26][23];
    ele[7][23] != ele[27][23];
    ele[7][23] != ele[28][23];
    ele[7][23] != ele[29][23];
    ele[7][23] != ele[30][23];
    ele[7][23] != ele[31][23];
    ele[7][23] != ele[32][23];
    ele[7][23] != ele[33][23];
    ele[7][23] != ele[34][23];
    ele[7][23] != ele[35][23];
    ele[7][23] != ele[7][24];
    ele[7][23] != ele[7][25];
    ele[7][23] != ele[7][26];
    ele[7][23] != ele[7][27];
    ele[7][23] != ele[7][28];
    ele[7][23] != ele[7][29];
    ele[7][23] != ele[7][30];
    ele[7][23] != ele[7][31];
    ele[7][23] != ele[7][32];
    ele[7][23] != ele[7][33];
    ele[7][23] != ele[7][34];
    ele[7][23] != ele[7][35];
    ele[7][23] != ele[8][18];
    ele[7][23] != ele[8][19];
    ele[7][23] != ele[8][20];
    ele[7][23] != ele[8][21];
    ele[7][23] != ele[8][22];
    ele[7][23] != ele[8][23];
    ele[7][23] != ele[9][18];
    ele[7][23] != ele[9][19];
    ele[7][23] != ele[9][20];
    ele[7][23] != ele[9][21];
    ele[7][23] != ele[9][22];
    ele[7][23] != ele[9][23];
    ele[7][24] != ele[10][24];
    ele[7][24] != ele[10][25];
    ele[7][24] != ele[10][26];
    ele[7][24] != ele[10][27];
    ele[7][24] != ele[10][28];
    ele[7][24] != ele[10][29];
    ele[7][24] != ele[11][24];
    ele[7][24] != ele[11][25];
    ele[7][24] != ele[11][26];
    ele[7][24] != ele[11][27];
    ele[7][24] != ele[11][28];
    ele[7][24] != ele[11][29];
    ele[7][24] != ele[12][24];
    ele[7][24] != ele[13][24];
    ele[7][24] != ele[14][24];
    ele[7][24] != ele[15][24];
    ele[7][24] != ele[16][24];
    ele[7][24] != ele[17][24];
    ele[7][24] != ele[18][24];
    ele[7][24] != ele[19][24];
    ele[7][24] != ele[20][24];
    ele[7][24] != ele[21][24];
    ele[7][24] != ele[22][24];
    ele[7][24] != ele[23][24];
    ele[7][24] != ele[24][24];
    ele[7][24] != ele[25][24];
    ele[7][24] != ele[26][24];
    ele[7][24] != ele[27][24];
    ele[7][24] != ele[28][24];
    ele[7][24] != ele[29][24];
    ele[7][24] != ele[30][24];
    ele[7][24] != ele[31][24];
    ele[7][24] != ele[32][24];
    ele[7][24] != ele[33][24];
    ele[7][24] != ele[34][24];
    ele[7][24] != ele[35][24];
    ele[7][24] != ele[7][25];
    ele[7][24] != ele[7][26];
    ele[7][24] != ele[7][27];
    ele[7][24] != ele[7][28];
    ele[7][24] != ele[7][29];
    ele[7][24] != ele[7][30];
    ele[7][24] != ele[7][31];
    ele[7][24] != ele[7][32];
    ele[7][24] != ele[7][33];
    ele[7][24] != ele[7][34];
    ele[7][24] != ele[7][35];
    ele[7][24] != ele[8][24];
    ele[7][24] != ele[8][25];
    ele[7][24] != ele[8][26];
    ele[7][24] != ele[8][27];
    ele[7][24] != ele[8][28];
    ele[7][24] != ele[8][29];
    ele[7][24] != ele[9][24];
    ele[7][24] != ele[9][25];
    ele[7][24] != ele[9][26];
    ele[7][24] != ele[9][27];
    ele[7][24] != ele[9][28];
    ele[7][24] != ele[9][29];
    ele[7][25] != ele[10][24];
    ele[7][25] != ele[10][25];
    ele[7][25] != ele[10][26];
    ele[7][25] != ele[10][27];
    ele[7][25] != ele[10][28];
    ele[7][25] != ele[10][29];
    ele[7][25] != ele[11][24];
    ele[7][25] != ele[11][25];
    ele[7][25] != ele[11][26];
    ele[7][25] != ele[11][27];
    ele[7][25] != ele[11][28];
    ele[7][25] != ele[11][29];
    ele[7][25] != ele[12][25];
    ele[7][25] != ele[13][25];
    ele[7][25] != ele[14][25];
    ele[7][25] != ele[15][25];
    ele[7][25] != ele[16][25];
    ele[7][25] != ele[17][25];
    ele[7][25] != ele[18][25];
    ele[7][25] != ele[19][25];
    ele[7][25] != ele[20][25];
    ele[7][25] != ele[21][25];
    ele[7][25] != ele[22][25];
    ele[7][25] != ele[23][25];
    ele[7][25] != ele[24][25];
    ele[7][25] != ele[25][25];
    ele[7][25] != ele[26][25];
    ele[7][25] != ele[27][25];
    ele[7][25] != ele[28][25];
    ele[7][25] != ele[29][25];
    ele[7][25] != ele[30][25];
    ele[7][25] != ele[31][25];
    ele[7][25] != ele[32][25];
    ele[7][25] != ele[33][25];
    ele[7][25] != ele[34][25];
    ele[7][25] != ele[35][25];
    ele[7][25] != ele[7][26];
    ele[7][25] != ele[7][27];
    ele[7][25] != ele[7][28];
    ele[7][25] != ele[7][29];
    ele[7][25] != ele[7][30];
    ele[7][25] != ele[7][31];
    ele[7][25] != ele[7][32];
    ele[7][25] != ele[7][33];
    ele[7][25] != ele[7][34];
    ele[7][25] != ele[7][35];
    ele[7][25] != ele[8][24];
    ele[7][25] != ele[8][25];
    ele[7][25] != ele[8][26];
    ele[7][25] != ele[8][27];
    ele[7][25] != ele[8][28];
    ele[7][25] != ele[8][29];
    ele[7][25] != ele[9][24];
    ele[7][25] != ele[9][25];
    ele[7][25] != ele[9][26];
    ele[7][25] != ele[9][27];
    ele[7][25] != ele[9][28];
    ele[7][25] != ele[9][29];
    ele[7][26] != ele[10][24];
    ele[7][26] != ele[10][25];
    ele[7][26] != ele[10][26];
    ele[7][26] != ele[10][27];
    ele[7][26] != ele[10][28];
    ele[7][26] != ele[10][29];
    ele[7][26] != ele[11][24];
    ele[7][26] != ele[11][25];
    ele[7][26] != ele[11][26];
    ele[7][26] != ele[11][27];
    ele[7][26] != ele[11][28];
    ele[7][26] != ele[11][29];
    ele[7][26] != ele[12][26];
    ele[7][26] != ele[13][26];
    ele[7][26] != ele[14][26];
    ele[7][26] != ele[15][26];
    ele[7][26] != ele[16][26];
    ele[7][26] != ele[17][26];
    ele[7][26] != ele[18][26];
    ele[7][26] != ele[19][26];
    ele[7][26] != ele[20][26];
    ele[7][26] != ele[21][26];
    ele[7][26] != ele[22][26];
    ele[7][26] != ele[23][26];
    ele[7][26] != ele[24][26];
    ele[7][26] != ele[25][26];
    ele[7][26] != ele[26][26];
    ele[7][26] != ele[27][26];
    ele[7][26] != ele[28][26];
    ele[7][26] != ele[29][26];
    ele[7][26] != ele[30][26];
    ele[7][26] != ele[31][26];
    ele[7][26] != ele[32][26];
    ele[7][26] != ele[33][26];
    ele[7][26] != ele[34][26];
    ele[7][26] != ele[35][26];
    ele[7][26] != ele[7][27];
    ele[7][26] != ele[7][28];
    ele[7][26] != ele[7][29];
    ele[7][26] != ele[7][30];
    ele[7][26] != ele[7][31];
    ele[7][26] != ele[7][32];
    ele[7][26] != ele[7][33];
    ele[7][26] != ele[7][34];
    ele[7][26] != ele[7][35];
    ele[7][26] != ele[8][24];
    ele[7][26] != ele[8][25];
    ele[7][26] != ele[8][26];
    ele[7][26] != ele[8][27];
    ele[7][26] != ele[8][28];
    ele[7][26] != ele[8][29];
    ele[7][26] != ele[9][24];
    ele[7][26] != ele[9][25];
    ele[7][26] != ele[9][26];
    ele[7][26] != ele[9][27];
    ele[7][26] != ele[9][28];
    ele[7][26] != ele[9][29];
    ele[7][27] != ele[10][24];
    ele[7][27] != ele[10][25];
    ele[7][27] != ele[10][26];
    ele[7][27] != ele[10][27];
    ele[7][27] != ele[10][28];
    ele[7][27] != ele[10][29];
    ele[7][27] != ele[11][24];
    ele[7][27] != ele[11][25];
    ele[7][27] != ele[11][26];
    ele[7][27] != ele[11][27];
    ele[7][27] != ele[11][28];
    ele[7][27] != ele[11][29];
    ele[7][27] != ele[12][27];
    ele[7][27] != ele[13][27];
    ele[7][27] != ele[14][27];
    ele[7][27] != ele[15][27];
    ele[7][27] != ele[16][27];
    ele[7][27] != ele[17][27];
    ele[7][27] != ele[18][27];
    ele[7][27] != ele[19][27];
    ele[7][27] != ele[20][27];
    ele[7][27] != ele[21][27];
    ele[7][27] != ele[22][27];
    ele[7][27] != ele[23][27];
    ele[7][27] != ele[24][27];
    ele[7][27] != ele[25][27];
    ele[7][27] != ele[26][27];
    ele[7][27] != ele[27][27];
    ele[7][27] != ele[28][27];
    ele[7][27] != ele[29][27];
    ele[7][27] != ele[30][27];
    ele[7][27] != ele[31][27];
    ele[7][27] != ele[32][27];
    ele[7][27] != ele[33][27];
    ele[7][27] != ele[34][27];
    ele[7][27] != ele[35][27];
    ele[7][27] != ele[7][28];
    ele[7][27] != ele[7][29];
    ele[7][27] != ele[7][30];
    ele[7][27] != ele[7][31];
    ele[7][27] != ele[7][32];
    ele[7][27] != ele[7][33];
    ele[7][27] != ele[7][34];
    ele[7][27] != ele[7][35];
    ele[7][27] != ele[8][24];
    ele[7][27] != ele[8][25];
    ele[7][27] != ele[8][26];
    ele[7][27] != ele[8][27];
    ele[7][27] != ele[8][28];
    ele[7][27] != ele[8][29];
    ele[7][27] != ele[9][24];
    ele[7][27] != ele[9][25];
    ele[7][27] != ele[9][26];
    ele[7][27] != ele[9][27];
    ele[7][27] != ele[9][28];
    ele[7][27] != ele[9][29];
    ele[7][28] != ele[10][24];
    ele[7][28] != ele[10][25];
    ele[7][28] != ele[10][26];
    ele[7][28] != ele[10][27];
    ele[7][28] != ele[10][28];
    ele[7][28] != ele[10][29];
    ele[7][28] != ele[11][24];
    ele[7][28] != ele[11][25];
    ele[7][28] != ele[11][26];
    ele[7][28] != ele[11][27];
    ele[7][28] != ele[11][28];
    ele[7][28] != ele[11][29];
    ele[7][28] != ele[12][28];
    ele[7][28] != ele[13][28];
    ele[7][28] != ele[14][28];
    ele[7][28] != ele[15][28];
    ele[7][28] != ele[16][28];
    ele[7][28] != ele[17][28];
    ele[7][28] != ele[18][28];
    ele[7][28] != ele[19][28];
    ele[7][28] != ele[20][28];
    ele[7][28] != ele[21][28];
    ele[7][28] != ele[22][28];
    ele[7][28] != ele[23][28];
    ele[7][28] != ele[24][28];
    ele[7][28] != ele[25][28];
    ele[7][28] != ele[26][28];
    ele[7][28] != ele[27][28];
    ele[7][28] != ele[28][28];
    ele[7][28] != ele[29][28];
    ele[7][28] != ele[30][28];
    ele[7][28] != ele[31][28];
    ele[7][28] != ele[32][28];
    ele[7][28] != ele[33][28];
    ele[7][28] != ele[34][28];
    ele[7][28] != ele[35][28];
    ele[7][28] != ele[7][29];
    ele[7][28] != ele[7][30];
    ele[7][28] != ele[7][31];
    ele[7][28] != ele[7][32];
    ele[7][28] != ele[7][33];
    ele[7][28] != ele[7][34];
    ele[7][28] != ele[7][35];
    ele[7][28] != ele[8][24];
    ele[7][28] != ele[8][25];
    ele[7][28] != ele[8][26];
    ele[7][28] != ele[8][27];
    ele[7][28] != ele[8][28];
    ele[7][28] != ele[8][29];
    ele[7][28] != ele[9][24];
    ele[7][28] != ele[9][25];
    ele[7][28] != ele[9][26];
    ele[7][28] != ele[9][27];
    ele[7][28] != ele[9][28];
    ele[7][28] != ele[9][29];
    ele[7][29] != ele[10][24];
    ele[7][29] != ele[10][25];
    ele[7][29] != ele[10][26];
    ele[7][29] != ele[10][27];
    ele[7][29] != ele[10][28];
    ele[7][29] != ele[10][29];
    ele[7][29] != ele[11][24];
    ele[7][29] != ele[11][25];
    ele[7][29] != ele[11][26];
    ele[7][29] != ele[11][27];
    ele[7][29] != ele[11][28];
    ele[7][29] != ele[11][29];
    ele[7][29] != ele[12][29];
    ele[7][29] != ele[13][29];
    ele[7][29] != ele[14][29];
    ele[7][29] != ele[15][29];
    ele[7][29] != ele[16][29];
    ele[7][29] != ele[17][29];
    ele[7][29] != ele[18][29];
    ele[7][29] != ele[19][29];
    ele[7][29] != ele[20][29];
    ele[7][29] != ele[21][29];
    ele[7][29] != ele[22][29];
    ele[7][29] != ele[23][29];
    ele[7][29] != ele[24][29];
    ele[7][29] != ele[25][29];
    ele[7][29] != ele[26][29];
    ele[7][29] != ele[27][29];
    ele[7][29] != ele[28][29];
    ele[7][29] != ele[29][29];
    ele[7][29] != ele[30][29];
    ele[7][29] != ele[31][29];
    ele[7][29] != ele[32][29];
    ele[7][29] != ele[33][29];
    ele[7][29] != ele[34][29];
    ele[7][29] != ele[35][29];
    ele[7][29] != ele[7][30];
    ele[7][29] != ele[7][31];
    ele[7][29] != ele[7][32];
    ele[7][29] != ele[7][33];
    ele[7][29] != ele[7][34];
    ele[7][29] != ele[7][35];
    ele[7][29] != ele[8][24];
    ele[7][29] != ele[8][25];
    ele[7][29] != ele[8][26];
    ele[7][29] != ele[8][27];
    ele[7][29] != ele[8][28];
    ele[7][29] != ele[8][29];
    ele[7][29] != ele[9][24];
    ele[7][29] != ele[9][25];
    ele[7][29] != ele[9][26];
    ele[7][29] != ele[9][27];
    ele[7][29] != ele[9][28];
    ele[7][29] != ele[9][29];
    ele[7][3] != ele[10][0];
    ele[7][3] != ele[10][1];
    ele[7][3] != ele[10][2];
    ele[7][3] != ele[10][3];
    ele[7][3] != ele[10][4];
    ele[7][3] != ele[10][5];
    ele[7][3] != ele[11][0];
    ele[7][3] != ele[11][1];
    ele[7][3] != ele[11][2];
    ele[7][3] != ele[11][3];
    ele[7][3] != ele[11][4];
    ele[7][3] != ele[11][5];
    ele[7][3] != ele[12][3];
    ele[7][3] != ele[13][3];
    ele[7][3] != ele[14][3];
    ele[7][3] != ele[15][3];
    ele[7][3] != ele[16][3];
    ele[7][3] != ele[17][3];
    ele[7][3] != ele[18][3];
    ele[7][3] != ele[19][3];
    ele[7][3] != ele[20][3];
    ele[7][3] != ele[21][3];
    ele[7][3] != ele[22][3];
    ele[7][3] != ele[23][3];
    ele[7][3] != ele[24][3];
    ele[7][3] != ele[25][3];
    ele[7][3] != ele[26][3];
    ele[7][3] != ele[27][3];
    ele[7][3] != ele[28][3];
    ele[7][3] != ele[29][3];
    ele[7][3] != ele[30][3];
    ele[7][3] != ele[31][3];
    ele[7][3] != ele[32][3];
    ele[7][3] != ele[33][3];
    ele[7][3] != ele[34][3];
    ele[7][3] != ele[35][3];
    ele[7][3] != ele[7][10];
    ele[7][3] != ele[7][11];
    ele[7][3] != ele[7][12];
    ele[7][3] != ele[7][13];
    ele[7][3] != ele[7][14];
    ele[7][3] != ele[7][15];
    ele[7][3] != ele[7][16];
    ele[7][3] != ele[7][17];
    ele[7][3] != ele[7][18];
    ele[7][3] != ele[7][19];
    ele[7][3] != ele[7][20];
    ele[7][3] != ele[7][21];
    ele[7][3] != ele[7][22];
    ele[7][3] != ele[7][23];
    ele[7][3] != ele[7][24];
    ele[7][3] != ele[7][25];
    ele[7][3] != ele[7][26];
    ele[7][3] != ele[7][27];
    ele[7][3] != ele[7][28];
    ele[7][3] != ele[7][29];
    ele[7][3] != ele[7][30];
    ele[7][3] != ele[7][31];
    ele[7][3] != ele[7][32];
    ele[7][3] != ele[7][33];
    ele[7][3] != ele[7][34];
    ele[7][3] != ele[7][35];
    ele[7][3] != ele[7][4];
    ele[7][3] != ele[7][5];
    ele[7][3] != ele[7][6];
    ele[7][3] != ele[7][7];
    ele[7][3] != ele[7][8];
    ele[7][3] != ele[7][9];
    ele[7][3] != ele[8][0];
    ele[7][3] != ele[8][1];
    ele[7][3] != ele[8][2];
    ele[7][3] != ele[8][3];
    ele[7][3] != ele[8][4];
    ele[7][3] != ele[8][5];
    ele[7][3] != ele[9][0];
    ele[7][3] != ele[9][1];
    ele[7][3] != ele[9][2];
    ele[7][3] != ele[9][3];
    ele[7][3] != ele[9][4];
    ele[7][3] != ele[9][5];
    ele[7][30] != ele[10][30];
    ele[7][30] != ele[10][31];
    ele[7][30] != ele[10][32];
    ele[7][30] != ele[10][33];
    ele[7][30] != ele[10][34];
    ele[7][30] != ele[10][35];
    ele[7][30] != ele[11][30];
    ele[7][30] != ele[11][31];
    ele[7][30] != ele[11][32];
    ele[7][30] != ele[11][33];
    ele[7][30] != ele[11][34];
    ele[7][30] != ele[11][35];
    ele[7][30] != ele[12][30];
    ele[7][30] != ele[13][30];
    ele[7][30] != ele[14][30];
    ele[7][30] != ele[15][30];
    ele[7][30] != ele[16][30];
    ele[7][30] != ele[17][30];
    ele[7][30] != ele[18][30];
    ele[7][30] != ele[19][30];
    ele[7][30] != ele[20][30];
    ele[7][30] != ele[21][30];
    ele[7][30] != ele[22][30];
    ele[7][30] != ele[23][30];
    ele[7][30] != ele[24][30];
    ele[7][30] != ele[25][30];
    ele[7][30] != ele[26][30];
    ele[7][30] != ele[27][30];
    ele[7][30] != ele[28][30];
    ele[7][30] != ele[29][30];
    ele[7][30] != ele[30][30];
    ele[7][30] != ele[31][30];
    ele[7][30] != ele[32][30];
    ele[7][30] != ele[33][30];
    ele[7][30] != ele[34][30];
    ele[7][30] != ele[35][30];
    ele[7][30] != ele[7][31];
    ele[7][30] != ele[7][32];
    ele[7][30] != ele[7][33];
    ele[7][30] != ele[7][34];
    ele[7][30] != ele[7][35];
    ele[7][30] != ele[8][30];
    ele[7][30] != ele[8][31];
    ele[7][30] != ele[8][32];
    ele[7][30] != ele[8][33];
    ele[7][30] != ele[8][34];
    ele[7][30] != ele[8][35];
    ele[7][30] != ele[9][30];
    ele[7][30] != ele[9][31];
    ele[7][30] != ele[9][32];
    ele[7][30] != ele[9][33];
    ele[7][30] != ele[9][34];
    ele[7][30] != ele[9][35];
    ele[7][31] != ele[10][30];
    ele[7][31] != ele[10][31];
    ele[7][31] != ele[10][32];
    ele[7][31] != ele[10][33];
    ele[7][31] != ele[10][34];
    ele[7][31] != ele[10][35];
    ele[7][31] != ele[11][30];
    ele[7][31] != ele[11][31];
    ele[7][31] != ele[11][32];
    ele[7][31] != ele[11][33];
    ele[7][31] != ele[11][34];
    ele[7][31] != ele[11][35];
    ele[7][31] != ele[12][31];
    ele[7][31] != ele[13][31];
    ele[7][31] != ele[14][31];
    ele[7][31] != ele[15][31];
    ele[7][31] != ele[16][31];
    ele[7][31] != ele[17][31];
    ele[7][31] != ele[18][31];
    ele[7][31] != ele[19][31];
    ele[7][31] != ele[20][31];
    ele[7][31] != ele[21][31];
    ele[7][31] != ele[22][31];
    ele[7][31] != ele[23][31];
    ele[7][31] != ele[24][31];
    ele[7][31] != ele[25][31];
    ele[7][31] != ele[26][31];
    ele[7][31] != ele[27][31];
    ele[7][31] != ele[28][31];
    ele[7][31] != ele[29][31];
    ele[7][31] != ele[30][31];
    ele[7][31] != ele[31][31];
    ele[7][31] != ele[32][31];
    ele[7][31] != ele[33][31];
    ele[7][31] != ele[34][31];
    ele[7][31] != ele[35][31];
    ele[7][31] != ele[7][32];
    ele[7][31] != ele[7][33];
    ele[7][31] != ele[7][34];
    ele[7][31] != ele[7][35];
    ele[7][31] != ele[8][30];
    ele[7][31] != ele[8][31];
    ele[7][31] != ele[8][32];
    ele[7][31] != ele[8][33];
    ele[7][31] != ele[8][34];
    ele[7][31] != ele[8][35];
    ele[7][31] != ele[9][30];
    ele[7][31] != ele[9][31];
    ele[7][31] != ele[9][32];
    ele[7][31] != ele[9][33];
    ele[7][31] != ele[9][34];
    ele[7][31] != ele[9][35];
    ele[7][32] != ele[10][30];
    ele[7][32] != ele[10][31];
    ele[7][32] != ele[10][32];
    ele[7][32] != ele[10][33];
    ele[7][32] != ele[10][34];
    ele[7][32] != ele[10][35];
    ele[7][32] != ele[11][30];
    ele[7][32] != ele[11][31];
    ele[7][32] != ele[11][32];
    ele[7][32] != ele[11][33];
    ele[7][32] != ele[11][34];
    ele[7][32] != ele[11][35];
    ele[7][32] != ele[12][32];
    ele[7][32] != ele[13][32];
    ele[7][32] != ele[14][32];
    ele[7][32] != ele[15][32];
    ele[7][32] != ele[16][32];
    ele[7][32] != ele[17][32];
    ele[7][32] != ele[18][32];
    ele[7][32] != ele[19][32];
    ele[7][32] != ele[20][32];
    ele[7][32] != ele[21][32];
    ele[7][32] != ele[22][32];
    ele[7][32] != ele[23][32];
    ele[7][32] != ele[24][32];
    ele[7][32] != ele[25][32];
    ele[7][32] != ele[26][32];
    ele[7][32] != ele[27][32];
    ele[7][32] != ele[28][32];
    ele[7][32] != ele[29][32];
    ele[7][32] != ele[30][32];
    ele[7][32] != ele[31][32];
    ele[7][32] != ele[32][32];
    ele[7][32] != ele[33][32];
    ele[7][32] != ele[34][32];
    ele[7][32] != ele[35][32];
    ele[7][32] != ele[7][33];
    ele[7][32] != ele[7][34];
    ele[7][32] != ele[7][35];
    ele[7][32] != ele[8][30];
    ele[7][32] != ele[8][31];
    ele[7][32] != ele[8][32];
    ele[7][32] != ele[8][33];
    ele[7][32] != ele[8][34];
    ele[7][32] != ele[8][35];
    ele[7][32] != ele[9][30];
    ele[7][32] != ele[9][31];
    ele[7][32] != ele[9][32];
    ele[7][32] != ele[9][33];
    ele[7][32] != ele[9][34];
    ele[7][32] != ele[9][35];
    ele[7][33] != ele[10][30];
    ele[7][33] != ele[10][31];
    ele[7][33] != ele[10][32];
    ele[7][33] != ele[10][33];
    ele[7][33] != ele[10][34];
    ele[7][33] != ele[10][35];
    ele[7][33] != ele[11][30];
    ele[7][33] != ele[11][31];
    ele[7][33] != ele[11][32];
    ele[7][33] != ele[11][33];
    ele[7][33] != ele[11][34];
    ele[7][33] != ele[11][35];
    ele[7][33] != ele[12][33];
    ele[7][33] != ele[13][33];
    ele[7][33] != ele[14][33];
    ele[7][33] != ele[15][33];
    ele[7][33] != ele[16][33];
    ele[7][33] != ele[17][33];
    ele[7][33] != ele[18][33];
    ele[7][33] != ele[19][33];
    ele[7][33] != ele[20][33];
    ele[7][33] != ele[21][33];
    ele[7][33] != ele[22][33];
    ele[7][33] != ele[23][33];
    ele[7][33] != ele[24][33];
    ele[7][33] != ele[25][33];
    ele[7][33] != ele[26][33];
    ele[7][33] != ele[27][33];
    ele[7][33] != ele[28][33];
    ele[7][33] != ele[29][33];
    ele[7][33] != ele[30][33];
    ele[7][33] != ele[31][33];
    ele[7][33] != ele[32][33];
    ele[7][33] != ele[33][33];
    ele[7][33] != ele[34][33];
    ele[7][33] != ele[35][33];
    ele[7][33] != ele[7][34];
    ele[7][33] != ele[7][35];
    ele[7][33] != ele[8][30];
    ele[7][33] != ele[8][31];
    ele[7][33] != ele[8][32];
    ele[7][33] != ele[8][33];
    ele[7][33] != ele[8][34];
    ele[7][33] != ele[8][35];
    ele[7][33] != ele[9][30];
    ele[7][33] != ele[9][31];
    ele[7][33] != ele[9][32];
    ele[7][33] != ele[9][33];
    ele[7][33] != ele[9][34];
    ele[7][33] != ele[9][35];
    ele[7][34] != ele[10][30];
    ele[7][34] != ele[10][31];
    ele[7][34] != ele[10][32];
    ele[7][34] != ele[10][33];
    ele[7][34] != ele[10][34];
    ele[7][34] != ele[10][35];
    ele[7][34] != ele[11][30];
    ele[7][34] != ele[11][31];
    ele[7][34] != ele[11][32];
    ele[7][34] != ele[11][33];
    ele[7][34] != ele[11][34];
    ele[7][34] != ele[11][35];
    ele[7][34] != ele[12][34];
    ele[7][34] != ele[13][34];
    ele[7][34] != ele[14][34];
    ele[7][34] != ele[15][34];
    ele[7][34] != ele[16][34];
    ele[7][34] != ele[17][34];
    ele[7][34] != ele[18][34];
    ele[7][34] != ele[19][34];
    ele[7][34] != ele[20][34];
    ele[7][34] != ele[21][34];
    ele[7][34] != ele[22][34];
    ele[7][34] != ele[23][34];
    ele[7][34] != ele[24][34];
    ele[7][34] != ele[25][34];
    ele[7][34] != ele[26][34];
    ele[7][34] != ele[27][34];
    ele[7][34] != ele[28][34];
    ele[7][34] != ele[29][34];
    ele[7][34] != ele[30][34];
    ele[7][34] != ele[31][34];
    ele[7][34] != ele[32][34];
    ele[7][34] != ele[33][34];
    ele[7][34] != ele[34][34];
    ele[7][34] != ele[35][34];
    ele[7][34] != ele[7][35];
    ele[7][34] != ele[8][30];
    ele[7][34] != ele[8][31];
    ele[7][34] != ele[8][32];
    ele[7][34] != ele[8][33];
    ele[7][34] != ele[8][34];
    ele[7][34] != ele[8][35];
    ele[7][34] != ele[9][30];
    ele[7][34] != ele[9][31];
    ele[7][34] != ele[9][32];
    ele[7][34] != ele[9][33];
    ele[7][34] != ele[9][34];
    ele[7][34] != ele[9][35];
    ele[7][35] != ele[10][30];
    ele[7][35] != ele[10][31];
    ele[7][35] != ele[10][32];
    ele[7][35] != ele[10][33];
    ele[7][35] != ele[10][34];
    ele[7][35] != ele[10][35];
    ele[7][35] != ele[11][30];
    ele[7][35] != ele[11][31];
    ele[7][35] != ele[11][32];
    ele[7][35] != ele[11][33];
    ele[7][35] != ele[11][34];
    ele[7][35] != ele[11][35];
    ele[7][35] != ele[12][35];
    ele[7][35] != ele[13][35];
    ele[7][35] != ele[14][35];
    ele[7][35] != ele[15][35];
    ele[7][35] != ele[16][35];
    ele[7][35] != ele[17][35];
    ele[7][35] != ele[18][35];
    ele[7][35] != ele[19][35];
    ele[7][35] != ele[20][35];
    ele[7][35] != ele[21][35];
    ele[7][35] != ele[22][35];
    ele[7][35] != ele[23][35];
    ele[7][35] != ele[24][35];
    ele[7][35] != ele[25][35];
    ele[7][35] != ele[26][35];
    ele[7][35] != ele[27][35];
    ele[7][35] != ele[28][35];
    ele[7][35] != ele[29][35];
    ele[7][35] != ele[30][35];
    ele[7][35] != ele[31][35];
    ele[7][35] != ele[32][35];
    ele[7][35] != ele[33][35];
    ele[7][35] != ele[34][35];
    ele[7][35] != ele[35][35];
    ele[7][35] != ele[8][30];
    ele[7][35] != ele[8][31];
    ele[7][35] != ele[8][32];
    ele[7][35] != ele[8][33];
    ele[7][35] != ele[8][34];
    ele[7][35] != ele[8][35];
    ele[7][35] != ele[9][30];
    ele[7][35] != ele[9][31];
    ele[7][35] != ele[9][32];
    ele[7][35] != ele[9][33];
    ele[7][35] != ele[9][34];
    ele[7][35] != ele[9][35];
    ele[7][4] != ele[10][0];
    ele[7][4] != ele[10][1];
    ele[7][4] != ele[10][2];
    ele[7][4] != ele[10][3];
    ele[7][4] != ele[10][4];
    ele[7][4] != ele[10][5];
    ele[7][4] != ele[11][0];
    ele[7][4] != ele[11][1];
    ele[7][4] != ele[11][2];
    ele[7][4] != ele[11][3];
    ele[7][4] != ele[11][4];
    ele[7][4] != ele[11][5];
    ele[7][4] != ele[12][4];
    ele[7][4] != ele[13][4];
    ele[7][4] != ele[14][4];
    ele[7][4] != ele[15][4];
    ele[7][4] != ele[16][4];
    ele[7][4] != ele[17][4];
    ele[7][4] != ele[18][4];
    ele[7][4] != ele[19][4];
    ele[7][4] != ele[20][4];
    ele[7][4] != ele[21][4];
    ele[7][4] != ele[22][4];
    ele[7][4] != ele[23][4];
    ele[7][4] != ele[24][4];
    ele[7][4] != ele[25][4];
    ele[7][4] != ele[26][4];
    ele[7][4] != ele[27][4];
    ele[7][4] != ele[28][4];
    ele[7][4] != ele[29][4];
    ele[7][4] != ele[30][4];
    ele[7][4] != ele[31][4];
    ele[7][4] != ele[32][4];
    ele[7][4] != ele[33][4];
    ele[7][4] != ele[34][4];
    ele[7][4] != ele[35][4];
    ele[7][4] != ele[7][10];
    ele[7][4] != ele[7][11];
    ele[7][4] != ele[7][12];
    ele[7][4] != ele[7][13];
    ele[7][4] != ele[7][14];
    ele[7][4] != ele[7][15];
    ele[7][4] != ele[7][16];
    ele[7][4] != ele[7][17];
    ele[7][4] != ele[7][18];
    ele[7][4] != ele[7][19];
    ele[7][4] != ele[7][20];
    ele[7][4] != ele[7][21];
    ele[7][4] != ele[7][22];
    ele[7][4] != ele[7][23];
    ele[7][4] != ele[7][24];
    ele[7][4] != ele[7][25];
    ele[7][4] != ele[7][26];
    ele[7][4] != ele[7][27];
    ele[7][4] != ele[7][28];
    ele[7][4] != ele[7][29];
    ele[7][4] != ele[7][30];
    ele[7][4] != ele[7][31];
    ele[7][4] != ele[7][32];
    ele[7][4] != ele[7][33];
    ele[7][4] != ele[7][34];
    ele[7][4] != ele[7][35];
    ele[7][4] != ele[7][5];
    ele[7][4] != ele[7][6];
    ele[7][4] != ele[7][7];
    ele[7][4] != ele[7][8];
    ele[7][4] != ele[7][9];
    ele[7][4] != ele[8][0];
    ele[7][4] != ele[8][1];
    ele[7][4] != ele[8][2];
    ele[7][4] != ele[8][3];
    ele[7][4] != ele[8][4];
    ele[7][4] != ele[8][5];
    ele[7][4] != ele[9][0];
    ele[7][4] != ele[9][1];
    ele[7][4] != ele[9][2];
    ele[7][4] != ele[9][3];
    ele[7][4] != ele[9][4];
    ele[7][4] != ele[9][5];
    ele[7][5] != ele[10][0];
    ele[7][5] != ele[10][1];
    ele[7][5] != ele[10][2];
    ele[7][5] != ele[10][3];
    ele[7][5] != ele[10][4];
    ele[7][5] != ele[10][5];
    ele[7][5] != ele[11][0];
    ele[7][5] != ele[11][1];
    ele[7][5] != ele[11][2];
    ele[7][5] != ele[11][3];
    ele[7][5] != ele[11][4];
    ele[7][5] != ele[11][5];
    ele[7][5] != ele[12][5];
    ele[7][5] != ele[13][5];
    ele[7][5] != ele[14][5];
    ele[7][5] != ele[15][5];
    ele[7][5] != ele[16][5];
    ele[7][5] != ele[17][5];
    ele[7][5] != ele[18][5];
    ele[7][5] != ele[19][5];
    ele[7][5] != ele[20][5];
    ele[7][5] != ele[21][5];
    ele[7][5] != ele[22][5];
    ele[7][5] != ele[23][5];
    ele[7][5] != ele[24][5];
    ele[7][5] != ele[25][5];
    ele[7][5] != ele[26][5];
    ele[7][5] != ele[27][5];
    ele[7][5] != ele[28][5];
    ele[7][5] != ele[29][5];
    ele[7][5] != ele[30][5];
    ele[7][5] != ele[31][5];
    ele[7][5] != ele[32][5];
    ele[7][5] != ele[33][5];
    ele[7][5] != ele[34][5];
    ele[7][5] != ele[35][5];
    ele[7][5] != ele[7][10];
    ele[7][5] != ele[7][11];
    ele[7][5] != ele[7][12];
    ele[7][5] != ele[7][13];
    ele[7][5] != ele[7][14];
    ele[7][5] != ele[7][15];
    ele[7][5] != ele[7][16];
    ele[7][5] != ele[7][17];
    ele[7][5] != ele[7][18];
    ele[7][5] != ele[7][19];
    ele[7][5] != ele[7][20];
    ele[7][5] != ele[7][21];
    ele[7][5] != ele[7][22];
    ele[7][5] != ele[7][23];
    ele[7][5] != ele[7][24];
    ele[7][5] != ele[7][25];
    ele[7][5] != ele[7][26];
    ele[7][5] != ele[7][27];
    ele[7][5] != ele[7][28];
    ele[7][5] != ele[7][29];
    ele[7][5] != ele[7][30];
    ele[7][5] != ele[7][31];
    ele[7][5] != ele[7][32];
    ele[7][5] != ele[7][33];
    ele[7][5] != ele[7][34];
    ele[7][5] != ele[7][35];
    ele[7][5] != ele[7][6];
    ele[7][5] != ele[7][7];
    ele[7][5] != ele[7][8];
    ele[7][5] != ele[7][9];
    ele[7][5] != ele[8][0];
    ele[7][5] != ele[8][1];
    ele[7][5] != ele[8][2];
    ele[7][5] != ele[8][3];
    ele[7][5] != ele[8][4];
    ele[7][5] != ele[8][5];
    ele[7][5] != ele[9][0];
    ele[7][5] != ele[9][1];
    ele[7][5] != ele[9][2];
    ele[7][5] != ele[9][3];
    ele[7][5] != ele[9][4];
    ele[7][5] != ele[9][5];
    ele[7][6] != ele[10][10];
    ele[7][6] != ele[10][11];
    ele[7][6] != ele[10][6];
    ele[7][6] != ele[10][7];
    ele[7][6] != ele[10][8];
    ele[7][6] != ele[10][9];
    ele[7][6] != ele[11][10];
    ele[7][6] != ele[11][11];
    ele[7][6] != ele[11][6];
    ele[7][6] != ele[11][7];
    ele[7][6] != ele[11][8];
    ele[7][6] != ele[11][9];
    ele[7][6] != ele[12][6];
    ele[7][6] != ele[13][6];
    ele[7][6] != ele[14][6];
    ele[7][6] != ele[15][6];
    ele[7][6] != ele[16][6];
    ele[7][6] != ele[17][6];
    ele[7][6] != ele[18][6];
    ele[7][6] != ele[19][6];
    ele[7][6] != ele[20][6];
    ele[7][6] != ele[21][6];
    ele[7][6] != ele[22][6];
    ele[7][6] != ele[23][6];
    ele[7][6] != ele[24][6];
    ele[7][6] != ele[25][6];
    ele[7][6] != ele[26][6];
    ele[7][6] != ele[27][6];
    ele[7][6] != ele[28][6];
    ele[7][6] != ele[29][6];
    ele[7][6] != ele[30][6];
    ele[7][6] != ele[31][6];
    ele[7][6] != ele[32][6];
    ele[7][6] != ele[33][6];
    ele[7][6] != ele[34][6];
    ele[7][6] != ele[35][6];
    ele[7][6] != ele[7][10];
    ele[7][6] != ele[7][11];
    ele[7][6] != ele[7][12];
    ele[7][6] != ele[7][13];
    ele[7][6] != ele[7][14];
    ele[7][6] != ele[7][15];
    ele[7][6] != ele[7][16];
    ele[7][6] != ele[7][17];
    ele[7][6] != ele[7][18];
    ele[7][6] != ele[7][19];
    ele[7][6] != ele[7][20];
    ele[7][6] != ele[7][21];
    ele[7][6] != ele[7][22];
    ele[7][6] != ele[7][23];
    ele[7][6] != ele[7][24];
    ele[7][6] != ele[7][25];
    ele[7][6] != ele[7][26];
    ele[7][6] != ele[7][27];
    ele[7][6] != ele[7][28];
    ele[7][6] != ele[7][29];
    ele[7][6] != ele[7][30];
    ele[7][6] != ele[7][31];
    ele[7][6] != ele[7][32];
    ele[7][6] != ele[7][33];
    ele[7][6] != ele[7][34];
    ele[7][6] != ele[7][35];
    ele[7][6] != ele[7][7];
    ele[7][6] != ele[7][8];
    ele[7][6] != ele[7][9];
    ele[7][6] != ele[8][10];
    ele[7][6] != ele[8][11];
    ele[7][6] != ele[8][6];
    ele[7][6] != ele[8][7];
    ele[7][6] != ele[8][8];
    ele[7][6] != ele[8][9];
    ele[7][6] != ele[9][10];
    ele[7][6] != ele[9][11];
    ele[7][6] != ele[9][6];
    ele[7][6] != ele[9][7];
    ele[7][6] != ele[9][8];
    ele[7][6] != ele[9][9];
    ele[7][7] != ele[10][10];
    ele[7][7] != ele[10][11];
    ele[7][7] != ele[10][6];
    ele[7][7] != ele[10][7];
    ele[7][7] != ele[10][8];
    ele[7][7] != ele[10][9];
    ele[7][7] != ele[11][10];
    ele[7][7] != ele[11][11];
    ele[7][7] != ele[11][6];
    ele[7][7] != ele[11][7];
    ele[7][7] != ele[11][8];
    ele[7][7] != ele[11][9];
    ele[7][7] != ele[12][7];
    ele[7][7] != ele[13][7];
    ele[7][7] != ele[14][7];
    ele[7][7] != ele[15][7];
    ele[7][7] != ele[16][7];
    ele[7][7] != ele[17][7];
    ele[7][7] != ele[18][7];
    ele[7][7] != ele[19][7];
    ele[7][7] != ele[20][7];
    ele[7][7] != ele[21][7];
    ele[7][7] != ele[22][7];
    ele[7][7] != ele[23][7];
    ele[7][7] != ele[24][7];
    ele[7][7] != ele[25][7];
    ele[7][7] != ele[26][7];
    ele[7][7] != ele[27][7];
    ele[7][7] != ele[28][7];
    ele[7][7] != ele[29][7];
    ele[7][7] != ele[30][7];
    ele[7][7] != ele[31][7];
    ele[7][7] != ele[32][7];
    ele[7][7] != ele[33][7];
    ele[7][7] != ele[34][7];
    ele[7][7] != ele[35][7];
    ele[7][7] != ele[7][10];
    ele[7][7] != ele[7][11];
    ele[7][7] != ele[7][12];
    ele[7][7] != ele[7][13];
    ele[7][7] != ele[7][14];
    ele[7][7] != ele[7][15];
    ele[7][7] != ele[7][16];
    ele[7][7] != ele[7][17];
    ele[7][7] != ele[7][18];
    ele[7][7] != ele[7][19];
    ele[7][7] != ele[7][20];
    ele[7][7] != ele[7][21];
    ele[7][7] != ele[7][22];
    ele[7][7] != ele[7][23];
    ele[7][7] != ele[7][24];
    ele[7][7] != ele[7][25];
    ele[7][7] != ele[7][26];
    ele[7][7] != ele[7][27];
    ele[7][7] != ele[7][28];
    ele[7][7] != ele[7][29];
    ele[7][7] != ele[7][30];
    ele[7][7] != ele[7][31];
    ele[7][7] != ele[7][32];
    ele[7][7] != ele[7][33];
    ele[7][7] != ele[7][34];
    ele[7][7] != ele[7][35];
    ele[7][7] != ele[7][8];
    ele[7][7] != ele[7][9];
    ele[7][7] != ele[8][10];
    ele[7][7] != ele[8][11];
    ele[7][7] != ele[8][6];
    ele[7][7] != ele[8][7];
    ele[7][7] != ele[8][8];
    ele[7][7] != ele[8][9];
    ele[7][7] != ele[9][10];
    ele[7][7] != ele[9][11];
    ele[7][7] != ele[9][6];
    ele[7][7] != ele[9][7];
    ele[7][7] != ele[9][8];
    ele[7][7] != ele[9][9];
    ele[7][8] != ele[10][10];
    ele[7][8] != ele[10][11];
    ele[7][8] != ele[10][6];
    ele[7][8] != ele[10][7];
    ele[7][8] != ele[10][8];
    ele[7][8] != ele[10][9];
    ele[7][8] != ele[11][10];
    ele[7][8] != ele[11][11];
    ele[7][8] != ele[11][6];
    ele[7][8] != ele[11][7];
    ele[7][8] != ele[11][8];
    ele[7][8] != ele[11][9];
    ele[7][8] != ele[12][8];
    ele[7][8] != ele[13][8];
    ele[7][8] != ele[14][8];
    ele[7][8] != ele[15][8];
    ele[7][8] != ele[16][8];
    ele[7][8] != ele[17][8];
    ele[7][8] != ele[18][8];
    ele[7][8] != ele[19][8];
    ele[7][8] != ele[20][8];
    ele[7][8] != ele[21][8];
    ele[7][8] != ele[22][8];
    ele[7][8] != ele[23][8];
    ele[7][8] != ele[24][8];
    ele[7][8] != ele[25][8];
    ele[7][8] != ele[26][8];
    ele[7][8] != ele[27][8];
    ele[7][8] != ele[28][8];
    ele[7][8] != ele[29][8];
    ele[7][8] != ele[30][8];
    ele[7][8] != ele[31][8];
    ele[7][8] != ele[32][8];
    ele[7][8] != ele[33][8];
    ele[7][8] != ele[34][8];
    ele[7][8] != ele[35][8];
    ele[7][8] != ele[7][10];
    ele[7][8] != ele[7][11];
    ele[7][8] != ele[7][12];
    ele[7][8] != ele[7][13];
    ele[7][8] != ele[7][14];
    ele[7][8] != ele[7][15];
    ele[7][8] != ele[7][16];
    ele[7][8] != ele[7][17];
    ele[7][8] != ele[7][18];
    ele[7][8] != ele[7][19];
    ele[7][8] != ele[7][20];
    ele[7][8] != ele[7][21];
    ele[7][8] != ele[7][22];
    ele[7][8] != ele[7][23];
    ele[7][8] != ele[7][24];
    ele[7][8] != ele[7][25];
    ele[7][8] != ele[7][26];
    ele[7][8] != ele[7][27];
    ele[7][8] != ele[7][28];
    ele[7][8] != ele[7][29];
    ele[7][8] != ele[7][30];
    ele[7][8] != ele[7][31];
    ele[7][8] != ele[7][32];
    ele[7][8] != ele[7][33];
    ele[7][8] != ele[7][34];
    ele[7][8] != ele[7][35];
    ele[7][8] != ele[7][9];
    ele[7][8] != ele[8][10];
    ele[7][8] != ele[8][11];
    ele[7][8] != ele[8][6];
    ele[7][8] != ele[8][7];
    ele[7][8] != ele[8][8];
    ele[7][8] != ele[8][9];
    ele[7][8] != ele[9][10];
    ele[7][8] != ele[9][11];
    ele[7][8] != ele[9][6];
    ele[7][8] != ele[9][7];
    ele[7][8] != ele[9][8];
    ele[7][8] != ele[9][9];
    ele[7][9] != ele[10][10];
    ele[7][9] != ele[10][11];
    ele[7][9] != ele[10][6];
    ele[7][9] != ele[10][7];
    ele[7][9] != ele[10][8];
    ele[7][9] != ele[10][9];
    ele[7][9] != ele[11][10];
    ele[7][9] != ele[11][11];
    ele[7][9] != ele[11][6];
    ele[7][9] != ele[11][7];
    ele[7][9] != ele[11][8];
    ele[7][9] != ele[11][9];
    ele[7][9] != ele[12][9];
    ele[7][9] != ele[13][9];
    ele[7][9] != ele[14][9];
    ele[7][9] != ele[15][9];
    ele[7][9] != ele[16][9];
    ele[7][9] != ele[17][9];
    ele[7][9] != ele[18][9];
    ele[7][9] != ele[19][9];
    ele[7][9] != ele[20][9];
    ele[7][9] != ele[21][9];
    ele[7][9] != ele[22][9];
    ele[7][9] != ele[23][9];
    ele[7][9] != ele[24][9];
    ele[7][9] != ele[25][9];
    ele[7][9] != ele[26][9];
    ele[7][9] != ele[27][9];
    ele[7][9] != ele[28][9];
    ele[7][9] != ele[29][9];
    ele[7][9] != ele[30][9];
    ele[7][9] != ele[31][9];
    ele[7][9] != ele[32][9];
    ele[7][9] != ele[33][9];
    ele[7][9] != ele[34][9];
    ele[7][9] != ele[35][9];
    ele[7][9] != ele[7][10];
    ele[7][9] != ele[7][11];
    ele[7][9] != ele[7][12];
    ele[7][9] != ele[7][13];
    ele[7][9] != ele[7][14];
    ele[7][9] != ele[7][15];
    ele[7][9] != ele[7][16];
    ele[7][9] != ele[7][17];
    ele[7][9] != ele[7][18];
    ele[7][9] != ele[7][19];
    ele[7][9] != ele[7][20];
    ele[7][9] != ele[7][21];
    ele[7][9] != ele[7][22];
    ele[7][9] != ele[7][23];
    ele[7][9] != ele[7][24];
    ele[7][9] != ele[7][25];
    ele[7][9] != ele[7][26];
    ele[7][9] != ele[7][27];
    ele[7][9] != ele[7][28];
    ele[7][9] != ele[7][29];
    ele[7][9] != ele[7][30];
    ele[7][9] != ele[7][31];
    ele[7][9] != ele[7][32];
    ele[7][9] != ele[7][33];
    ele[7][9] != ele[7][34];
    ele[7][9] != ele[7][35];
    ele[7][9] != ele[8][10];
    ele[7][9] != ele[8][11];
    ele[7][9] != ele[8][6];
    ele[7][9] != ele[8][7];
    ele[7][9] != ele[8][8];
    ele[7][9] != ele[8][9];
    ele[7][9] != ele[9][10];
    ele[7][9] != ele[9][11];
    ele[7][9] != ele[9][6];
    ele[7][9] != ele[9][7];
    ele[7][9] != ele[9][8];
    ele[7][9] != ele[9][9];
    ele[8][0] != ele[10][0];
    ele[8][0] != ele[10][1];
    ele[8][0] != ele[10][2];
    ele[8][0] != ele[10][3];
    ele[8][0] != ele[10][4];
    ele[8][0] != ele[10][5];
    ele[8][0] != ele[11][0];
    ele[8][0] != ele[11][1];
    ele[8][0] != ele[11][2];
    ele[8][0] != ele[11][3];
    ele[8][0] != ele[11][4];
    ele[8][0] != ele[11][5];
    ele[8][0] != ele[12][0];
    ele[8][0] != ele[13][0];
    ele[8][0] != ele[14][0];
    ele[8][0] != ele[15][0];
    ele[8][0] != ele[16][0];
    ele[8][0] != ele[17][0];
    ele[8][0] != ele[18][0];
    ele[8][0] != ele[19][0];
    ele[8][0] != ele[20][0];
    ele[8][0] != ele[21][0];
    ele[8][0] != ele[22][0];
    ele[8][0] != ele[23][0];
    ele[8][0] != ele[24][0];
    ele[8][0] != ele[25][0];
    ele[8][0] != ele[26][0];
    ele[8][0] != ele[27][0];
    ele[8][0] != ele[28][0];
    ele[8][0] != ele[29][0];
    ele[8][0] != ele[30][0];
    ele[8][0] != ele[31][0];
    ele[8][0] != ele[32][0];
    ele[8][0] != ele[33][0];
    ele[8][0] != ele[34][0];
    ele[8][0] != ele[35][0];
    ele[8][0] != ele[8][1];
    ele[8][0] != ele[8][10];
    ele[8][0] != ele[8][11];
    ele[8][0] != ele[8][12];
    ele[8][0] != ele[8][13];
    ele[8][0] != ele[8][14];
    ele[8][0] != ele[8][15];
    ele[8][0] != ele[8][16];
    ele[8][0] != ele[8][17];
    ele[8][0] != ele[8][18];
    ele[8][0] != ele[8][19];
    ele[8][0] != ele[8][2];
    ele[8][0] != ele[8][20];
    ele[8][0] != ele[8][21];
    ele[8][0] != ele[8][22];
    ele[8][0] != ele[8][23];
    ele[8][0] != ele[8][24];
    ele[8][0] != ele[8][25];
    ele[8][0] != ele[8][26];
    ele[8][0] != ele[8][27];
    ele[8][0] != ele[8][28];
    ele[8][0] != ele[8][29];
    ele[8][0] != ele[8][3];
    ele[8][0] != ele[8][30];
    ele[8][0] != ele[8][31];
    ele[8][0] != ele[8][32];
    ele[8][0] != ele[8][33];
    ele[8][0] != ele[8][34];
    ele[8][0] != ele[8][35];
    ele[8][0] != ele[8][4];
    ele[8][0] != ele[8][5];
    ele[8][0] != ele[8][6];
    ele[8][0] != ele[8][7];
    ele[8][0] != ele[8][8];
    ele[8][0] != ele[8][9];
    ele[8][0] != ele[9][0];
    ele[8][0] != ele[9][1];
    ele[8][0] != ele[9][2];
    ele[8][0] != ele[9][3];
    ele[8][0] != ele[9][4];
    ele[8][0] != ele[9][5];
    ele[8][1] != ele[10][0];
    ele[8][1] != ele[10][1];
    ele[8][1] != ele[10][2];
    ele[8][1] != ele[10][3];
    ele[8][1] != ele[10][4];
    ele[8][1] != ele[10][5];
    ele[8][1] != ele[11][0];
    ele[8][1] != ele[11][1];
    ele[8][1] != ele[11][2];
    ele[8][1] != ele[11][3];
    ele[8][1] != ele[11][4];
    ele[8][1] != ele[11][5];
    ele[8][1] != ele[12][1];
    ele[8][1] != ele[13][1];
    ele[8][1] != ele[14][1];
    ele[8][1] != ele[15][1];
    ele[8][1] != ele[16][1];
    ele[8][1] != ele[17][1];
    ele[8][1] != ele[18][1];
    ele[8][1] != ele[19][1];
    ele[8][1] != ele[20][1];
    ele[8][1] != ele[21][1];
    ele[8][1] != ele[22][1];
    ele[8][1] != ele[23][1];
    ele[8][1] != ele[24][1];
    ele[8][1] != ele[25][1];
    ele[8][1] != ele[26][1];
    ele[8][1] != ele[27][1];
    ele[8][1] != ele[28][1];
    ele[8][1] != ele[29][1];
    ele[8][1] != ele[30][1];
    ele[8][1] != ele[31][1];
    ele[8][1] != ele[32][1];
    ele[8][1] != ele[33][1];
    ele[8][1] != ele[34][1];
    ele[8][1] != ele[35][1];
    ele[8][1] != ele[8][10];
    ele[8][1] != ele[8][11];
    ele[8][1] != ele[8][12];
    ele[8][1] != ele[8][13];
    ele[8][1] != ele[8][14];
    ele[8][1] != ele[8][15];
    ele[8][1] != ele[8][16];
    ele[8][1] != ele[8][17];
    ele[8][1] != ele[8][18];
    ele[8][1] != ele[8][19];
    ele[8][1] != ele[8][2];
    ele[8][1] != ele[8][20];
    ele[8][1] != ele[8][21];
    ele[8][1] != ele[8][22];
    ele[8][1] != ele[8][23];
    ele[8][1] != ele[8][24];
    ele[8][1] != ele[8][25];
    ele[8][1] != ele[8][26];
    ele[8][1] != ele[8][27];
    ele[8][1] != ele[8][28];
    ele[8][1] != ele[8][29];
    ele[8][1] != ele[8][3];
    ele[8][1] != ele[8][30];
    ele[8][1] != ele[8][31];
    ele[8][1] != ele[8][32];
    ele[8][1] != ele[8][33];
    ele[8][1] != ele[8][34];
    ele[8][1] != ele[8][35];
    ele[8][1] != ele[8][4];
    ele[8][1] != ele[8][5];
    ele[8][1] != ele[8][6];
    ele[8][1] != ele[8][7];
    ele[8][1] != ele[8][8];
    ele[8][1] != ele[8][9];
    ele[8][1] != ele[9][0];
    ele[8][1] != ele[9][1];
    ele[8][1] != ele[9][2];
    ele[8][1] != ele[9][3];
    ele[8][1] != ele[9][4];
    ele[8][1] != ele[9][5];
    ele[8][10] != ele[10][10];
    ele[8][10] != ele[10][11];
    ele[8][10] != ele[10][6];
    ele[8][10] != ele[10][7];
    ele[8][10] != ele[10][8];
    ele[8][10] != ele[10][9];
    ele[8][10] != ele[11][10];
    ele[8][10] != ele[11][11];
    ele[8][10] != ele[11][6];
    ele[8][10] != ele[11][7];
    ele[8][10] != ele[11][8];
    ele[8][10] != ele[11][9];
    ele[8][10] != ele[12][10];
    ele[8][10] != ele[13][10];
    ele[8][10] != ele[14][10];
    ele[8][10] != ele[15][10];
    ele[8][10] != ele[16][10];
    ele[8][10] != ele[17][10];
    ele[8][10] != ele[18][10];
    ele[8][10] != ele[19][10];
    ele[8][10] != ele[20][10];
    ele[8][10] != ele[21][10];
    ele[8][10] != ele[22][10];
    ele[8][10] != ele[23][10];
    ele[8][10] != ele[24][10];
    ele[8][10] != ele[25][10];
    ele[8][10] != ele[26][10];
    ele[8][10] != ele[27][10];
    ele[8][10] != ele[28][10];
    ele[8][10] != ele[29][10];
    ele[8][10] != ele[30][10];
    ele[8][10] != ele[31][10];
    ele[8][10] != ele[32][10];
    ele[8][10] != ele[33][10];
    ele[8][10] != ele[34][10];
    ele[8][10] != ele[35][10];
    ele[8][10] != ele[8][11];
    ele[8][10] != ele[8][12];
    ele[8][10] != ele[8][13];
    ele[8][10] != ele[8][14];
    ele[8][10] != ele[8][15];
    ele[8][10] != ele[8][16];
    ele[8][10] != ele[8][17];
    ele[8][10] != ele[8][18];
    ele[8][10] != ele[8][19];
    ele[8][10] != ele[8][20];
    ele[8][10] != ele[8][21];
    ele[8][10] != ele[8][22];
    ele[8][10] != ele[8][23];
    ele[8][10] != ele[8][24];
    ele[8][10] != ele[8][25];
    ele[8][10] != ele[8][26];
    ele[8][10] != ele[8][27];
    ele[8][10] != ele[8][28];
    ele[8][10] != ele[8][29];
    ele[8][10] != ele[8][30];
    ele[8][10] != ele[8][31];
    ele[8][10] != ele[8][32];
    ele[8][10] != ele[8][33];
    ele[8][10] != ele[8][34];
    ele[8][10] != ele[8][35];
    ele[8][10] != ele[9][10];
    ele[8][10] != ele[9][11];
    ele[8][10] != ele[9][6];
    ele[8][10] != ele[9][7];
    ele[8][10] != ele[9][8];
    ele[8][10] != ele[9][9];
    ele[8][11] != ele[10][10];
    ele[8][11] != ele[10][11];
    ele[8][11] != ele[10][6];
    ele[8][11] != ele[10][7];
    ele[8][11] != ele[10][8];
    ele[8][11] != ele[10][9];
    ele[8][11] != ele[11][10];
    ele[8][11] != ele[11][11];
    ele[8][11] != ele[11][6];
    ele[8][11] != ele[11][7];
    ele[8][11] != ele[11][8];
    ele[8][11] != ele[11][9];
    ele[8][11] != ele[12][11];
    ele[8][11] != ele[13][11];
    ele[8][11] != ele[14][11];
    ele[8][11] != ele[15][11];
    ele[8][11] != ele[16][11];
    ele[8][11] != ele[17][11];
    ele[8][11] != ele[18][11];
    ele[8][11] != ele[19][11];
    ele[8][11] != ele[20][11];
    ele[8][11] != ele[21][11];
    ele[8][11] != ele[22][11];
    ele[8][11] != ele[23][11];
    ele[8][11] != ele[24][11];
    ele[8][11] != ele[25][11];
    ele[8][11] != ele[26][11];
    ele[8][11] != ele[27][11];
    ele[8][11] != ele[28][11];
    ele[8][11] != ele[29][11];
    ele[8][11] != ele[30][11];
    ele[8][11] != ele[31][11];
    ele[8][11] != ele[32][11];
    ele[8][11] != ele[33][11];
    ele[8][11] != ele[34][11];
    ele[8][11] != ele[35][11];
    ele[8][11] != ele[8][12];
    ele[8][11] != ele[8][13];
    ele[8][11] != ele[8][14];
    ele[8][11] != ele[8][15];
    ele[8][11] != ele[8][16];
    ele[8][11] != ele[8][17];
    ele[8][11] != ele[8][18];
    ele[8][11] != ele[8][19];
    ele[8][11] != ele[8][20];
    ele[8][11] != ele[8][21];
    ele[8][11] != ele[8][22];
    ele[8][11] != ele[8][23];
    ele[8][11] != ele[8][24];
    ele[8][11] != ele[8][25];
    ele[8][11] != ele[8][26];
    ele[8][11] != ele[8][27];
    ele[8][11] != ele[8][28];
    ele[8][11] != ele[8][29];
    ele[8][11] != ele[8][30];
    ele[8][11] != ele[8][31];
    ele[8][11] != ele[8][32];
    ele[8][11] != ele[8][33];
    ele[8][11] != ele[8][34];
    ele[8][11] != ele[8][35];
    ele[8][11] != ele[9][10];
    ele[8][11] != ele[9][11];
    ele[8][11] != ele[9][6];
    ele[8][11] != ele[9][7];
    ele[8][11] != ele[9][8];
    ele[8][11] != ele[9][9];
    ele[8][12] != ele[10][12];
    ele[8][12] != ele[10][13];
    ele[8][12] != ele[10][14];
    ele[8][12] != ele[10][15];
    ele[8][12] != ele[10][16];
    ele[8][12] != ele[10][17];
    ele[8][12] != ele[11][12];
    ele[8][12] != ele[11][13];
    ele[8][12] != ele[11][14];
    ele[8][12] != ele[11][15];
    ele[8][12] != ele[11][16];
    ele[8][12] != ele[11][17];
    ele[8][12] != ele[12][12];
    ele[8][12] != ele[13][12];
    ele[8][12] != ele[14][12];
    ele[8][12] != ele[15][12];
    ele[8][12] != ele[16][12];
    ele[8][12] != ele[17][12];
    ele[8][12] != ele[18][12];
    ele[8][12] != ele[19][12];
    ele[8][12] != ele[20][12];
    ele[8][12] != ele[21][12];
    ele[8][12] != ele[22][12];
    ele[8][12] != ele[23][12];
    ele[8][12] != ele[24][12];
    ele[8][12] != ele[25][12];
    ele[8][12] != ele[26][12];
    ele[8][12] != ele[27][12];
    ele[8][12] != ele[28][12];
    ele[8][12] != ele[29][12];
    ele[8][12] != ele[30][12];
    ele[8][12] != ele[31][12];
    ele[8][12] != ele[32][12];
    ele[8][12] != ele[33][12];
    ele[8][12] != ele[34][12];
    ele[8][12] != ele[35][12];
    ele[8][12] != ele[8][13];
    ele[8][12] != ele[8][14];
    ele[8][12] != ele[8][15];
    ele[8][12] != ele[8][16];
    ele[8][12] != ele[8][17];
    ele[8][12] != ele[8][18];
    ele[8][12] != ele[8][19];
    ele[8][12] != ele[8][20];
    ele[8][12] != ele[8][21];
    ele[8][12] != ele[8][22];
    ele[8][12] != ele[8][23];
    ele[8][12] != ele[8][24];
    ele[8][12] != ele[8][25];
    ele[8][12] != ele[8][26];
    ele[8][12] != ele[8][27];
    ele[8][12] != ele[8][28];
    ele[8][12] != ele[8][29];
    ele[8][12] != ele[8][30];
    ele[8][12] != ele[8][31];
    ele[8][12] != ele[8][32];
    ele[8][12] != ele[8][33];
    ele[8][12] != ele[8][34];
    ele[8][12] != ele[8][35];
    ele[8][12] != ele[9][12];
    ele[8][12] != ele[9][13];
    ele[8][12] != ele[9][14];
    ele[8][12] != ele[9][15];
    ele[8][12] != ele[9][16];
    ele[8][12] != ele[9][17];
    ele[8][13] != ele[10][12];
    ele[8][13] != ele[10][13];
    ele[8][13] != ele[10][14];
    ele[8][13] != ele[10][15];
    ele[8][13] != ele[10][16];
    ele[8][13] != ele[10][17];
    ele[8][13] != ele[11][12];
    ele[8][13] != ele[11][13];
    ele[8][13] != ele[11][14];
    ele[8][13] != ele[11][15];
    ele[8][13] != ele[11][16];
    ele[8][13] != ele[11][17];
    ele[8][13] != ele[12][13];
    ele[8][13] != ele[13][13];
    ele[8][13] != ele[14][13];
    ele[8][13] != ele[15][13];
    ele[8][13] != ele[16][13];
    ele[8][13] != ele[17][13];
    ele[8][13] != ele[18][13];
    ele[8][13] != ele[19][13];
    ele[8][13] != ele[20][13];
    ele[8][13] != ele[21][13];
    ele[8][13] != ele[22][13];
    ele[8][13] != ele[23][13];
    ele[8][13] != ele[24][13];
    ele[8][13] != ele[25][13];
    ele[8][13] != ele[26][13];
    ele[8][13] != ele[27][13];
    ele[8][13] != ele[28][13];
    ele[8][13] != ele[29][13];
    ele[8][13] != ele[30][13];
    ele[8][13] != ele[31][13];
    ele[8][13] != ele[32][13];
    ele[8][13] != ele[33][13];
    ele[8][13] != ele[34][13];
    ele[8][13] != ele[35][13];
    ele[8][13] != ele[8][14];
    ele[8][13] != ele[8][15];
    ele[8][13] != ele[8][16];
    ele[8][13] != ele[8][17];
    ele[8][13] != ele[8][18];
    ele[8][13] != ele[8][19];
    ele[8][13] != ele[8][20];
    ele[8][13] != ele[8][21];
    ele[8][13] != ele[8][22];
    ele[8][13] != ele[8][23];
    ele[8][13] != ele[8][24];
    ele[8][13] != ele[8][25];
    ele[8][13] != ele[8][26];
    ele[8][13] != ele[8][27];
    ele[8][13] != ele[8][28];
    ele[8][13] != ele[8][29];
    ele[8][13] != ele[8][30];
    ele[8][13] != ele[8][31];
    ele[8][13] != ele[8][32];
    ele[8][13] != ele[8][33];
    ele[8][13] != ele[8][34];
    ele[8][13] != ele[8][35];
    ele[8][13] != ele[9][12];
    ele[8][13] != ele[9][13];
    ele[8][13] != ele[9][14];
    ele[8][13] != ele[9][15];
    ele[8][13] != ele[9][16];
    ele[8][13] != ele[9][17];
    ele[8][14] != ele[10][12];
    ele[8][14] != ele[10][13];
    ele[8][14] != ele[10][14];
    ele[8][14] != ele[10][15];
    ele[8][14] != ele[10][16];
    ele[8][14] != ele[10][17];
    ele[8][14] != ele[11][12];
    ele[8][14] != ele[11][13];
    ele[8][14] != ele[11][14];
    ele[8][14] != ele[11][15];
    ele[8][14] != ele[11][16];
    ele[8][14] != ele[11][17];
    ele[8][14] != ele[12][14];
    ele[8][14] != ele[13][14];
    ele[8][14] != ele[14][14];
    ele[8][14] != ele[15][14];
    ele[8][14] != ele[16][14];
    ele[8][14] != ele[17][14];
    ele[8][14] != ele[18][14];
    ele[8][14] != ele[19][14];
    ele[8][14] != ele[20][14];
    ele[8][14] != ele[21][14];
    ele[8][14] != ele[22][14];
    ele[8][14] != ele[23][14];
    ele[8][14] != ele[24][14];
    ele[8][14] != ele[25][14];
    ele[8][14] != ele[26][14];
    ele[8][14] != ele[27][14];
    ele[8][14] != ele[28][14];
    ele[8][14] != ele[29][14];
    ele[8][14] != ele[30][14];
    ele[8][14] != ele[31][14];
    ele[8][14] != ele[32][14];
    ele[8][14] != ele[33][14];
    ele[8][14] != ele[34][14];
    ele[8][14] != ele[35][14];
    ele[8][14] != ele[8][15];
    ele[8][14] != ele[8][16];
    ele[8][14] != ele[8][17];
    ele[8][14] != ele[8][18];
    ele[8][14] != ele[8][19];
    ele[8][14] != ele[8][20];
    ele[8][14] != ele[8][21];
    ele[8][14] != ele[8][22];
    ele[8][14] != ele[8][23];
    ele[8][14] != ele[8][24];
    ele[8][14] != ele[8][25];
    ele[8][14] != ele[8][26];
    ele[8][14] != ele[8][27];
    ele[8][14] != ele[8][28];
    ele[8][14] != ele[8][29];
    ele[8][14] != ele[8][30];
    ele[8][14] != ele[8][31];
    ele[8][14] != ele[8][32];
    ele[8][14] != ele[8][33];
    ele[8][14] != ele[8][34];
    ele[8][14] != ele[8][35];
    ele[8][14] != ele[9][12];
    ele[8][14] != ele[9][13];
    ele[8][14] != ele[9][14];
    ele[8][14] != ele[9][15];
    ele[8][14] != ele[9][16];
    ele[8][14] != ele[9][17];
    ele[8][15] != ele[10][12];
    ele[8][15] != ele[10][13];
    ele[8][15] != ele[10][14];
    ele[8][15] != ele[10][15];
    ele[8][15] != ele[10][16];
    ele[8][15] != ele[10][17];
    ele[8][15] != ele[11][12];
    ele[8][15] != ele[11][13];
    ele[8][15] != ele[11][14];
    ele[8][15] != ele[11][15];
    ele[8][15] != ele[11][16];
    ele[8][15] != ele[11][17];
    ele[8][15] != ele[12][15];
    ele[8][15] != ele[13][15];
    ele[8][15] != ele[14][15];
    ele[8][15] != ele[15][15];
    ele[8][15] != ele[16][15];
    ele[8][15] != ele[17][15];
    ele[8][15] != ele[18][15];
    ele[8][15] != ele[19][15];
    ele[8][15] != ele[20][15];
    ele[8][15] != ele[21][15];
    ele[8][15] != ele[22][15];
    ele[8][15] != ele[23][15];
    ele[8][15] != ele[24][15];
    ele[8][15] != ele[25][15];
    ele[8][15] != ele[26][15];
    ele[8][15] != ele[27][15];
    ele[8][15] != ele[28][15];
    ele[8][15] != ele[29][15];
    ele[8][15] != ele[30][15];
    ele[8][15] != ele[31][15];
    ele[8][15] != ele[32][15];
    ele[8][15] != ele[33][15];
    ele[8][15] != ele[34][15];
    ele[8][15] != ele[35][15];
    ele[8][15] != ele[8][16];
    ele[8][15] != ele[8][17];
    ele[8][15] != ele[8][18];
    ele[8][15] != ele[8][19];
    ele[8][15] != ele[8][20];
    ele[8][15] != ele[8][21];
    ele[8][15] != ele[8][22];
    ele[8][15] != ele[8][23];
    ele[8][15] != ele[8][24];
    ele[8][15] != ele[8][25];
    ele[8][15] != ele[8][26];
    ele[8][15] != ele[8][27];
    ele[8][15] != ele[8][28];
    ele[8][15] != ele[8][29];
    ele[8][15] != ele[8][30];
    ele[8][15] != ele[8][31];
    ele[8][15] != ele[8][32];
    ele[8][15] != ele[8][33];
    ele[8][15] != ele[8][34];
    ele[8][15] != ele[8][35];
    ele[8][15] != ele[9][12];
    ele[8][15] != ele[9][13];
    ele[8][15] != ele[9][14];
    ele[8][15] != ele[9][15];
    ele[8][15] != ele[9][16];
    ele[8][15] != ele[9][17];
    ele[8][16] != ele[10][12];
    ele[8][16] != ele[10][13];
    ele[8][16] != ele[10][14];
    ele[8][16] != ele[10][15];
    ele[8][16] != ele[10][16];
    ele[8][16] != ele[10][17];
    ele[8][16] != ele[11][12];
    ele[8][16] != ele[11][13];
    ele[8][16] != ele[11][14];
    ele[8][16] != ele[11][15];
    ele[8][16] != ele[11][16];
    ele[8][16] != ele[11][17];
    ele[8][16] != ele[12][16];
    ele[8][16] != ele[13][16];
    ele[8][16] != ele[14][16];
    ele[8][16] != ele[15][16];
    ele[8][16] != ele[16][16];
    ele[8][16] != ele[17][16];
    ele[8][16] != ele[18][16];
    ele[8][16] != ele[19][16];
    ele[8][16] != ele[20][16];
    ele[8][16] != ele[21][16];
    ele[8][16] != ele[22][16];
    ele[8][16] != ele[23][16];
    ele[8][16] != ele[24][16];
    ele[8][16] != ele[25][16];
    ele[8][16] != ele[26][16];
    ele[8][16] != ele[27][16];
    ele[8][16] != ele[28][16];
    ele[8][16] != ele[29][16];
    ele[8][16] != ele[30][16];
    ele[8][16] != ele[31][16];
    ele[8][16] != ele[32][16];
    ele[8][16] != ele[33][16];
    ele[8][16] != ele[34][16];
    ele[8][16] != ele[35][16];
    ele[8][16] != ele[8][17];
    ele[8][16] != ele[8][18];
    ele[8][16] != ele[8][19];
    ele[8][16] != ele[8][20];
    ele[8][16] != ele[8][21];
    ele[8][16] != ele[8][22];
    ele[8][16] != ele[8][23];
    ele[8][16] != ele[8][24];
    ele[8][16] != ele[8][25];
    ele[8][16] != ele[8][26];
    ele[8][16] != ele[8][27];
    ele[8][16] != ele[8][28];
    ele[8][16] != ele[8][29];
    ele[8][16] != ele[8][30];
    ele[8][16] != ele[8][31];
    ele[8][16] != ele[8][32];
    ele[8][16] != ele[8][33];
    ele[8][16] != ele[8][34];
    ele[8][16] != ele[8][35];
    ele[8][16] != ele[9][12];
    ele[8][16] != ele[9][13];
    ele[8][16] != ele[9][14];
    ele[8][16] != ele[9][15];
    ele[8][16] != ele[9][16];
    ele[8][16] != ele[9][17];
    ele[8][17] != ele[10][12];
    ele[8][17] != ele[10][13];
    ele[8][17] != ele[10][14];
    ele[8][17] != ele[10][15];
    ele[8][17] != ele[10][16];
    ele[8][17] != ele[10][17];
    ele[8][17] != ele[11][12];
    ele[8][17] != ele[11][13];
    ele[8][17] != ele[11][14];
    ele[8][17] != ele[11][15];
    ele[8][17] != ele[11][16];
    ele[8][17] != ele[11][17];
    ele[8][17] != ele[12][17];
    ele[8][17] != ele[13][17];
    ele[8][17] != ele[14][17];
    ele[8][17] != ele[15][17];
    ele[8][17] != ele[16][17];
    ele[8][17] != ele[17][17];
    ele[8][17] != ele[18][17];
    ele[8][17] != ele[19][17];
    ele[8][17] != ele[20][17];
    ele[8][17] != ele[21][17];
    ele[8][17] != ele[22][17];
    ele[8][17] != ele[23][17];
    ele[8][17] != ele[24][17];
    ele[8][17] != ele[25][17];
    ele[8][17] != ele[26][17];
    ele[8][17] != ele[27][17];
    ele[8][17] != ele[28][17];
    ele[8][17] != ele[29][17];
    ele[8][17] != ele[30][17];
    ele[8][17] != ele[31][17];
    ele[8][17] != ele[32][17];
    ele[8][17] != ele[33][17];
    ele[8][17] != ele[34][17];
    ele[8][17] != ele[35][17];
    ele[8][17] != ele[8][18];
    ele[8][17] != ele[8][19];
    ele[8][17] != ele[8][20];
    ele[8][17] != ele[8][21];
    ele[8][17] != ele[8][22];
    ele[8][17] != ele[8][23];
    ele[8][17] != ele[8][24];
    ele[8][17] != ele[8][25];
    ele[8][17] != ele[8][26];
    ele[8][17] != ele[8][27];
    ele[8][17] != ele[8][28];
    ele[8][17] != ele[8][29];
    ele[8][17] != ele[8][30];
    ele[8][17] != ele[8][31];
    ele[8][17] != ele[8][32];
    ele[8][17] != ele[8][33];
    ele[8][17] != ele[8][34];
    ele[8][17] != ele[8][35];
    ele[8][17] != ele[9][12];
    ele[8][17] != ele[9][13];
    ele[8][17] != ele[9][14];
    ele[8][17] != ele[9][15];
    ele[8][17] != ele[9][16];
    ele[8][17] != ele[9][17];
    ele[8][18] != ele[10][18];
    ele[8][18] != ele[10][19];
    ele[8][18] != ele[10][20];
    ele[8][18] != ele[10][21];
    ele[8][18] != ele[10][22];
    ele[8][18] != ele[10][23];
    ele[8][18] != ele[11][18];
    ele[8][18] != ele[11][19];
    ele[8][18] != ele[11][20];
    ele[8][18] != ele[11][21];
    ele[8][18] != ele[11][22];
    ele[8][18] != ele[11][23];
    ele[8][18] != ele[12][18];
    ele[8][18] != ele[13][18];
    ele[8][18] != ele[14][18];
    ele[8][18] != ele[15][18];
    ele[8][18] != ele[16][18];
    ele[8][18] != ele[17][18];
    ele[8][18] != ele[18][18];
    ele[8][18] != ele[19][18];
    ele[8][18] != ele[20][18];
    ele[8][18] != ele[21][18];
    ele[8][18] != ele[22][18];
    ele[8][18] != ele[23][18];
    ele[8][18] != ele[24][18];
    ele[8][18] != ele[25][18];
    ele[8][18] != ele[26][18];
    ele[8][18] != ele[27][18];
    ele[8][18] != ele[28][18];
    ele[8][18] != ele[29][18];
    ele[8][18] != ele[30][18];
    ele[8][18] != ele[31][18];
    ele[8][18] != ele[32][18];
    ele[8][18] != ele[33][18];
    ele[8][18] != ele[34][18];
    ele[8][18] != ele[35][18];
    ele[8][18] != ele[8][19];
    ele[8][18] != ele[8][20];
    ele[8][18] != ele[8][21];
    ele[8][18] != ele[8][22];
    ele[8][18] != ele[8][23];
    ele[8][18] != ele[8][24];
    ele[8][18] != ele[8][25];
    ele[8][18] != ele[8][26];
    ele[8][18] != ele[8][27];
    ele[8][18] != ele[8][28];
    ele[8][18] != ele[8][29];
    ele[8][18] != ele[8][30];
    ele[8][18] != ele[8][31];
    ele[8][18] != ele[8][32];
    ele[8][18] != ele[8][33];
    ele[8][18] != ele[8][34];
    ele[8][18] != ele[8][35];
    ele[8][18] != ele[9][18];
    ele[8][18] != ele[9][19];
    ele[8][18] != ele[9][20];
    ele[8][18] != ele[9][21];
    ele[8][18] != ele[9][22];
    ele[8][18] != ele[9][23];
    ele[8][19] != ele[10][18];
    ele[8][19] != ele[10][19];
    ele[8][19] != ele[10][20];
    ele[8][19] != ele[10][21];
    ele[8][19] != ele[10][22];
    ele[8][19] != ele[10][23];
    ele[8][19] != ele[11][18];
    ele[8][19] != ele[11][19];
    ele[8][19] != ele[11][20];
    ele[8][19] != ele[11][21];
    ele[8][19] != ele[11][22];
    ele[8][19] != ele[11][23];
    ele[8][19] != ele[12][19];
    ele[8][19] != ele[13][19];
    ele[8][19] != ele[14][19];
    ele[8][19] != ele[15][19];
    ele[8][19] != ele[16][19];
    ele[8][19] != ele[17][19];
    ele[8][19] != ele[18][19];
    ele[8][19] != ele[19][19];
    ele[8][19] != ele[20][19];
    ele[8][19] != ele[21][19];
    ele[8][19] != ele[22][19];
    ele[8][19] != ele[23][19];
    ele[8][19] != ele[24][19];
    ele[8][19] != ele[25][19];
    ele[8][19] != ele[26][19];
    ele[8][19] != ele[27][19];
    ele[8][19] != ele[28][19];
    ele[8][19] != ele[29][19];
    ele[8][19] != ele[30][19];
    ele[8][19] != ele[31][19];
    ele[8][19] != ele[32][19];
    ele[8][19] != ele[33][19];
    ele[8][19] != ele[34][19];
    ele[8][19] != ele[35][19];
    ele[8][19] != ele[8][20];
    ele[8][19] != ele[8][21];
    ele[8][19] != ele[8][22];
    ele[8][19] != ele[8][23];
    ele[8][19] != ele[8][24];
    ele[8][19] != ele[8][25];
    ele[8][19] != ele[8][26];
    ele[8][19] != ele[8][27];
    ele[8][19] != ele[8][28];
    ele[8][19] != ele[8][29];
    ele[8][19] != ele[8][30];
    ele[8][19] != ele[8][31];
    ele[8][19] != ele[8][32];
    ele[8][19] != ele[8][33];
    ele[8][19] != ele[8][34];
    ele[8][19] != ele[8][35];
    ele[8][19] != ele[9][18];
    ele[8][19] != ele[9][19];
    ele[8][19] != ele[9][20];
    ele[8][19] != ele[9][21];
    ele[8][19] != ele[9][22];
    ele[8][19] != ele[9][23];
    ele[8][2] != ele[10][0];
    ele[8][2] != ele[10][1];
    ele[8][2] != ele[10][2];
    ele[8][2] != ele[10][3];
    ele[8][2] != ele[10][4];
    ele[8][2] != ele[10][5];
    ele[8][2] != ele[11][0];
    ele[8][2] != ele[11][1];
    ele[8][2] != ele[11][2];
    ele[8][2] != ele[11][3];
    ele[8][2] != ele[11][4];
    ele[8][2] != ele[11][5];
    ele[8][2] != ele[12][2];
    ele[8][2] != ele[13][2];
    ele[8][2] != ele[14][2];
    ele[8][2] != ele[15][2];
    ele[8][2] != ele[16][2];
    ele[8][2] != ele[17][2];
    ele[8][2] != ele[18][2];
    ele[8][2] != ele[19][2];
    ele[8][2] != ele[20][2];
    ele[8][2] != ele[21][2];
    ele[8][2] != ele[22][2];
    ele[8][2] != ele[23][2];
    ele[8][2] != ele[24][2];
    ele[8][2] != ele[25][2];
    ele[8][2] != ele[26][2];
    ele[8][2] != ele[27][2];
    ele[8][2] != ele[28][2];
    ele[8][2] != ele[29][2];
    ele[8][2] != ele[30][2];
    ele[8][2] != ele[31][2];
    ele[8][2] != ele[32][2];
    ele[8][2] != ele[33][2];
    ele[8][2] != ele[34][2];
    ele[8][2] != ele[35][2];
    ele[8][2] != ele[8][10];
    ele[8][2] != ele[8][11];
    ele[8][2] != ele[8][12];
    ele[8][2] != ele[8][13];
    ele[8][2] != ele[8][14];
    ele[8][2] != ele[8][15];
    ele[8][2] != ele[8][16];
    ele[8][2] != ele[8][17];
    ele[8][2] != ele[8][18];
    ele[8][2] != ele[8][19];
    ele[8][2] != ele[8][20];
    ele[8][2] != ele[8][21];
    ele[8][2] != ele[8][22];
    ele[8][2] != ele[8][23];
    ele[8][2] != ele[8][24];
    ele[8][2] != ele[8][25];
    ele[8][2] != ele[8][26];
    ele[8][2] != ele[8][27];
    ele[8][2] != ele[8][28];
    ele[8][2] != ele[8][29];
    ele[8][2] != ele[8][3];
    ele[8][2] != ele[8][30];
    ele[8][2] != ele[8][31];
    ele[8][2] != ele[8][32];
    ele[8][2] != ele[8][33];
    ele[8][2] != ele[8][34];
    ele[8][2] != ele[8][35];
    ele[8][2] != ele[8][4];
    ele[8][2] != ele[8][5];
    ele[8][2] != ele[8][6];
    ele[8][2] != ele[8][7];
    ele[8][2] != ele[8][8];
    ele[8][2] != ele[8][9];
    ele[8][2] != ele[9][0];
    ele[8][2] != ele[9][1];
    ele[8][2] != ele[9][2];
    ele[8][2] != ele[9][3];
    ele[8][2] != ele[9][4];
    ele[8][2] != ele[9][5];
    ele[8][20] != ele[10][18];
    ele[8][20] != ele[10][19];
    ele[8][20] != ele[10][20];
    ele[8][20] != ele[10][21];
    ele[8][20] != ele[10][22];
    ele[8][20] != ele[10][23];
    ele[8][20] != ele[11][18];
    ele[8][20] != ele[11][19];
    ele[8][20] != ele[11][20];
    ele[8][20] != ele[11][21];
    ele[8][20] != ele[11][22];
    ele[8][20] != ele[11][23];
    ele[8][20] != ele[12][20];
    ele[8][20] != ele[13][20];
    ele[8][20] != ele[14][20];
    ele[8][20] != ele[15][20];
    ele[8][20] != ele[16][20];
    ele[8][20] != ele[17][20];
    ele[8][20] != ele[18][20];
    ele[8][20] != ele[19][20];
    ele[8][20] != ele[20][20];
    ele[8][20] != ele[21][20];
    ele[8][20] != ele[22][20];
    ele[8][20] != ele[23][20];
    ele[8][20] != ele[24][20];
    ele[8][20] != ele[25][20];
    ele[8][20] != ele[26][20];
    ele[8][20] != ele[27][20];
    ele[8][20] != ele[28][20];
    ele[8][20] != ele[29][20];
    ele[8][20] != ele[30][20];
    ele[8][20] != ele[31][20];
    ele[8][20] != ele[32][20];
    ele[8][20] != ele[33][20];
    ele[8][20] != ele[34][20];
    ele[8][20] != ele[35][20];
    ele[8][20] != ele[8][21];
    ele[8][20] != ele[8][22];
    ele[8][20] != ele[8][23];
    ele[8][20] != ele[8][24];
    ele[8][20] != ele[8][25];
    ele[8][20] != ele[8][26];
    ele[8][20] != ele[8][27];
    ele[8][20] != ele[8][28];
    ele[8][20] != ele[8][29];
    ele[8][20] != ele[8][30];
    ele[8][20] != ele[8][31];
    ele[8][20] != ele[8][32];
    ele[8][20] != ele[8][33];
    ele[8][20] != ele[8][34];
    ele[8][20] != ele[8][35];
    ele[8][20] != ele[9][18];
    ele[8][20] != ele[9][19];
    ele[8][20] != ele[9][20];
    ele[8][20] != ele[9][21];
    ele[8][20] != ele[9][22];
    ele[8][20] != ele[9][23];
    ele[8][21] != ele[10][18];
    ele[8][21] != ele[10][19];
    ele[8][21] != ele[10][20];
    ele[8][21] != ele[10][21];
    ele[8][21] != ele[10][22];
    ele[8][21] != ele[10][23];
    ele[8][21] != ele[11][18];
    ele[8][21] != ele[11][19];
    ele[8][21] != ele[11][20];
    ele[8][21] != ele[11][21];
    ele[8][21] != ele[11][22];
    ele[8][21] != ele[11][23];
    ele[8][21] != ele[12][21];
    ele[8][21] != ele[13][21];
    ele[8][21] != ele[14][21];
    ele[8][21] != ele[15][21];
    ele[8][21] != ele[16][21];
    ele[8][21] != ele[17][21];
    ele[8][21] != ele[18][21];
    ele[8][21] != ele[19][21];
    ele[8][21] != ele[20][21];
    ele[8][21] != ele[21][21];
    ele[8][21] != ele[22][21];
    ele[8][21] != ele[23][21];
    ele[8][21] != ele[24][21];
    ele[8][21] != ele[25][21];
    ele[8][21] != ele[26][21];
    ele[8][21] != ele[27][21];
    ele[8][21] != ele[28][21];
    ele[8][21] != ele[29][21];
    ele[8][21] != ele[30][21];
    ele[8][21] != ele[31][21];
    ele[8][21] != ele[32][21];
    ele[8][21] != ele[33][21];
    ele[8][21] != ele[34][21];
    ele[8][21] != ele[35][21];
    ele[8][21] != ele[8][22];
    ele[8][21] != ele[8][23];
    ele[8][21] != ele[8][24];
    ele[8][21] != ele[8][25];
    ele[8][21] != ele[8][26];
    ele[8][21] != ele[8][27];
    ele[8][21] != ele[8][28];
    ele[8][21] != ele[8][29];
    ele[8][21] != ele[8][30];
    ele[8][21] != ele[8][31];
    ele[8][21] != ele[8][32];
    ele[8][21] != ele[8][33];
    ele[8][21] != ele[8][34];
    ele[8][21] != ele[8][35];
    ele[8][21] != ele[9][18];
    ele[8][21] != ele[9][19];
    ele[8][21] != ele[9][20];
    ele[8][21] != ele[9][21];
    ele[8][21] != ele[9][22];
    ele[8][21] != ele[9][23];
    ele[8][22] != ele[10][18];
    ele[8][22] != ele[10][19];
    ele[8][22] != ele[10][20];
    ele[8][22] != ele[10][21];
    ele[8][22] != ele[10][22];
    ele[8][22] != ele[10][23];
    ele[8][22] != ele[11][18];
    ele[8][22] != ele[11][19];
    ele[8][22] != ele[11][20];
    ele[8][22] != ele[11][21];
    ele[8][22] != ele[11][22];
    ele[8][22] != ele[11][23];
    ele[8][22] != ele[12][22];
    ele[8][22] != ele[13][22];
    ele[8][22] != ele[14][22];
    ele[8][22] != ele[15][22];
    ele[8][22] != ele[16][22];
    ele[8][22] != ele[17][22];
    ele[8][22] != ele[18][22];
    ele[8][22] != ele[19][22];
    ele[8][22] != ele[20][22];
    ele[8][22] != ele[21][22];
    ele[8][22] != ele[22][22];
    ele[8][22] != ele[23][22];
    ele[8][22] != ele[24][22];
    ele[8][22] != ele[25][22];
    ele[8][22] != ele[26][22];
    ele[8][22] != ele[27][22];
    ele[8][22] != ele[28][22];
    ele[8][22] != ele[29][22];
    ele[8][22] != ele[30][22];
    ele[8][22] != ele[31][22];
    ele[8][22] != ele[32][22];
    ele[8][22] != ele[33][22];
    ele[8][22] != ele[34][22];
    ele[8][22] != ele[35][22];
    ele[8][22] != ele[8][23];
    ele[8][22] != ele[8][24];
    ele[8][22] != ele[8][25];
    ele[8][22] != ele[8][26];
    ele[8][22] != ele[8][27];
    ele[8][22] != ele[8][28];
    ele[8][22] != ele[8][29];
    ele[8][22] != ele[8][30];
    ele[8][22] != ele[8][31];
    ele[8][22] != ele[8][32];
    ele[8][22] != ele[8][33];
    ele[8][22] != ele[8][34];
    ele[8][22] != ele[8][35];
    ele[8][22] != ele[9][18];
    ele[8][22] != ele[9][19];
    ele[8][22] != ele[9][20];
    ele[8][22] != ele[9][21];
    ele[8][22] != ele[9][22];
    ele[8][22] != ele[9][23];
    ele[8][23] != ele[10][18];
    ele[8][23] != ele[10][19];
    ele[8][23] != ele[10][20];
    ele[8][23] != ele[10][21];
    ele[8][23] != ele[10][22];
    ele[8][23] != ele[10][23];
    ele[8][23] != ele[11][18];
    ele[8][23] != ele[11][19];
    ele[8][23] != ele[11][20];
    ele[8][23] != ele[11][21];
    ele[8][23] != ele[11][22];
    ele[8][23] != ele[11][23];
    ele[8][23] != ele[12][23];
    ele[8][23] != ele[13][23];
    ele[8][23] != ele[14][23];
    ele[8][23] != ele[15][23];
    ele[8][23] != ele[16][23];
    ele[8][23] != ele[17][23];
    ele[8][23] != ele[18][23];
    ele[8][23] != ele[19][23];
    ele[8][23] != ele[20][23];
    ele[8][23] != ele[21][23];
    ele[8][23] != ele[22][23];
    ele[8][23] != ele[23][23];
    ele[8][23] != ele[24][23];
    ele[8][23] != ele[25][23];
    ele[8][23] != ele[26][23];
    ele[8][23] != ele[27][23];
    ele[8][23] != ele[28][23];
    ele[8][23] != ele[29][23];
    ele[8][23] != ele[30][23];
    ele[8][23] != ele[31][23];
    ele[8][23] != ele[32][23];
    ele[8][23] != ele[33][23];
    ele[8][23] != ele[34][23];
    ele[8][23] != ele[35][23];
    ele[8][23] != ele[8][24];
    ele[8][23] != ele[8][25];
    ele[8][23] != ele[8][26];
    ele[8][23] != ele[8][27];
    ele[8][23] != ele[8][28];
    ele[8][23] != ele[8][29];
    ele[8][23] != ele[8][30];
    ele[8][23] != ele[8][31];
    ele[8][23] != ele[8][32];
    ele[8][23] != ele[8][33];
    ele[8][23] != ele[8][34];
    ele[8][23] != ele[8][35];
    ele[8][23] != ele[9][18];
    ele[8][23] != ele[9][19];
    ele[8][23] != ele[9][20];
    ele[8][23] != ele[9][21];
    ele[8][23] != ele[9][22];
    ele[8][23] != ele[9][23];
    ele[8][24] != ele[10][24];
    ele[8][24] != ele[10][25];
    ele[8][24] != ele[10][26];
    ele[8][24] != ele[10][27];
    ele[8][24] != ele[10][28];
    ele[8][24] != ele[10][29];
    ele[8][24] != ele[11][24];
    ele[8][24] != ele[11][25];
    ele[8][24] != ele[11][26];
    ele[8][24] != ele[11][27];
    ele[8][24] != ele[11][28];
    ele[8][24] != ele[11][29];
    ele[8][24] != ele[12][24];
    ele[8][24] != ele[13][24];
    ele[8][24] != ele[14][24];
    ele[8][24] != ele[15][24];
    ele[8][24] != ele[16][24];
    ele[8][24] != ele[17][24];
    ele[8][24] != ele[18][24];
    ele[8][24] != ele[19][24];
    ele[8][24] != ele[20][24];
    ele[8][24] != ele[21][24];
    ele[8][24] != ele[22][24];
    ele[8][24] != ele[23][24];
    ele[8][24] != ele[24][24];
    ele[8][24] != ele[25][24];
    ele[8][24] != ele[26][24];
    ele[8][24] != ele[27][24];
    ele[8][24] != ele[28][24];
    ele[8][24] != ele[29][24];
    ele[8][24] != ele[30][24];
    ele[8][24] != ele[31][24];
    ele[8][24] != ele[32][24];
    ele[8][24] != ele[33][24];
    ele[8][24] != ele[34][24];
    ele[8][24] != ele[35][24];
    ele[8][24] != ele[8][25];
    ele[8][24] != ele[8][26];
    ele[8][24] != ele[8][27];
    ele[8][24] != ele[8][28];
    ele[8][24] != ele[8][29];
    ele[8][24] != ele[8][30];
    ele[8][24] != ele[8][31];
    ele[8][24] != ele[8][32];
    ele[8][24] != ele[8][33];
    ele[8][24] != ele[8][34];
    ele[8][24] != ele[8][35];
    ele[8][24] != ele[9][24];
    ele[8][24] != ele[9][25];
    ele[8][24] != ele[9][26];
    ele[8][24] != ele[9][27];
    ele[8][24] != ele[9][28];
    ele[8][24] != ele[9][29];
    ele[8][25] != ele[10][24];
    ele[8][25] != ele[10][25];
    ele[8][25] != ele[10][26];
    ele[8][25] != ele[10][27];
    ele[8][25] != ele[10][28];
    ele[8][25] != ele[10][29];
    ele[8][25] != ele[11][24];
    ele[8][25] != ele[11][25];
    ele[8][25] != ele[11][26];
    ele[8][25] != ele[11][27];
    ele[8][25] != ele[11][28];
    ele[8][25] != ele[11][29];
    ele[8][25] != ele[12][25];
    ele[8][25] != ele[13][25];
    ele[8][25] != ele[14][25];
    ele[8][25] != ele[15][25];
    ele[8][25] != ele[16][25];
    ele[8][25] != ele[17][25];
    ele[8][25] != ele[18][25];
    ele[8][25] != ele[19][25];
    ele[8][25] != ele[20][25];
    ele[8][25] != ele[21][25];
    ele[8][25] != ele[22][25];
    ele[8][25] != ele[23][25];
    ele[8][25] != ele[24][25];
    ele[8][25] != ele[25][25];
    ele[8][25] != ele[26][25];
    ele[8][25] != ele[27][25];
    ele[8][25] != ele[28][25];
    ele[8][25] != ele[29][25];
    ele[8][25] != ele[30][25];
    ele[8][25] != ele[31][25];
    ele[8][25] != ele[32][25];
    ele[8][25] != ele[33][25];
    ele[8][25] != ele[34][25];
    ele[8][25] != ele[35][25];
    ele[8][25] != ele[8][26];
    ele[8][25] != ele[8][27];
    ele[8][25] != ele[8][28];
    ele[8][25] != ele[8][29];
    ele[8][25] != ele[8][30];
    ele[8][25] != ele[8][31];
    ele[8][25] != ele[8][32];
    ele[8][25] != ele[8][33];
    ele[8][25] != ele[8][34];
    ele[8][25] != ele[8][35];
    ele[8][25] != ele[9][24];
    ele[8][25] != ele[9][25];
    ele[8][25] != ele[9][26];
    ele[8][25] != ele[9][27];
    ele[8][25] != ele[9][28];
    ele[8][25] != ele[9][29];
    ele[8][26] != ele[10][24];
    ele[8][26] != ele[10][25];
    ele[8][26] != ele[10][26];
    ele[8][26] != ele[10][27];
    ele[8][26] != ele[10][28];
    ele[8][26] != ele[10][29];
    ele[8][26] != ele[11][24];
    ele[8][26] != ele[11][25];
    ele[8][26] != ele[11][26];
    ele[8][26] != ele[11][27];
    ele[8][26] != ele[11][28];
    ele[8][26] != ele[11][29];
    ele[8][26] != ele[12][26];
    ele[8][26] != ele[13][26];
    ele[8][26] != ele[14][26];
    ele[8][26] != ele[15][26];
    ele[8][26] != ele[16][26];
    ele[8][26] != ele[17][26];
    ele[8][26] != ele[18][26];
    ele[8][26] != ele[19][26];
    ele[8][26] != ele[20][26];
    ele[8][26] != ele[21][26];
    ele[8][26] != ele[22][26];
    ele[8][26] != ele[23][26];
    ele[8][26] != ele[24][26];
    ele[8][26] != ele[25][26];
    ele[8][26] != ele[26][26];
    ele[8][26] != ele[27][26];
    ele[8][26] != ele[28][26];
    ele[8][26] != ele[29][26];
    ele[8][26] != ele[30][26];
    ele[8][26] != ele[31][26];
    ele[8][26] != ele[32][26];
    ele[8][26] != ele[33][26];
    ele[8][26] != ele[34][26];
    ele[8][26] != ele[35][26];
    ele[8][26] != ele[8][27];
    ele[8][26] != ele[8][28];
    ele[8][26] != ele[8][29];
    ele[8][26] != ele[8][30];
    ele[8][26] != ele[8][31];
    ele[8][26] != ele[8][32];
    ele[8][26] != ele[8][33];
    ele[8][26] != ele[8][34];
    ele[8][26] != ele[8][35];
    ele[8][26] != ele[9][24];
    ele[8][26] != ele[9][25];
    ele[8][26] != ele[9][26];
    ele[8][26] != ele[9][27];
    ele[8][26] != ele[9][28];
    ele[8][26] != ele[9][29];
    ele[8][27] != ele[10][24];
    ele[8][27] != ele[10][25];
    ele[8][27] != ele[10][26];
    ele[8][27] != ele[10][27];
    ele[8][27] != ele[10][28];
    ele[8][27] != ele[10][29];
    ele[8][27] != ele[11][24];
    ele[8][27] != ele[11][25];
    ele[8][27] != ele[11][26];
    ele[8][27] != ele[11][27];
    ele[8][27] != ele[11][28];
    ele[8][27] != ele[11][29];
    ele[8][27] != ele[12][27];
    ele[8][27] != ele[13][27];
    ele[8][27] != ele[14][27];
    ele[8][27] != ele[15][27];
    ele[8][27] != ele[16][27];
    ele[8][27] != ele[17][27];
    ele[8][27] != ele[18][27];
    ele[8][27] != ele[19][27];
    ele[8][27] != ele[20][27];
    ele[8][27] != ele[21][27];
    ele[8][27] != ele[22][27];
    ele[8][27] != ele[23][27];
    ele[8][27] != ele[24][27];
    ele[8][27] != ele[25][27];
    ele[8][27] != ele[26][27];
    ele[8][27] != ele[27][27];
    ele[8][27] != ele[28][27];
    ele[8][27] != ele[29][27];
    ele[8][27] != ele[30][27];
    ele[8][27] != ele[31][27];
    ele[8][27] != ele[32][27];
    ele[8][27] != ele[33][27];
    ele[8][27] != ele[34][27];
    ele[8][27] != ele[35][27];
    ele[8][27] != ele[8][28];
    ele[8][27] != ele[8][29];
    ele[8][27] != ele[8][30];
    ele[8][27] != ele[8][31];
    ele[8][27] != ele[8][32];
    ele[8][27] != ele[8][33];
    ele[8][27] != ele[8][34];
    ele[8][27] != ele[8][35];
    ele[8][27] != ele[9][24];
    ele[8][27] != ele[9][25];
    ele[8][27] != ele[9][26];
    ele[8][27] != ele[9][27];
    ele[8][27] != ele[9][28];
    ele[8][27] != ele[9][29];
    ele[8][28] != ele[10][24];
    ele[8][28] != ele[10][25];
    ele[8][28] != ele[10][26];
    ele[8][28] != ele[10][27];
    ele[8][28] != ele[10][28];
    ele[8][28] != ele[10][29];
    ele[8][28] != ele[11][24];
    ele[8][28] != ele[11][25];
    ele[8][28] != ele[11][26];
    ele[8][28] != ele[11][27];
    ele[8][28] != ele[11][28];
    ele[8][28] != ele[11][29];
    ele[8][28] != ele[12][28];
    ele[8][28] != ele[13][28];
    ele[8][28] != ele[14][28];
    ele[8][28] != ele[15][28];
    ele[8][28] != ele[16][28];
    ele[8][28] != ele[17][28];
    ele[8][28] != ele[18][28];
    ele[8][28] != ele[19][28];
    ele[8][28] != ele[20][28];
    ele[8][28] != ele[21][28];
    ele[8][28] != ele[22][28];
    ele[8][28] != ele[23][28];
    ele[8][28] != ele[24][28];
    ele[8][28] != ele[25][28];
    ele[8][28] != ele[26][28];
    ele[8][28] != ele[27][28];
    ele[8][28] != ele[28][28];
    ele[8][28] != ele[29][28];
    ele[8][28] != ele[30][28];
    ele[8][28] != ele[31][28];
    ele[8][28] != ele[32][28];
    ele[8][28] != ele[33][28];
    ele[8][28] != ele[34][28];
    ele[8][28] != ele[35][28];
    ele[8][28] != ele[8][29];
    ele[8][28] != ele[8][30];
    ele[8][28] != ele[8][31];
    ele[8][28] != ele[8][32];
    ele[8][28] != ele[8][33];
    ele[8][28] != ele[8][34];
    ele[8][28] != ele[8][35];
    ele[8][28] != ele[9][24];
    ele[8][28] != ele[9][25];
    ele[8][28] != ele[9][26];
    ele[8][28] != ele[9][27];
    ele[8][28] != ele[9][28];
    ele[8][28] != ele[9][29];
    ele[8][29] != ele[10][24];
    ele[8][29] != ele[10][25];
    ele[8][29] != ele[10][26];
    ele[8][29] != ele[10][27];
    ele[8][29] != ele[10][28];
    ele[8][29] != ele[10][29];
    ele[8][29] != ele[11][24];
    ele[8][29] != ele[11][25];
    ele[8][29] != ele[11][26];
    ele[8][29] != ele[11][27];
    ele[8][29] != ele[11][28];
    ele[8][29] != ele[11][29];
    ele[8][29] != ele[12][29];
    ele[8][29] != ele[13][29];
    ele[8][29] != ele[14][29];
    ele[8][29] != ele[15][29];
    ele[8][29] != ele[16][29];
    ele[8][29] != ele[17][29];
    ele[8][29] != ele[18][29];
    ele[8][29] != ele[19][29];
    ele[8][29] != ele[20][29];
    ele[8][29] != ele[21][29];
    ele[8][29] != ele[22][29];
    ele[8][29] != ele[23][29];
    ele[8][29] != ele[24][29];
    ele[8][29] != ele[25][29];
    ele[8][29] != ele[26][29];
    ele[8][29] != ele[27][29];
    ele[8][29] != ele[28][29];
    ele[8][29] != ele[29][29];
    ele[8][29] != ele[30][29];
    ele[8][29] != ele[31][29];
    ele[8][29] != ele[32][29];
    ele[8][29] != ele[33][29];
    ele[8][29] != ele[34][29];
    ele[8][29] != ele[35][29];
    ele[8][29] != ele[8][30];
    ele[8][29] != ele[8][31];
    ele[8][29] != ele[8][32];
    ele[8][29] != ele[8][33];
    ele[8][29] != ele[8][34];
    ele[8][29] != ele[8][35];
    ele[8][29] != ele[9][24];
    ele[8][29] != ele[9][25];
    ele[8][29] != ele[9][26];
    ele[8][29] != ele[9][27];
    ele[8][29] != ele[9][28];
    ele[8][29] != ele[9][29];
    ele[8][3] != ele[10][0];
    ele[8][3] != ele[10][1];
    ele[8][3] != ele[10][2];
    ele[8][3] != ele[10][3];
    ele[8][3] != ele[10][4];
    ele[8][3] != ele[10][5];
    ele[8][3] != ele[11][0];
    ele[8][3] != ele[11][1];
    ele[8][3] != ele[11][2];
    ele[8][3] != ele[11][3];
    ele[8][3] != ele[11][4];
    ele[8][3] != ele[11][5];
    ele[8][3] != ele[12][3];
    ele[8][3] != ele[13][3];
    ele[8][3] != ele[14][3];
    ele[8][3] != ele[15][3];
    ele[8][3] != ele[16][3];
    ele[8][3] != ele[17][3];
    ele[8][3] != ele[18][3];
    ele[8][3] != ele[19][3];
    ele[8][3] != ele[20][3];
    ele[8][3] != ele[21][3];
    ele[8][3] != ele[22][3];
    ele[8][3] != ele[23][3];
    ele[8][3] != ele[24][3];
    ele[8][3] != ele[25][3];
    ele[8][3] != ele[26][3];
    ele[8][3] != ele[27][3];
    ele[8][3] != ele[28][3];
    ele[8][3] != ele[29][3];
    ele[8][3] != ele[30][3];
    ele[8][3] != ele[31][3];
    ele[8][3] != ele[32][3];
    ele[8][3] != ele[33][3];
    ele[8][3] != ele[34][3];
    ele[8][3] != ele[35][3];
    ele[8][3] != ele[8][10];
    ele[8][3] != ele[8][11];
    ele[8][3] != ele[8][12];
    ele[8][3] != ele[8][13];
    ele[8][3] != ele[8][14];
    ele[8][3] != ele[8][15];
    ele[8][3] != ele[8][16];
    ele[8][3] != ele[8][17];
    ele[8][3] != ele[8][18];
    ele[8][3] != ele[8][19];
    ele[8][3] != ele[8][20];
    ele[8][3] != ele[8][21];
    ele[8][3] != ele[8][22];
    ele[8][3] != ele[8][23];
    ele[8][3] != ele[8][24];
    ele[8][3] != ele[8][25];
    ele[8][3] != ele[8][26];
    ele[8][3] != ele[8][27];
    ele[8][3] != ele[8][28];
    ele[8][3] != ele[8][29];
    ele[8][3] != ele[8][30];
    ele[8][3] != ele[8][31];
    ele[8][3] != ele[8][32];
    ele[8][3] != ele[8][33];
    ele[8][3] != ele[8][34];
    ele[8][3] != ele[8][35];
    ele[8][3] != ele[8][4];
    ele[8][3] != ele[8][5];
    ele[8][3] != ele[8][6];
    ele[8][3] != ele[8][7];
    ele[8][3] != ele[8][8];
    ele[8][3] != ele[8][9];
    ele[8][3] != ele[9][0];
    ele[8][3] != ele[9][1];
    ele[8][3] != ele[9][2];
    ele[8][3] != ele[9][3];
    ele[8][3] != ele[9][4];
    ele[8][3] != ele[9][5];
    ele[8][30] != ele[10][30];
    ele[8][30] != ele[10][31];
    ele[8][30] != ele[10][32];
    ele[8][30] != ele[10][33];
    ele[8][30] != ele[10][34];
    ele[8][30] != ele[10][35];
    ele[8][30] != ele[11][30];
    ele[8][30] != ele[11][31];
    ele[8][30] != ele[11][32];
    ele[8][30] != ele[11][33];
    ele[8][30] != ele[11][34];
    ele[8][30] != ele[11][35];
    ele[8][30] != ele[12][30];
    ele[8][30] != ele[13][30];
    ele[8][30] != ele[14][30];
    ele[8][30] != ele[15][30];
    ele[8][30] != ele[16][30];
    ele[8][30] != ele[17][30];
    ele[8][30] != ele[18][30];
    ele[8][30] != ele[19][30];
    ele[8][30] != ele[20][30];
    ele[8][30] != ele[21][30];
    ele[8][30] != ele[22][30];
    ele[8][30] != ele[23][30];
    ele[8][30] != ele[24][30];
    ele[8][30] != ele[25][30];
    ele[8][30] != ele[26][30];
    ele[8][30] != ele[27][30];
    ele[8][30] != ele[28][30];
    ele[8][30] != ele[29][30];
    ele[8][30] != ele[30][30];
    ele[8][30] != ele[31][30];
    ele[8][30] != ele[32][30];
    ele[8][30] != ele[33][30];
    ele[8][30] != ele[34][30];
    ele[8][30] != ele[35][30];
    ele[8][30] != ele[8][31];
    ele[8][30] != ele[8][32];
    ele[8][30] != ele[8][33];
    ele[8][30] != ele[8][34];
    ele[8][30] != ele[8][35];
    ele[8][30] != ele[9][30];
    ele[8][30] != ele[9][31];
    ele[8][30] != ele[9][32];
    ele[8][30] != ele[9][33];
    ele[8][30] != ele[9][34];
    ele[8][30] != ele[9][35];
    ele[8][31] != ele[10][30];
    ele[8][31] != ele[10][31];
    ele[8][31] != ele[10][32];
    ele[8][31] != ele[10][33];
    ele[8][31] != ele[10][34];
    ele[8][31] != ele[10][35];
    ele[8][31] != ele[11][30];
    ele[8][31] != ele[11][31];
    ele[8][31] != ele[11][32];
    ele[8][31] != ele[11][33];
    ele[8][31] != ele[11][34];
    ele[8][31] != ele[11][35];
    ele[8][31] != ele[12][31];
    ele[8][31] != ele[13][31];
    ele[8][31] != ele[14][31];
    ele[8][31] != ele[15][31];
    ele[8][31] != ele[16][31];
    ele[8][31] != ele[17][31];
    ele[8][31] != ele[18][31];
    ele[8][31] != ele[19][31];
    ele[8][31] != ele[20][31];
    ele[8][31] != ele[21][31];
    ele[8][31] != ele[22][31];
    ele[8][31] != ele[23][31];
    ele[8][31] != ele[24][31];
    ele[8][31] != ele[25][31];
    ele[8][31] != ele[26][31];
    ele[8][31] != ele[27][31];
    ele[8][31] != ele[28][31];
    ele[8][31] != ele[29][31];
    ele[8][31] != ele[30][31];
    ele[8][31] != ele[31][31];
    ele[8][31] != ele[32][31];
    ele[8][31] != ele[33][31];
    ele[8][31] != ele[34][31];
    ele[8][31] != ele[35][31];
    ele[8][31] != ele[8][32];
    ele[8][31] != ele[8][33];
    ele[8][31] != ele[8][34];
    ele[8][31] != ele[8][35];
    ele[8][31] != ele[9][30];
    ele[8][31] != ele[9][31];
    ele[8][31] != ele[9][32];
    ele[8][31] != ele[9][33];
    ele[8][31] != ele[9][34];
    ele[8][31] != ele[9][35];
    ele[8][32] != ele[10][30];
    ele[8][32] != ele[10][31];
    ele[8][32] != ele[10][32];
    ele[8][32] != ele[10][33];
    ele[8][32] != ele[10][34];
    ele[8][32] != ele[10][35];
    ele[8][32] != ele[11][30];
    ele[8][32] != ele[11][31];
    ele[8][32] != ele[11][32];
    ele[8][32] != ele[11][33];
    ele[8][32] != ele[11][34];
    ele[8][32] != ele[11][35];
    ele[8][32] != ele[12][32];
    ele[8][32] != ele[13][32];
    ele[8][32] != ele[14][32];
    ele[8][32] != ele[15][32];
    ele[8][32] != ele[16][32];
    ele[8][32] != ele[17][32];
    ele[8][32] != ele[18][32];
    ele[8][32] != ele[19][32];
    ele[8][32] != ele[20][32];
    ele[8][32] != ele[21][32];
    ele[8][32] != ele[22][32];
    ele[8][32] != ele[23][32];
    ele[8][32] != ele[24][32];
    ele[8][32] != ele[25][32];
    ele[8][32] != ele[26][32];
    ele[8][32] != ele[27][32];
    ele[8][32] != ele[28][32];
    ele[8][32] != ele[29][32];
    ele[8][32] != ele[30][32];
    ele[8][32] != ele[31][32];
    ele[8][32] != ele[32][32];
    ele[8][32] != ele[33][32];
    ele[8][32] != ele[34][32];
    ele[8][32] != ele[35][32];
    ele[8][32] != ele[8][33];
    ele[8][32] != ele[8][34];
    ele[8][32] != ele[8][35];
    ele[8][32] != ele[9][30];
    ele[8][32] != ele[9][31];
    ele[8][32] != ele[9][32];
    ele[8][32] != ele[9][33];
    ele[8][32] != ele[9][34];
    ele[8][32] != ele[9][35];
    ele[8][33] != ele[10][30];
    ele[8][33] != ele[10][31];
    ele[8][33] != ele[10][32];
    ele[8][33] != ele[10][33];
    ele[8][33] != ele[10][34];
    ele[8][33] != ele[10][35];
    ele[8][33] != ele[11][30];
    ele[8][33] != ele[11][31];
    ele[8][33] != ele[11][32];
    ele[8][33] != ele[11][33];
    ele[8][33] != ele[11][34];
    ele[8][33] != ele[11][35];
    ele[8][33] != ele[12][33];
    ele[8][33] != ele[13][33];
    ele[8][33] != ele[14][33];
    ele[8][33] != ele[15][33];
    ele[8][33] != ele[16][33];
    ele[8][33] != ele[17][33];
    ele[8][33] != ele[18][33];
    ele[8][33] != ele[19][33];
    ele[8][33] != ele[20][33];
    ele[8][33] != ele[21][33];
    ele[8][33] != ele[22][33];
    ele[8][33] != ele[23][33];
    ele[8][33] != ele[24][33];
    ele[8][33] != ele[25][33];
    ele[8][33] != ele[26][33];
    ele[8][33] != ele[27][33];
    ele[8][33] != ele[28][33];
    ele[8][33] != ele[29][33];
    ele[8][33] != ele[30][33];
    ele[8][33] != ele[31][33];
    ele[8][33] != ele[32][33];
    ele[8][33] != ele[33][33];
    ele[8][33] != ele[34][33];
    ele[8][33] != ele[35][33];
    ele[8][33] != ele[8][34];
    ele[8][33] != ele[8][35];
    ele[8][33] != ele[9][30];
    ele[8][33] != ele[9][31];
    ele[8][33] != ele[9][32];
    ele[8][33] != ele[9][33];
    ele[8][33] != ele[9][34];
    ele[8][33] != ele[9][35];
    ele[8][34] != ele[10][30];
    ele[8][34] != ele[10][31];
    ele[8][34] != ele[10][32];
    ele[8][34] != ele[10][33];
    ele[8][34] != ele[10][34];
    ele[8][34] != ele[10][35];
    ele[8][34] != ele[11][30];
    ele[8][34] != ele[11][31];
    ele[8][34] != ele[11][32];
    ele[8][34] != ele[11][33];
    ele[8][34] != ele[11][34];
    ele[8][34] != ele[11][35];
    ele[8][34] != ele[12][34];
    ele[8][34] != ele[13][34];
    ele[8][34] != ele[14][34];
    ele[8][34] != ele[15][34];
    ele[8][34] != ele[16][34];
    ele[8][34] != ele[17][34];
    ele[8][34] != ele[18][34];
    ele[8][34] != ele[19][34];
    ele[8][34] != ele[20][34];
    ele[8][34] != ele[21][34];
    ele[8][34] != ele[22][34];
    ele[8][34] != ele[23][34];
    ele[8][34] != ele[24][34];
    ele[8][34] != ele[25][34];
    ele[8][34] != ele[26][34];
    ele[8][34] != ele[27][34];
    ele[8][34] != ele[28][34];
    ele[8][34] != ele[29][34];
    ele[8][34] != ele[30][34];
    ele[8][34] != ele[31][34];
    ele[8][34] != ele[32][34];
    ele[8][34] != ele[33][34];
    ele[8][34] != ele[34][34];
    ele[8][34] != ele[35][34];
    ele[8][34] != ele[8][35];
    ele[8][34] != ele[9][30];
    ele[8][34] != ele[9][31];
    ele[8][34] != ele[9][32];
    ele[8][34] != ele[9][33];
    ele[8][34] != ele[9][34];
    ele[8][34] != ele[9][35];
    ele[8][35] != ele[10][30];
    ele[8][35] != ele[10][31];
    ele[8][35] != ele[10][32];
    ele[8][35] != ele[10][33];
    ele[8][35] != ele[10][34];
    ele[8][35] != ele[10][35];
    ele[8][35] != ele[11][30];
    ele[8][35] != ele[11][31];
    ele[8][35] != ele[11][32];
    ele[8][35] != ele[11][33];
    ele[8][35] != ele[11][34];
    ele[8][35] != ele[11][35];
    ele[8][35] != ele[12][35];
    ele[8][35] != ele[13][35];
    ele[8][35] != ele[14][35];
    ele[8][35] != ele[15][35];
    ele[8][35] != ele[16][35];
    ele[8][35] != ele[17][35];
    ele[8][35] != ele[18][35];
    ele[8][35] != ele[19][35];
    ele[8][35] != ele[20][35];
    ele[8][35] != ele[21][35];
    ele[8][35] != ele[22][35];
    ele[8][35] != ele[23][35];
    ele[8][35] != ele[24][35];
    ele[8][35] != ele[25][35];
    ele[8][35] != ele[26][35];
    ele[8][35] != ele[27][35];
    ele[8][35] != ele[28][35];
    ele[8][35] != ele[29][35];
    ele[8][35] != ele[30][35];
    ele[8][35] != ele[31][35];
    ele[8][35] != ele[32][35];
    ele[8][35] != ele[33][35];
    ele[8][35] != ele[34][35];
    ele[8][35] != ele[35][35];
    ele[8][35] != ele[9][30];
    ele[8][35] != ele[9][31];
    ele[8][35] != ele[9][32];
    ele[8][35] != ele[9][33];
    ele[8][35] != ele[9][34];
    ele[8][35] != ele[9][35];
    ele[8][4] != ele[10][0];
    ele[8][4] != ele[10][1];
    ele[8][4] != ele[10][2];
    ele[8][4] != ele[10][3];
    ele[8][4] != ele[10][4];
    ele[8][4] != ele[10][5];
    ele[8][4] != ele[11][0];
    ele[8][4] != ele[11][1];
    ele[8][4] != ele[11][2];
    ele[8][4] != ele[11][3];
    ele[8][4] != ele[11][4];
    ele[8][4] != ele[11][5];
    ele[8][4] != ele[12][4];
    ele[8][4] != ele[13][4];
    ele[8][4] != ele[14][4];
    ele[8][4] != ele[15][4];
    ele[8][4] != ele[16][4];
    ele[8][4] != ele[17][4];
    ele[8][4] != ele[18][4];
    ele[8][4] != ele[19][4];
    ele[8][4] != ele[20][4];
    ele[8][4] != ele[21][4];
    ele[8][4] != ele[22][4];
    ele[8][4] != ele[23][4];
    ele[8][4] != ele[24][4];
    ele[8][4] != ele[25][4];
    ele[8][4] != ele[26][4];
    ele[8][4] != ele[27][4];
    ele[8][4] != ele[28][4];
    ele[8][4] != ele[29][4];
    ele[8][4] != ele[30][4];
    ele[8][4] != ele[31][4];
    ele[8][4] != ele[32][4];
    ele[8][4] != ele[33][4];
    ele[8][4] != ele[34][4];
    ele[8][4] != ele[35][4];
    ele[8][4] != ele[8][10];
    ele[8][4] != ele[8][11];
    ele[8][4] != ele[8][12];
    ele[8][4] != ele[8][13];
    ele[8][4] != ele[8][14];
    ele[8][4] != ele[8][15];
    ele[8][4] != ele[8][16];
    ele[8][4] != ele[8][17];
    ele[8][4] != ele[8][18];
    ele[8][4] != ele[8][19];
    ele[8][4] != ele[8][20];
    ele[8][4] != ele[8][21];
    ele[8][4] != ele[8][22];
    ele[8][4] != ele[8][23];
    ele[8][4] != ele[8][24];
    ele[8][4] != ele[8][25];
    ele[8][4] != ele[8][26];
    ele[8][4] != ele[8][27];
    ele[8][4] != ele[8][28];
    ele[8][4] != ele[8][29];
    ele[8][4] != ele[8][30];
    ele[8][4] != ele[8][31];
    ele[8][4] != ele[8][32];
    ele[8][4] != ele[8][33];
    ele[8][4] != ele[8][34];
    ele[8][4] != ele[8][35];
    ele[8][4] != ele[8][5];
    ele[8][4] != ele[8][6];
    ele[8][4] != ele[8][7];
    ele[8][4] != ele[8][8];
    ele[8][4] != ele[8][9];
    ele[8][4] != ele[9][0];
    ele[8][4] != ele[9][1];
    ele[8][4] != ele[9][2];
    ele[8][4] != ele[9][3];
    ele[8][4] != ele[9][4];
    ele[8][4] != ele[9][5];
    ele[8][5] != ele[10][0];
    ele[8][5] != ele[10][1];
    ele[8][5] != ele[10][2];
    ele[8][5] != ele[10][3];
    ele[8][5] != ele[10][4];
    ele[8][5] != ele[10][5];
    ele[8][5] != ele[11][0];
    ele[8][5] != ele[11][1];
    ele[8][5] != ele[11][2];
    ele[8][5] != ele[11][3];
    ele[8][5] != ele[11][4];
    ele[8][5] != ele[11][5];
    ele[8][5] != ele[12][5];
    ele[8][5] != ele[13][5];
    ele[8][5] != ele[14][5];
    ele[8][5] != ele[15][5];
    ele[8][5] != ele[16][5];
    ele[8][5] != ele[17][5];
    ele[8][5] != ele[18][5];
    ele[8][5] != ele[19][5];
    ele[8][5] != ele[20][5];
    ele[8][5] != ele[21][5];
    ele[8][5] != ele[22][5];
    ele[8][5] != ele[23][5];
    ele[8][5] != ele[24][5];
    ele[8][5] != ele[25][5];
    ele[8][5] != ele[26][5];
    ele[8][5] != ele[27][5];
    ele[8][5] != ele[28][5];
    ele[8][5] != ele[29][5];
    ele[8][5] != ele[30][5];
    ele[8][5] != ele[31][5];
    ele[8][5] != ele[32][5];
    ele[8][5] != ele[33][5];
    ele[8][5] != ele[34][5];
    ele[8][5] != ele[35][5];
    ele[8][5] != ele[8][10];
    ele[8][5] != ele[8][11];
    ele[8][5] != ele[8][12];
    ele[8][5] != ele[8][13];
    ele[8][5] != ele[8][14];
    ele[8][5] != ele[8][15];
    ele[8][5] != ele[8][16];
    ele[8][5] != ele[8][17];
    ele[8][5] != ele[8][18];
    ele[8][5] != ele[8][19];
    ele[8][5] != ele[8][20];
    ele[8][5] != ele[8][21];
    ele[8][5] != ele[8][22];
    ele[8][5] != ele[8][23];
    ele[8][5] != ele[8][24];
    ele[8][5] != ele[8][25];
    ele[8][5] != ele[8][26];
    ele[8][5] != ele[8][27];
    ele[8][5] != ele[8][28];
    ele[8][5] != ele[8][29];
    ele[8][5] != ele[8][30];
    ele[8][5] != ele[8][31];
    ele[8][5] != ele[8][32];
    ele[8][5] != ele[8][33];
    ele[8][5] != ele[8][34];
    ele[8][5] != ele[8][35];
    ele[8][5] != ele[8][6];
    ele[8][5] != ele[8][7];
    ele[8][5] != ele[8][8];
    ele[8][5] != ele[8][9];
    ele[8][5] != ele[9][0];
    ele[8][5] != ele[9][1];
    ele[8][5] != ele[9][2];
    ele[8][5] != ele[9][3];
    ele[8][5] != ele[9][4];
    ele[8][5] != ele[9][5];
    ele[8][6] != ele[10][10];
    ele[8][6] != ele[10][11];
    ele[8][6] != ele[10][6];
    ele[8][6] != ele[10][7];
    ele[8][6] != ele[10][8];
    ele[8][6] != ele[10][9];
    ele[8][6] != ele[11][10];
    ele[8][6] != ele[11][11];
    ele[8][6] != ele[11][6];
    ele[8][6] != ele[11][7];
    ele[8][6] != ele[11][8];
    ele[8][6] != ele[11][9];
    ele[8][6] != ele[12][6];
    ele[8][6] != ele[13][6];
    ele[8][6] != ele[14][6];
    ele[8][6] != ele[15][6];
    ele[8][6] != ele[16][6];
    ele[8][6] != ele[17][6];
    ele[8][6] != ele[18][6];
    ele[8][6] != ele[19][6];
    ele[8][6] != ele[20][6];
    ele[8][6] != ele[21][6];
    ele[8][6] != ele[22][6];
    ele[8][6] != ele[23][6];
    ele[8][6] != ele[24][6];
    ele[8][6] != ele[25][6];
    ele[8][6] != ele[26][6];
    ele[8][6] != ele[27][6];
    ele[8][6] != ele[28][6];
    ele[8][6] != ele[29][6];
    ele[8][6] != ele[30][6];
    ele[8][6] != ele[31][6];
    ele[8][6] != ele[32][6];
    ele[8][6] != ele[33][6];
    ele[8][6] != ele[34][6];
    ele[8][6] != ele[35][6];
    ele[8][6] != ele[8][10];
    ele[8][6] != ele[8][11];
    ele[8][6] != ele[8][12];
    ele[8][6] != ele[8][13];
    ele[8][6] != ele[8][14];
    ele[8][6] != ele[8][15];
    ele[8][6] != ele[8][16];
    ele[8][6] != ele[8][17];
    ele[8][6] != ele[8][18];
    ele[8][6] != ele[8][19];
    ele[8][6] != ele[8][20];
    ele[8][6] != ele[8][21];
    ele[8][6] != ele[8][22];
    ele[8][6] != ele[8][23];
    ele[8][6] != ele[8][24];
    ele[8][6] != ele[8][25];
    ele[8][6] != ele[8][26];
    ele[8][6] != ele[8][27];
    ele[8][6] != ele[8][28];
    ele[8][6] != ele[8][29];
    ele[8][6] != ele[8][30];
    ele[8][6] != ele[8][31];
    ele[8][6] != ele[8][32];
    ele[8][6] != ele[8][33];
    ele[8][6] != ele[8][34];
    ele[8][6] != ele[8][35];
    ele[8][6] != ele[8][7];
    ele[8][6] != ele[8][8];
    ele[8][6] != ele[8][9];
    ele[8][6] != ele[9][10];
    ele[8][6] != ele[9][11];
    ele[8][6] != ele[9][6];
    ele[8][6] != ele[9][7];
    ele[8][6] != ele[9][8];
    ele[8][6] != ele[9][9];
    ele[8][7] != ele[10][10];
    ele[8][7] != ele[10][11];
    ele[8][7] != ele[10][6];
    ele[8][7] != ele[10][7];
    ele[8][7] != ele[10][8];
    ele[8][7] != ele[10][9];
    ele[8][7] != ele[11][10];
    ele[8][7] != ele[11][11];
    ele[8][7] != ele[11][6];
    ele[8][7] != ele[11][7];
    ele[8][7] != ele[11][8];
    ele[8][7] != ele[11][9];
    ele[8][7] != ele[12][7];
    ele[8][7] != ele[13][7];
    ele[8][7] != ele[14][7];
    ele[8][7] != ele[15][7];
    ele[8][7] != ele[16][7];
    ele[8][7] != ele[17][7];
    ele[8][7] != ele[18][7];
    ele[8][7] != ele[19][7];
    ele[8][7] != ele[20][7];
    ele[8][7] != ele[21][7];
    ele[8][7] != ele[22][7];
    ele[8][7] != ele[23][7];
    ele[8][7] != ele[24][7];
    ele[8][7] != ele[25][7];
    ele[8][7] != ele[26][7];
    ele[8][7] != ele[27][7];
    ele[8][7] != ele[28][7];
    ele[8][7] != ele[29][7];
    ele[8][7] != ele[30][7];
    ele[8][7] != ele[31][7];
    ele[8][7] != ele[32][7];
    ele[8][7] != ele[33][7];
    ele[8][7] != ele[34][7];
    ele[8][7] != ele[35][7];
    ele[8][7] != ele[8][10];
    ele[8][7] != ele[8][11];
    ele[8][7] != ele[8][12];
    ele[8][7] != ele[8][13];
    ele[8][7] != ele[8][14];
    ele[8][7] != ele[8][15];
    ele[8][7] != ele[8][16];
    ele[8][7] != ele[8][17];
    ele[8][7] != ele[8][18];
    ele[8][7] != ele[8][19];
    ele[8][7] != ele[8][20];
    ele[8][7] != ele[8][21];
    ele[8][7] != ele[8][22];
    ele[8][7] != ele[8][23];
    ele[8][7] != ele[8][24];
    ele[8][7] != ele[8][25];
    ele[8][7] != ele[8][26];
    ele[8][7] != ele[8][27];
    ele[8][7] != ele[8][28];
    ele[8][7] != ele[8][29];
    ele[8][7] != ele[8][30];
    ele[8][7] != ele[8][31];
    ele[8][7] != ele[8][32];
    ele[8][7] != ele[8][33];
    ele[8][7] != ele[8][34];
    ele[8][7] != ele[8][35];
    ele[8][7] != ele[8][8];
    ele[8][7] != ele[8][9];
    ele[8][7] != ele[9][10];
    ele[8][7] != ele[9][11];
    ele[8][7] != ele[9][6];
    ele[8][7] != ele[9][7];
    ele[8][7] != ele[9][8];
    ele[8][7] != ele[9][9];
    ele[8][8] != ele[10][10];
    ele[8][8] != ele[10][11];
    ele[8][8] != ele[10][6];
    ele[8][8] != ele[10][7];
    ele[8][8] != ele[10][8];
    ele[8][8] != ele[10][9];
    ele[8][8] != ele[11][10];
    ele[8][8] != ele[11][11];
    ele[8][8] != ele[11][6];
    ele[8][8] != ele[11][7];
    ele[8][8] != ele[11][8];
    ele[8][8] != ele[11][9];
    ele[8][8] != ele[12][8];
    ele[8][8] != ele[13][8];
    ele[8][8] != ele[14][8];
    ele[8][8] != ele[15][8];
    ele[8][8] != ele[16][8];
    ele[8][8] != ele[17][8];
    ele[8][8] != ele[18][8];
    ele[8][8] != ele[19][8];
    ele[8][8] != ele[20][8];
    ele[8][8] != ele[21][8];
    ele[8][8] != ele[22][8];
    ele[8][8] != ele[23][8];
    ele[8][8] != ele[24][8];
    ele[8][8] != ele[25][8];
    ele[8][8] != ele[26][8];
    ele[8][8] != ele[27][8];
    ele[8][8] != ele[28][8];
    ele[8][8] != ele[29][8];
    ele[8][8] != ele[30][8];
    ele[8][8] != ele[31][8];
    ele[8][8] != ele[32][8];
    ele[8][8] != ele[33][8];
    ele[8][8] != ele[34][8];
    ele[8][8] != ele[35][8];
    ele[8][8] != ele[8][10];
    ele[8][8] != ele[8][11];
    ele[8][8] != ele[8][12];
    ele[8][8] != ele[8][13];
    ele[8][8] != ele[8][14];
    ele[8][8] != ele[8][15];
    ele[8][8] != ele[8][16];
    ele[8][8] != ele[8][17];
    ele[8][8] != ele[8][18];
    ele[8][8] != ele[8][19];
    ele[8][8] != ele[8][20];
    ele[8][8] != ele[8][21];
    ele[8][8] != ele[8][22];
    ele[8][8] != ele[8][23];
    ele[8][8] != ele[8][24];
    ele[8][8] != ele[8][25];
    ele[8][8] != ele[8][26];
    ele[8][8] != ele[8][27];
    ele[8][8] != ele[8][28];
    ele[8][8] != ele[8][29];
    ele[8][8] != ele[8][30];
    ele[8][8] != ele[8][31];
    ele[8][8] != ele[8][32];
    ele[8][8] != ele[8][33];
    ele[8][8] != ele[8][34];
    ele[8][8] != ele[8][35];
    ele[8][8] != ele[8][9];
    ele[8][8] != ele[9][10];
    ele[8][8] != ele[9][11];
    ele[8][8] != ele[9][6];
    ele[8][8] != ele[9][7];
    ele[8][8] != ele[9][8];
    ele[8][8] != ele[9][9];
    ele[8][9] != ele[10][10];
    ele[8][9] != ele[10][11];
    ele[8][9] != ele[10][6];
    ele[8][9] != ele[10][7];
    ele[8][9] != ele[10][8];
    ele[8][9] != ele[10][9];
    ele[8][9] != ele[11][10];
    ele[8][9] != ele[11][11];
    ele[8][9] != ele[11][6];
    ele[8][9] != ele[11][7];
    ele[8][9] != ele[11][8];
    ele[8][9] != ele[11][9];
    ele[8][9] != ele[12][9];
    ele[8][9] != ele[13][9];
    ele[8][9] != ele[14][9];
    ele[8][9] != ele[15][9];
    ele[8][9] != ele[16][9];
    ele[8][9] != ele[17][9];
    ele[8][9] != ele[18][9];
    ele[8][9] != ele[19][9];
    ele[8][9] != ele[20][9];
    ele[8][9] != ele[21][9];
    ele[8][9] != ele[22][9];
    ele[8][9] != ele[23][9];
    ele[8][9] != ele[24][9];
    ele[8][9] != ele[25][9];
    ele[8][9] != ele[26][9];
    ele[8][9] != ele[27][9];
    ele[8][9] != ele[28][9];
    ele[8][9] != ele[29][9];
    ele[8][9] != ele[30][9];
    ele[8][9] != ele[31][9];
    ele[8][9] != ele[32][9];
    ele[8][9] != ele[33][9];
    ele[8][9] != ele[34][9];
    ele[8][9] != ele[35][9];
    ele[8][9] != ele[8][10];
    ele[8][9] != ele[8][11];
    ele[8][9] != ele[8][12];
    ele[8][9] != ele[8][13];
    ele[8][9] != ele[8][14];
    ele[8][9] != ele[8][15];
    ele[8][9] != ele[8][16];
    ele[8][9] != ele[8][17];
    ele[8][9] != ele[8][18];
    ele[8][9] != ele[8][19];
    ele[8][9] != ele[8][20];
    ele[8][9] != ele[8][21];
    ele[8][9] != ele[8][22];
    ele[8][9] != ele[8][23];
    ele[8][9] != ele[8][24];
    ele[8][9] != ele[8][25];
    ele[8][9] != ele[8][26];
    ele[8][9] != ele[8][27];
    ele[8][9] != ele[8][28];
    ele[8][9] != ele[8][29];
    ele[8][9] != ele[8][30];
    ele[8][9] != ele[8][31];
    ele[8][9] != ele[8][32];
    ele[8][9] != ele[8][33];
    ele[8][9] != ele[8][34];
    ele[8][9] != ele[8][35];
    ele[8][9] != ele[9][10];
    ele[8][9] != ele[9][11];
    ele[8][9] != ele[9][6];
    ele[8][9] != ele[9][7];
    ele[8][9] != ele[9][8];
    ele[8][9] != ele[9][9];
    ele[9][0] != ele[10][0];
    ele[9][0] != ele[10][1];
    ele[9][0] != ele[10][2];
    ele[9][0] != ele[10][3];
    ele[9][0] != ele[10][4];
    ele[9][0] != ele[10][5];
    ele[9][0] != ele[11][0];
    ele[9][0] != ele[11][1];
    ele[9][0] != ele[11][2];
    ele[9][0] != ele[11][3];
    ele[9][0] != ele[11][4];
    ele[9][0] != ele[11][5];
    ele[9][0] != ele[12][0];
    ele[9][0] != ele[13][0];
    ele[9][0] != ele[14][0];
    ele[9][0] != ele[15][0];
    ele[9][0] != ele[16][0];
    ele[9][0] != ele[17][0];
    ele[9][0] != ele[18][0];
    ele[9][0] != ele[19][0];
    ele[9][0] != ele[20][0];
    ele[9][0] != ele[21][0];
    ele[9][0] != ele[22][0];
    ele[9][0] != ele[23][0];
    ele[9][0] != ele[24][0];
    ele[9][0] != ele[25][0];
    ele[9][0] != ele[26][0];
    ele[9][0] != ele[27][0];
    ele[9][0] != ele[28][0];
    ele[9][0] != ele[29][0];
    ele[9][0] != ele[30][0];
    ele[9][0] != ele[31][0];
    ele[9][0] != ele[32][0];
    ele[9][0] != ele[33][0];
    ele[9][0] != ele[34][0];
    ele[9][0] != ele[35][0];
    ele[9][0] != ele[9][1];
    ele[9][0] != ele[9][10];
    ele[9][0] != ele[9][11];
    ele[9][0] != ele[9][12];
    ele[9][0] != ele[9][13];
    ele[9][0] != ele[9][14];
    ele[9][0] != ele[9][15];
    ele[9][0] != ele[9][16];
    ele[9][0] != ele[9][17];
    ele[9][0] != ele[9][18];
    ele[9][0] != ele[9][19];
    ele[9][0] != ele[9][2];
    ele[9][0] != ele[9][20];
    ele[9][0] != ele[9][21];
    ele[9][0] != ele[9][22];
    ele[9][0] != ele[9][23];
    ele[9][0] != ele[9][24];
    ele[9][0] != ele[9][25];
    ele[9][0] != ele[9][26];
    ele[9][0] != ele[9][27];
    ele[9][0] != ele[9][28];
    ele[9][0] != ele[9][29];
    ele[9][0] != ele[9][3];
    ele[9][0] != ele[9][30];
    ele[9][0] != ele[9][31];
    ele[9][0] != ele[9][32];
    ele[9][0] != ele[9][33];
    ele[9][0] != ele[9][34];
    ele[9][0] != ele[9][35];
    ele[9][0] != ele[9][4];
    ele[9][0] != ele[9][5];
    ele[9][0] != ele[9][6];
    ele[9][0] != ele[9][7];
    ele[9][0] != ele[9][8];
    ele[9][0] != ele[9][9];
    ele[9][1] != ele[10][0];
    ele[9][1] != ele[10][1];
    ele[9][1] != ele[10][2];
    ele[9][1] != ele[10][3];
    ele[9][1] != ele[10][4];
    ele[9][1] != ele[10][5];
    ele[9][1] != ele[11][0];
    ele[9][1] != ele[11][1];
    ele[9][1] != ele[11][2];
    ele[9][1] != ele[11][3];
    ele[9][1] != ele[11][4];
    ele[9][1] != ele[11][5];
    ele[9][1] != ele[12][1];
    ele[9][1] != ele[13][1];
    ele[9][1] != ele[14][1];
    ele[9][1] != ele[15][1];
    ele[9][1] != ele[16][1];
    ele[9][1] != ele[17][1];
    ele[9][1] != ele[18][1];
    ele[9][1] != ele[19][1];
    ele[9][1] != ele[20][1];
    ele[9][1] != ele[21][1];
    ele[9][1] != ele[22][1];
    ele[9][1] != ele[23][1];
    ele[9][1] != ele[24][1];
    ele[9][1] != ele[25][1];
    ele[9][1] != ele[26][1];
    ele[9][1] != ele[27][1];
    ele[9][1] != ele[28][1];
    ele[9][1] != ele[29][1];
    ele[9][1] != ele[30][1];
    ele[9][1] != ele[31][1];
    ele[9][1] != ele[32][1];
    ele[9][1] != ele[33][1];
    ele[9][1] != ele[34][1];
    ele[9][1] != ele[35][1];
    ele[9][1] != ele[9][10];
    ele[9][1] != ele[9][11];
    ele[9][1] != ele[9][12];
    ele[9][1] != ele[9][13];
    ele[9][1] != ele[9][14];
    ele[9][1] != ele[9][15];
    ele[9][1] != ele[9][16];
    ele[9][1] != ele[9][17];
    ele[9][1] != ele[9][18];
    ele[9][1] != ele[9][19];
    ele[9][1] != ele[9][2];
    ele[9][1] != ele[9][20];
    ele[9][1] != ele[9][21];
    ele[9][1] != ele[9][22];
    ele[9][1] != ele[9][23];
    ele[9][1] != ele[9][24];
    ele[9][1] != ele[9][25];
    ele[9][1] != ele[9][26];
    ele[9][1] != ele[9][27];
    ele[9][1] != ele[9][28];
    ele[9][1] != ele[9][29];
    ele[9][1] != ele[9][3];
    ele[9][1] != ele[9][30];
    ele[9][1] != ele[9][31];
    ele[9][1] != ele[9][32];
    ele[9][1] != ele[9][33];
    ele[9][1] != ele[9][34];
    ele[9][1] != ele[9][35];
    ele[9][1] != ele[9][4];
    ele[9][1] != ele[9][5];
    ele[9][1] != ele[9][6];
    ele[9][1] != ele[9][7];
    ele[9][1] != ele[9][8];
    ele[9][1] != ele[9][9];
    ele[9][10] != ele[10][10];
    ele[9][10] != ele[10][11];
    ele[9][10] != ele[10][6];
    ele[9][10] != ele[10][7];
    ele[9][10] != ele[10][8];
    ele[9][10] != ele[10][9];
    ele[9][10] != ele[11][10];
    ele[9][10] != ele[11][11];
    ele[9][10] != ele[11][6];
    ele[9][10] != ele[11][7];
    ele[9][10] != ele[11][8];
    ele[9][10] != ele[11][9];
    ele[9][10] != ele[12][10];
    ele[9][10] != ele[13][10];
    ele[9][10] != ele[14][10];
    ele[9][10] != ele[15][10];
    ele[9][10] != ele[16][10];
    ele[9][10] != ele[17][10];
    ele[9][10] != ele[18][10];
    ele[9][10] != ele[19][10];
    ele[9][10] != ele[20][10];
    ele[9][10] != ele[21][10];
    ele[9][10] != ele[22][10];
    ele[9][10] != ele[23][10];
    ele[9][10] != ele[24][10];
    ele[9][10] != ele[25][10];
    ele[9][10] != ele[26][10];
    ele[9][10] != ele[27][10];
    ele[9][10] != ele[28][10];
    ele[9][10] != ele[29][10];
    ele[9][10] != ele[30][10];
    ele[9][10] != ele[31][10];
    ele[9][10] != ele[32][10];
    ele[9][10] != ele[33][10];
    ele[9][10] != ele[34][10];
    ele[9][10] != ele[35][10];
    ele[9][10] != ele[9][11];
    ele[9][10] != ele[9][12];
    ele[9][10] != ele[9][13];
    ele[9][10] != ele[9][14];
    ele[9][10] != ele[9][15];
    ele[9][10] != ele[9][16];
    ele[9][10] != ele[9][17];
    ele[9][10] != ele[9][18];
    ele[9][10] != ele[9][19];
    ele[9][10] != ele[9][20];
    ele[9][10] != ele[9][21];
    ele[9][10] != ele[9][22];
    ele[9][10] != ele[9][23];
    ele[9][10] != ele[9][24];
    ele[9][10] != ele[9][25];
    ele[9][10] != ele[9][26];
    ele[9][10] != ele[9][27];
    ele[9][10] != ele[9][28];
    ele[9][10] != ele[9][29];
    ele[9][10] != ele[9][30];
    ele[9][10] != ele[9][31];
    ele[9][10] != ele[9][32];
    ele[9][10] != ele[9][33];
    ele[9][10] != ele[9][34];
    ele[9][10] != ele[9][35];
    ele[9][11] != ele[10][10];
    ele[9][11] != ele[10][11];
    ele[9][11] != ele[10][6];
    ele[9][11] != ele[10][7];
    ele[9][11] != ele[10][8];
    ele[9][11] != ele[10][9];
    ele[9][11] != ele[11][10];
    ele[9][11] != ele[11][11];
    ele[9][11] != ele[11][6];
    ele[9][11] != ele[11][7];
    ele[9][11] != ele[11][8];
    ele[9][11] != ele[11][9];
    ele[9][11] != ele[12][11];
    ele[9][11] != ele[13][11];
    ele[9][11] != ele[14][11];
    ele[9][11] != ele[15][11];
    ele[9][11] != ele[16][11];
    ele[9][11] != ele[17][11];
    ele[9][11] != ele[18][11];
    ele[9][11] != ele[19][11];
    ele[9][11] != ele[20][11];
    ele[9][11] != ele[21][11];
    ele[9][11] != ele[22][11];
    ele[9][11] != ele[23][11];
    ele[9][11] != ele[24][11];
    ele[9][11] != ele[25][11];
    ele[9][11] != ele[26][11];
    ele[9][11] != ele[27][11];
    ele[9][11] != ele[28][11];
    ele[9][11] != ele[29][11];
    ele[9][11] != ele[30][11];
    ele[9][11] != ele[31][11];
    ele[9][11] != ele[32][11];
    ele[9][11] != ele[33][11];
    ele[9][11] != ele[34][11];
    ele[9][11] != ele[35][11];
    ele[9][11] != ele[9][12];
    ele[9][11] != ele[9][13];
    ele[9][11] != ele[9][14];
    ele[9][11] != ele[9][15];
    ele[9][11] != ele[9][16];
    ele[9][11] != ele[9][17];
    ele[9][11] != ele[9][18];
    ele[9][11] != ele[9][19];
    ele[9][11] != ele[9][20];
    ele[9][11] != ele[9][21];
    ele[9][11] != ele[9][22];
    ele[9][11] != ele[9][23];
    ele[9][11] != ele[9][24];
    ele[9][11] != ele[9][25];
    ele[9][11] != ele[9][26];
    ele[9][11] != ele[9][27];
    ele[9][11] != ele[9][28];
    ele[9][11] != ele[9][29];
    ele[9][11] != ele[9][30];
    ele[9][11] != ele[9][31];
    ele[9][11] != ele[9][32];
    ele[9][11] != ele[9][33];
    ele[9][11] != ele[9][34];
    ele[9][11] != ele[9][35];
    ele[9][12] != ele[10][12];
    ele[9][12] != ele[10][13];
    ele[9][12] != ele[10][14];
    ele[9][12] != ele[10][15];
    ele[9][12] != ele[10][16];
    ele[9][12] != ele[10][17];
    ele[9][12] != ele[11][12];
    ele[9][12] != ele[11][13];
    ele[9][12] != ele[11][14];
    ele[9][12] != ele[11][15];
    ele[9][12] != ele[11][16];
    ele[9][12] != ele[11][17];
    ele[9][12] != ele[12][12];
    ele[9][12] != ele[13][12];
    ele[9][12] != ele[14][12];
    ele[9][12] != ele[15][12];
    ele[9][12] != ele[16][12];
    ele[9][12] != ele[17][12];
    ele[9][12] != ele[18][12];
    ele[9][12] != ele[19][12];
    ele[9][12] != ele[20][12];
    ele[9][12] != ele[21][12];
    ele[9][12] != ele[22][12];
    ele[9][12] != ele[23][12];
    ele[9][12] != ele[24][12];
    ele[9][12] != ele[25][12];
    ele[9][12] != ele[26][12];
    ele[9][12] != ele[27][12];
    ele[9][12] != ele[28][12];
    ele[9][12] != ele[29][12];
    ele[9][12] != ele[30][12];
    ele[9][12] != ele[31][12];
    ele[9][12] != ele[32][12];
    ele[9][12] != ele[33][12];
    ele[9][12] != ele[34][12];
    ele[9][12] != ele[35][12];
    ele[9][12] != ele[9][13];
    ele[9][12] != ele[9][14];
    ele[9][12] != ele[9][15];
    ele[9][12] != ele[9][16];
    ele[9][12] != ele[9][17];
    ele[9][12] != ele[9][18];
    ele[9][12] != ele[9][19];
    ele[9][12] != ele[9][20];
    ele[9][12] != ele[9][21];
    ele[9][12] != ele[9][22];
    ele[9][12] != ele[9][23];
    ele[9][12] != ele[9][24];
    ele[9][12] != ele[9][25];
    ele[9][12] != ele[9][26];
    ele[9][12] != ele[9][27];
    ele[9][12] != ele[9][28];
    ele[9][12] != ele[9][29];
    ele[9][12] != ele[9][30];
    ele[9][12] != ele[9][31];
    ele[9][12] != ele[9][32];
    ele[9][12] != ele[9][33];
    ele[9][12] != ele[9][34];
    ele[9][12] != ele[9][35];
    ele[9][13] != ele[10][12];
    ele[9][13] != ele[10][13];
    ele[9][13] != ele[10][14];
    ele[9][13] != ele[10][15];
    ele[9][13] != ele[10][16];
    ele[9][13] != ele[10][17];
    ele[9][13] != ele[11][12];
    ele[9][13] != ele[11][13];
    ele[9][13] != ele[11][14];
    ele[9][13] != ele[11][15];
    ele[9][13] != ele[11][16];
    ele[9][13] != ele[11][17];
    ele[9][13] != ele[12][13];
    ele[9][13] != ele[13][13];
    ele[9][13] != ele[14][13];
    ele[9][13] != ele[15][13];
    ele[9][13] != ele[16][13];
    ele[9][13] != ele[17][13];
    ele[9][13] != ele[18][13];
    ele[9][13] != ele[19][13];
    ele[9][13] != ele[20][13];
    ele[9][13] != ele[21][13];
    ele[9][13] != ele[22][13];
    ele[9][13] != ele[23][13];
    ele[9][13] != ele[24][13];
    ele[9][13] != ele[25][13];
    ele[9][13] != ele[26][13];
    ele[9][13] != ele[27][13];
    ele[9][13] != ele[28][13];
    ele[9][13] != ele[29][13];
    ele[9][13] != ele[30][13];
    ele[9][13] != ele[31][13];
    ele[9][13] != ele[32][13];
    ele[9][13] != ele[33][13];
    ele[9][13] != ele[34][13];
    ele[9][13] != ele[35][13];
    ele[9][13] != ele[9][14];
    ele[9][13] != ele[9][15];
    ele[9][13] != ele[9][16];
    ele[9][13] != ele[9][17];
    ele[9][13] != ele[9][18];
    ele[9][13] != ele[9][19];
    ele[9][13] != ele[9][20];
    ele[9][13] != ele[9][21];
    ele[9][13] != ele[9][22];
    ele[9][13] != ele[9][23];
    ele[9][13] != ele[9][24];
    ele[9][13] != ele[9][25];
    ele[9][13] != ele[9][26];
    ele[9][13] != ele[9][27];
    ele[9][13] != ele[9][28];
    ele[9][13] != ele[9][29];
    ele[9][13] != ele[9][30];
    ele[9][13] != ele[9][31];
    ele[9][13] != ele[9][32];
    ele[9][13] != ele[9][33];
    ele[9][13] != ele[9][34];
    ele[9][13] != ele[9][35];
    ele[9][14] != ele[10][12];
    ele[9][14] != ele[10][13];
    ele[9][14] != ele[10][14];
    ele[9][14] != ele[10][15];
    ele[9][14] != ele[10][16];
    ele[9][14] != ele[10][17];
    ele[9][14] != ele[11][12];
    ele[9][14] != ele[11][13];
    ele[9][14] != ele[11][14];
    ele[9][14] != ele[11][15];
    ele[9][14] != ele[11][16];
    ele[9][14] != ele[11][17];
    ele[9][14] != ele[12][14];
    ele[9][14] != ele[13][14];
    ele[9][14] != ele[14][14];
    ele[9][14] != ele[15][14];
    ele[9][14] != ele[16][14];
    ele[9][14] != ele[17][14];
    ele[9][14] != ele[18][14];
    ele[9][14] != ele[19][14];
    ele[9][14] != ele[20][14];
    ele[9][14] != ele[21][14];
    ele[9][14] != ele[22][14];
    ele[9][14] != ele[23][14];
    ele[9][14] != ele[24][14];
    ele[9][14] != ele[25][14];
    ele[9][14] != ele[26][14];
    ele[9][14] != ele[27][14];
    ele[9][14] != ele[28][14];
    ele[9][14] != ele[29][14];
    ele[9][14] != ele[30][14];
    ele[9][14] != ele[31][14];
    ele[9][14] != ele[32][14];
    ele[9][14] != ele[33][14];
    ele[9][14] != ele[34][14];
    ele[9][14] != ele[35][14];
    ele[9][14] != ele[9][15];
    ele[9][14] != ele[9][16];
    ele[9][14] != ele[9][17];
    ele[9][14] != ele[9][18];
    ele[9][14] != ele[9][19];
    ele[9][14] != ele[9][20];
    ele[9][14] != ele[9][21];
    ele[9][14] != ele[9][22];
    ele[9][14] != ele[9][23];
    ele[9][14] != ele[9][24];
    ele[9][14] != ele[9][25];
    ele[9][14] != ele[9][26];
    ele[9][14] != ele[9][27];
    ele[9][14] != ele[9][28];
    ele[9][14] != ele[9][29];
    ele[9][14] != ele[9][30];
    ele[9][14] != ele[9][31];
    ele[9][14] != ele[9][32];
    ele[9][14] != ele[9][33];
    ele[9][14] != ele[9][34];
    ele[9][14] != ele[9][35];
    ele[9][15] != ele[10][12];
    ele[9][15] != ele[10][13];
    ele[9][15] != ele[10][14];
    ele[9][15] != ele[10][15];
    ele[9][15] != ele[10][16];
    ele[9][15] != ele[10][17];
    ele[9][15] != ele[11][12];
    ele[9][15] != ele[11][13];
    ele[9][15] != ele[11][14];
    ele[9][15] != ele[11][15];
    ele[9][15] != ele[11][16];
    ele[9][15] != ele[11][17];
    ele[9][15] != ele[12][15];
    ele[9][15] != ele[13][15];
    ele[9][15] != ele[14][15];
    ele[9][15] != ele[15][15];
    ele[9][15] != ele[16][15];
    ele[9][15] != ele[17][15];
    ele[9][15] != ele[18][15];
    ele[9][15] != ele[19][15];
    ele[9][15] != ele[20][15];
    ele[9][15] != ele[21][15];
    ele[9][15] != ele[22][15];
    ele[9][15] != ele[23][15];
    ele[9][15] != ele[24][15];
    ele[9][15] != ele[25][15];
    ele[9][15] != ele[26][15];
    ele[9][15] != ele[27][15];
    ele[9][15] != ele[28][15];
    ele[9][15] != ele[29][15];
    ele[9][15] != ele[30][15];
    ele[9][15] != ele[31][15];
    ele[9][15] != ele[32][15];
    ele[9][15] != ele[33][15];
    ele[9][15] != ele[34][15];
    ele[9][15] != ele[35][15];
    ele[9][15] != ele[9][16];
    ele[9][15] != ele[9][17];
    ele[9][15] != ele[9][18];
    ele[9][15] != ele[9][19];
    ele[9][15] != ele[9][20];
    ele[9][15] != ele[9][21];
    ele[9][15] != ele[9][22];
    ele[9][15] != ele[9][23];
    ele[9][15] != ele[9][24];
    ele[9][15] != ele[9][25];
    ele[9][15] != ele[9][26];
    ele[9][15] != ele[9][27];
    ele[9][15] != ele[9][28];
    ele[9][15] != ele[9][29];
    ele[9][15] != ele[9][30];
    ele[9][15] != ele[9][31];
    ele[9][15] != ele[9][32];
    ele[9][15] != ele[9][33];
    ele[9][15] != ele[9][34];
    ele[9][15] != ele[9][35];
    ele[9][16] != ele[10][12];
    ele[9][16] != ele[10][13];
    ele[9][16] != ele[10][14];
    ele[9][16] != ele[10][15];
    ele[9][16] != ele[10][16];
    ele[9][16] != ele[10][17];
    ele[9][16] != ele[11][12];
    ele[9][16] != ele[11][13];
    ele[9][16] != ele[11][14];
    ele[9][16] != ele[11][15];
    ele[9][16] != ele[11][16];
    ele[9][16] != ele[11][17];
    ele[9][16] != ele[12][16];
    ele[9][16] != ele[13][16];
    ele[9][16] != ele[14][16];
    ele[9][16] != ele[15][16];
    ele[9][16] != ele[16][16];
    ele[9][16] != ele[17][16];
    ele[9][16] != ele[18][16];
    ele[9][16] != ele[19][16];
    ele[9][16] != ele[20][16];
    ele[9][16] != ele[21][16];
    ele[9][16] != ele[22][16];
    ele[9][16] != ele[23][16];
    ele[9][16] != ele[24][16];
    ele[9][16] != ele[25][16];
    ele[9][16] != ele[26][16];
    ele[9][16] != ele[27][16];
    ele[9][16] != ele[28][16];
    ele[9][16] != ele[29][16];
    ele[9][16] != ele[30][16];
    ele[9][16] != ele[31][16];
    ele[9][16] != ele[32][16];
    ele[9][16] != ele[33][16];
    ele[9][16] != ele[34][16];
    ele[9][16] != ele[35][16];
    ele[9][16] != ele[9][17];
    ele[9][16] != ele[9][18];
    ele[9][16] != ele[9][19];
    ele[9][16] != ele[9][20];
    ele[9][16] != ele[9][21];
    ele[9][16] != ele[9][22];
    ele[9][16] != ele[9][23];
    ele[9][16] != ele[9][24];
    ele[9][16] != ele[9][25];
    ele[9][16] != ele[9][26];
    ele[9][16] != ele[9][27];
    ele[9][16] != ele[9][28];
    ele[9][16] != ele[9][29];
    ele[9][16] != ele[9][30];
    ele[9][16] != ele[9][31];
    ele[9][16] != ele[9][32];
    ele[9][16] != ele[9][33];
    ele[9][16] != ele[9][34];
    ele[9][16] != ele[9][35];
    ele[9][17] != ele[10][12];
    ele[9][17] != ele[10][13];
    ele[9][17] != ele[10][14];
    ele[9][17] != ele[10][15];
    ele[9][17] != ele[10][16];
    ele[9][17] != ele[10][17];
    ele[9][17] != ele[11][12];
    ele[9][17] != ele[11][13];
    ele[9][17] != ele[11][14];
    ele[9][17] != ele[11][15];
    ele[9][17] != ele[11][16];
    ele[9][17] != ele[11][17];
    ele[9][17] != ele[12][17];
    ele[9][17] != ele[13][17];
    ele[9][17] != ele[14][17];
    ele[9][17] != ele[15][17];
    ele[9][17] != ele[16][17];
    ele[9][17] != ele[17][17];
    ele[9][17] != ele[18][17];
    ele[9][17] != ele[19][17];
    ele[9][17] != ele[20][17];
    ele[9][17] != ele[21][17];
    ele[9][17] != ele[22][17];
    ele[9][17] != ele[23][17];
    ele[9][17] != ele[24][17];
    ele[9][17] != ele[25][17];
    ele[9][17] != ele[26][17];
    ele[9][17] != ele[27][17];
    ele[9][17] != ele[28][17];
    ele[9][17] != ele[29][17];
    ele[9][17] != ele[30][17];
    ele[9][17] != ele[31][17];
    ele[9][17] != ele[32][17];
    ele[9][17] != ele[33][17];
    ele[9][17] != ele[34][17];
    ele[9][17] != ele[35][17];
    ele[9][17] != ele[9][18];
    ele[9][17] != ele[9][19];
    ele[9][17] != ele[9][20];
    ele[9][17] != ele[9][21];
    ele[9][17] != ele[9][22];
    ele[9][17] != ele[9][23];
    ele[9][17] != ele[9][24];
    ele[9][17] != ele[9][25];
    ele[9][17] != ele[9][26];
    ele[9][17] != ele[9][27];
    ele[9][17] != ele[9][28];
    ele[9][17] != ele[9][29];
    ele[9][17] != ele[9][30];
    ele[9][17] != ele[9][31];
    ele[9][17] != ele[9][32];
    ele[9][17] != ele[9][33];
    ele[9][17] != ele[9][34];
    ele[9][17] != ele[9][35];
    ele[9][18] != ele[10][18];
    ele[9][18] != ele[10][19];
    ele[9][18] != ele[10][20];
    ele[9][18] != ele[10][21];
    ele[9][18] != ele[10][22];
    ele[9][18] != ele[10][23];
    ele[9][18] != ele[11][18];
    ele[9][18] != ele[11][19];
    ele[9][18] != ele[11][20];
    ele[9][18] != ele[11][21];
    ele[9][18] != ele[11][22];
    ele[9][18] != ele[11][23];
    ele[9][18] != ele[12][18];
    ele[9][18] != ele[13][18];
    ele[9][18] != ele[14][18];
    ele[9][18] != ele[15][18];
    ele[9][18] != ele[16][18];
    ele[9][18] != ele[17][18];
    ele[9][18] != ele[18][18];
    ele[9][18] != ele[19][18];
    ele[9][18] != ele[20][18];
    ele[9][18] != ele[21][18];
    ele[9][18] != ele[22][18];
    ele[9][18] != ele[23][18];
    ele[9][18] != ele[24][18];
    ele[9][18] != ele[25][18];
    ele[9][18] != ele[26][18];
    ele[9][18] != ele[27][18];
    ele[9][18] != ele[28][18];
    ele[9][18] != ele[29][18];
    ele[9][18] != ele[30][18];
    ele[9][18] != ele[31][18];
    ele[9][18] != ele[32][18];
    ele[9][18] != ele[33][18];
    ele[9][18] != ele[34][18];
    ele[9][18] != ele[35][18];
    ele[9][18] != ele[9][19];
    ele[9][18] != ele[9][20];
    ele[9][18] != ele[9][21];
    ele[9][18] != ele[9][22];
    ele[9][18] != ele[9][23];
    ele[9][18] != ele[9][24];
    ele[9][18] != ele[9][25];
    ele[9][18] != ele[9][26];
    ele[9][18] != ele[9][27];
    ele[9][18] != ele[9][28];
    ele[9][18] != ele[9][29];
    ele[9][18] != ele[9][30];
    ele[9][18] != ele[9][31];
    ele[9][18] != ele[9][32];
    ele[9][18] != ele[9][33];
    ele[9][18] != ele[9][34];
    ele[9][18] != ele[9][35];
    ele[9][19] != ele[10][18];
    ele[9][19] != ele[10][19];
    ele[9][19] != ele[10][20];
    ele[9][19] != ele[10][21];
    ele[9][19] != ele[10][22];
    ele[9][19] != ele[10][23];
    ele[9][19] != ele[11][18];
    ele[9][19] != ele[11][19];
    ele[9][19] != ele[11][20];
    ele[9][19] != ele[11][21];
    ele[9][19] != ele[11][22];
    ele[9][19] != ele[11][23];
    ele[9][19] != ele[12][19];
    ele[9][19] != ele[13][19];
    ele[9][19] != ele[14][19];
    ele[9][19] != ele[15][19];
    ele[9][19] != ele[16][19];
    ele[9][19] != ele[17][19];
    ele[9][19] != ele[18][19];
    ele[9][19] != ele[19][19];
    ele[9][19] != ele[20][19];
    ele[9][19] != ele[21][19];
    ele[9][19] != ele[22][19];
    ele[9][19] != ele[23][19];
    ele[9][19] != ele[24][19];
    ele[9][19] != ele[25][19];
    ele[9][19] != ele[26][19];
    ele[9][19] != ele[27][19];
    ele[9][19] != ele[28][19];
    ele[9][19] != ele[29][19];
    ele[9][19] != ele[30][19];
    ele[9][19] != ele[31][19];
    ele[9][19] != ele[32][19];
    ele[9][19] != ele[33][19];
    ele[9][19] != ele[34][19];
    ele[9][19] != ele[35][19];
    ele[9][19] != ele[9][20];
    ele[9][19] != ele[9][21];
    ele[9][19] != ele[9][22];
    ele[9][19] != ele[9][23];
    ele[9][19] != ele[9][24];
    ele[9][19] != ele[9][25];
    ele[9][19] != ele[9][26];
    ele[9][19] != ele[9][27];
    ele[9][19] != ele[9][28];
    ele[9][19] != ele[9][29];
    ele[9][19] != ele[9][30];
    ele[9][19] != ele[9][31];
    ele[9][19] != ele[9][32];
    ele[9][19] != ele[9][33];
    ele[9][19] != ele[9][34];
    ele[9][19] != ele[9][35];
    ele[9][2] != ele[10][0];
    ele[9][2] != ele[10][1];
    ele[9][2] != ele[10][2];
    ele[9][2] != ele[10][3];
    ele[9][2] != ele[10][4];
    ele[9][2] != ele[10][5];
    ele[9][2] != ele[11][0];
    ele[9][2] != ele[11][1];
    ele[9][2] != ele[11][2];
    ele[9][2] != ele[11][3];
    ele[9][2] != ele[11][4];
    ele[9][2] != ele[11][5];
    ele[9][2] != ele[12][2];
    ele[9][2] != ele[13][2];
    ele[9][2] != ele[14][2];
    ele[9][2] != ele[15][2];
    ele[9][2] != ele[16][2];
    ele[9][2] != ele[17][2];
    ele[9][2] != ele[18][2];
    ele[9][2] != ele[19][2];
    ele[9][2] != ele[20][2];
    ele[9][2] != ele[21][2];
    ele[9][2] != ele[22][2];
    ele[9][2] != ele[23][2];
    ele[9][2] != ele[24][2];
    ele[9][2] != ele[25][2];
    ele[9][2] != ele[26][2];
    ele[9][2] != ele[27][2];
    ele[9][2] != ele[28][2];
    ele[9][2] != ele[29][2];
    ele[9][2] != ele[30][2];
    ele[9][2] != ele[31][2];
    ele[9][2] != ele[32][2];
    ele[9][2] != ele[33][2];
    ele[9][2] != ele[34][2];
    ele[9][2] != ele[35][2];
    ele[9][2] != ele[9][10];
    ele[9][2] != ele[9][11];
    ele[9][2] != ele[9][12];
    ele[9][2] != ele[9][13];
    ele[9][2] != ele[9][14];
    ele[9][2] != ele[9][15];
    ele[9][2] != ele[9][16];
    ele[9][2] != ele[9][17];
    ele[9][2] != ele[9][18];
    ele[9][2] != ele[9][19];
    ele[9][2] != ele[9][20];
    ele[9][2] != ele[9][21];
    ele[9][2] != ele[9][22];
    ele[9][2] != ele[9][23];
    ele[9][2] != ele[9][24];
    ele[9][2] != ele[9][25];
    ele[9][2] != ele[9][26];
    ele[9][2] != ele[9][27];
    ele[9][2] != ele[9][28];
    ele[9][2] != ele[9][29];
    ele[9][2] != ele[9][3];
    ele[9][2] != ele[9][30];
    ele[9][2] != ele[9][31];
    ele[9][2] != ele[9][32];
    ele[9][2] != ele[9][33];
    ele[9][2] != ele[9][34];
    ele[9][2] != ele[9][35];
    ele[9][2] != ele[9][4];
    ele[9][2] != ele[9][5];
    ele[9][2] != ele[9][6];
    ele[9][2] != ele[9][7];
    ele[9][2] != ele[9][8];
    ele[9][2] != ele[9][9];
    ele[9][20] != ele[10][18];
    ele[9][20] != ele[10][19];
    ele[9][20] != ele[10][20];
    ele[9][20] != ele[10][21];
    ele[9][20] != ele[10][22];
    ele[9][20] != ele[10][23];
    ele[9][20] != ele[11][18];
    ele[9][20] != ele[11][19];
    ele[9][20] != ele[11][20];
    ele[9][20] != ele[11][21];
    ele[9][20] != ele[11][22];
    ele[9][20] != ele[11][23];
    ele[9][20] != ele[12][20];
    ele[9][20] != ele[13][20];
    ele[9][20] != ele[14][20];
    ele[9][20] != ele[15][20];
    ele[9][20] != ele[16][20];
    ele[9][20] != ele[17][20];
    ele[9][20] != ele[18][20];
    ele[9][20] != ele[19][20];
    ele[9][20] != ele[20][20];
    ele[9][20] != ele[21][20];
    ele[9][20] != ele[22][20];
    ele[9][20] != ele[23][20];
    ele[9][20] != ele[24][20];
    ele[9][20] != ele[25][20];
    ele[9][20] != ele[26][20];
    ele[9][20] != ele[27][20];
    ele[9][20] != ele[28][20];
    ele[9][20] != ele[29][20];
    ele[9][20] != ele[30][20];
    ele[9][20] != ele[31][20];
    ele[9][20] != ele[32][20];
    ele[9][20] != ele[33][20];
    ele[9][20] != ele[34][20];
    ele[9][20] != ele[35][20];
    ele[9][20] != ele[9][21];
    ele[9][20] != ele[9][22];
    ele[9][20] != ele[9][23];
    ele[9][20] != ele[9][24];
    ele[9][20] != ele[9][25];
    ele[9][20] != ele[9][26];
    ele[9][20] != ele[9][27];
    ele[9][20] != ele[9][28];
    ele[9][20] != ele[9][29];
    ele[9][20] != ele[9][30];
    ele[9][20] != ele[9][31];
    ele[9][20] != ele[9][32];
    ele[9][20] != ele[9][33];
    ele[9][20] != ele[9][34];
    ele[9][20] != ele[9][35];
    ele[9][21] != ele[10][18];
    ele[9][21] != ele[10][19];
    ele[9][21] != ele[10][20];
    ele[9][21] != ele[10][21];
    ele[9][21] != ele[10][22];
    ele[9][21] != ele[10][23];
    ele[9][21] != ele[11][18];
    ele[9][21] != ele[11][19];
    ele[9][21] != ele[11][20];
    ele[9][21] != ele[11][21];
    ele[9][21] != ele[11][22];
    ele[9][21] != ele[11][23];
    ele[9][21] != ele[12][21];
    ele[9][21] != ele[13][21];
    ele[9][21] != ele[14][21];
    ele[9][21] != ele[15][21];
    ele[9][21] != ele[16][21];
    ele[9][21] != ele[17][21];
    ele[9][21] != ele[18][21];
    ele[9][21] != ele[19][21];
    ele[9][21] != ele[20][21];
    ele[9][21] != ele[21][21];
    ele[9][21] != ele[22][21];
    ele[9][21] != ele[23][21];
    ele[9][21] != ele[24][21];
    ele[9][21] != ele[25][21];
    ele[9][21] != ele[26][21];
    ele[9][21] != ele[27][21];
    ele[9][21] != ele[28][21];
    ele[9][21] != ele[29][21];
    ele[9][21] != ele[30][21];
    ele[9][21] != ele[31][21];
    ele[9][21] != ele[32][21];
    ele[9][21] != ele[33][21];
    ele[9][21] != ele[34][21];
    ele[9][21] != ele[35][21];
    ele[9][21] != ele[9][22];
    ele[9][21] != ele[9][23];
    ele[9][21] != ele[9][24];
    ele[9][21] != ele[9][25];
    ele[9][21] != ele[9][26];
    ele[9][21] != ele[9][27];
    ele[9][21] != ele[9][28];
    ele[9][21] != ele[9][29];
    ele[9][21] != ele[9][30];
    ele[9][21] != ele[9][31];
    ele[9][21] != ele[9][32];
    ele[9][21] != ele[9][33];
    ele[9][21] != ele[9][34];
    ele[9][21] != ele[9][35];
    ele[9][22] != ele[10][18];
    ele[9][22] != ele[10][19];
    ele[9][22] != ele[10][20];
    ele[9][22] != ele[10][21];
    ele[9][22] != ele[10][22];
    ele[9][22] != ele[10][23];
    ele[9][22] != ele[11][18];
    ele[9][22] != ele[11][19];
    ele[9][22] != ele[11][20];
    ele[9][22] != ele[11][21];
    ele[9][22] != ele[11][22];
    ele[9][22] != ele[11][23];
    ele[9][22] != ele[12][22];
    ele[9][22] != ele[13][22];
    ele[9][22] != ele[14][22];
    ele[9][22] != ele[15][22];
    ele[9][22] != ele[16][22];
    ele[9][22] != ele[17][22];
    ele[9][22] != ele[18][22];
    ele[9][22] != ele[19][22];
    ele[9][22] != ele[20][22];
    ele[9][22] != ele[21][22];
    ele[9][22] != ele[22][22];
    ele[9][22] != ele[23][22];
    ele[9][22] != ele[24][22];
    ele[9][22] != ele[25][22];
    ele[9][22] != ele[26][22];
    ele[9][22] != ele[27][22];
    ele[9][22] != ele[28][22];
    ele[9][22] != ele[29][22];
    ele[9][22] != ele[30][22];
    ele[9][22] != ele[31][22];
    ele[9][22] != ele[32][22];
    ele[9][22] != ele[33][22];
    ele[9][22] != ele[34][22];
    ele[9][22] != ele[35][22];
    ele[9][22] != ele[9][23];
    ele[9][22] != ele[9][24];
    ele[9][22] != ele[9][25];
    ele[9][22] != ele[9][26];
    ele[9][22] != ele[9][27];
    ele[9][22] != ele[9][28];
    ele[9][22] != ele[9][29];
    ele[9][22] != ele[9][30];
    ele[9][22] != ele[9][31];
    ele[9][22] != ele[9][32];
    ele[9][22] != ele[9][33];
    ele[9][22] != ele[9][34];
    ele[9][22] != ele[9][35];
    ele[9][23] != ele[10][18];
    ele[9][23] != ele[10][19];
    ele[9][23] != ele[10][20];
    ele[9][23] != ele[10][21];
    ele[9][23] != ele[10][22];
    ele[9][23] != ele[10][23];
    ele[9][23] != ele[11][18];
    ele[9][23] != ele[11][19];
    ele[9][23] != ele[11][20];
    ele[9][23] != ele[11][21];
    ele[9][23] != ele[11][22];
    ele[9][23] != ele[11][23];
    ele[9][23] != ele[12][23];
    ele[9][23] != ele[13][23];
    ele[9][23] != ele[14][23];
    ele[9][23] != ele[15][23];
    ele[9][23] != ele[16][23];
    ele[9][23] != ele[17][23];
    ele[9][23] != ele[18][23];
    ele[9][23] != ele[19][23];
    ele[9][23] != ele[20][23];
    ele[9][23] != ele[21][23];
    ele[9][23] != ele[22][23];
    ele[9][23] != ele[23][23];
    ele[9][23] != ele[24][23];
    ele[9][23] != ele[25][23];
    ele[9][23] != ele[26][23];
    ele[9][23] != ele[27][23];
    ele[9][23] != ele[28][23];
    ele[9][23] != ele[29][23];
    ele[9][23] != ele[30][23];
    ele[9][23] != ele[31][23];
    ele[9][23] != ele[32][23];
    ele[9][23] != ele[33][23];
    ele[9][23] != ele[34][23];
    ele[9][23] != ele[35][23];
    ele[9][23] != ele[9][24];
    ele[9][23] != ele[9][25];
    ele[9][23] != ele[9][26];
    ele[9][23] != ele[9][27];
    ele[9][23] != ele[9][28];
    ele[9][23] != ele[9][29];
    ele[9][23] != ele[9][30];
    ele[9][23] != ele[9][31];
    ele[9][23] != ele[9][32];
    ele[9][23] != ele[9][33];
    ele[9][23] != ele[9][34];
    ele[9][23] != ele[9][35];
    ele[9][24] != ele[10][24];
    ele[9][24] != ele[10][25];
    ele[9][24] != ele[10][26];
    ele[9][24] != ele[10][27];
    ele[9][24] != ele[10][28];
    ele[9][24] != ele[10][29];
    ele[9][24] != ele[11][24];
    ele[9][24] != ele[11][25];
    ele[9][24] != ele[11][26];
    ele[9][24] != ele[11][27];
    ele[9][24] != ele[11][28];
    ele[9][24] != ele[11][29];
    ele[9][24] != ele[12][24];
    ele[9][24] != ele[13][24];
    ele[9][24] != ele[14][24];
    ele[9][24] != ele[15][24];
    ele[9][24] != ele[16][24];
    ele[9][24] != ele[17][24];
    ele[9][24] != ele[18][24];
    ele[9][24] != ele[19][24];
    ele[9][24] != ele[20][24];
    ele[9][24] != ele[21][24];
    ele[9][24] != ele[22][24];
    ele[9][24] != ele[23][24];
    ele[9][24] != ele[24][24];
    ele[9][24] != ele[25][24];
    ele[9][24] != ele[26][24];
    ele[9][24] != ele[27][24];
    ele[9][24] != ele[28][24];
    ele[9][24] != ele[29][24];
    ele[9][24] != ele[30][24];
    ele[9][24] != ele[31][24];
    ele[9][24] != ele[32][24];
    ele[9][24] != ele[33][24];
    ele[9][24] != ele[34][24];
    ele[9][24] != ele[35][24];
    ele[9][24] != ele[9][25];
    ele[9][24] != ele[9][26];
    ele[9][24] != ele[9][27];
    ele[9][24] != ele[9][28];
    ele[9][24] != ele[9][29];
    ele[9][24] != ele[9][30];
    ele[9][24] != ele[9][31];
    ele[9][24] != ele[9][32];
    ele[9][24] != ele[9][33];
    ele[9][24] != ele[9][34];
    ele[9][24] != ele[9][35];
    ele[9][25] != ele[10][24];
    ele[9][25] != ele[10][25];
    ele[9][25] != ele[10][26];
    ele[9][25] != ele[10][27];
    ele[9][25] != ele[10][28];
    ele[9][25] != ele[10][29];
    ele[9][25] != ele[11][24];
    ele[9][25] != ele[11][25];
    ele[9][25] != ele[11][26];
    ele[9][25] != ele[11][27];
    ele[9][25] != ele[11][28];
    ele[9][25] != ele[11][29];
    ele[9][25] != ele[12][25];
    ele[9][25] != ele[13][25];
    ele[9][25] != ele[14][25];
    ele[9][25] != ele[15][25];
    ele[9][25] != ele[16][25];
    ele[9][25] != ele[17][25];
    ele[9][25] != ele[18][25];
    ele[9][25] != ele[19][25];
    ele[9][25] != ele[20][25];
    ele[9][25] != ele[21][25];
    ele[9][25] != ele[22][25];
    ele[9][25] != ele[23][25];
    ele[9][25] != ele[24][25];
    ele[9][25] != ele[25][25];
    ele[9][25] != ele[26][25];
    ele[9][25] != ele[27][25];
    ele[9][25] != ele[28][25];
    ele[9][25] != ele[29][25];
    ele[9][25] != ele[30][25];
    ele[9][25] != ele[31][25];
    ele[9][25] != ele[32][25];
    ele[9][25] != ele[33][25];
    ele[9][25] != ele[34][25];
    ele[9][25] != ele[35][25];
    ele[9][25] != ele[9][26];
    ele[9][25] != ele[9][27];
    ele[9][25] != ele[9][28];
    ele[9][25] != ele[9][29];
    ele[9][25] != ele[9][30];
    ele[9][25] != ele[9][31];
    ele[9][25] != ele[9][32];
    ele[9][25] != ele[9][33];
    ele[9][25] != ele[9][34];
    ele[9][25] != ele[9][35];
    ele[9][26] != ele[10][24];
    ele[9][26] != ele[10][25];
    ele[9][26] != ele[10][26];
    ele[9][26] != ele[10][27];
    ele[9][26] != ele[10][28];
    ele[9][26] != ele[10][29];
    ele[9][26] != ele[11][24];
    ele[9][26] != ele[11][25];
    ele[9][26] != ele[11][26];
    ele[9][26] != ele[11][27];
    ele[9][26] != ele[11][28];
    ele[9][26] != ele[11][29];
    ele[9][26] != ele[12][26];
    ele[9][26] != ele[13][26];
    ele[9][26] != ele[14][26];
    ele[9][26] != ele[15][26];
    ele[9][26] != ele[16][26];
    ele[9][26] != ele[17][26];
    ele[9][26] != ele[18][26];
    ele[9][26] != ele[19][26];
    ele[9][26] != ele[20][26];
    ele[9][26] != ele[21][26];
    ele[9][26] != ele[22][26];
    ele[9][26] != ele[23][26];
    ele[9][26] != ele[24][26];
    ele[9][26] != ele[25][26];
    ele[9][26] != ele[26][26];
    ele[9][26] != ele[27][26];
    ele[9][26] != ele[28][26];
    ele[9][26] != ele[29][26];
    ele[9][26] != ele[30][26];
    ele[9][26] != ele[31][26];
    ele[9][26] != ele[32][26];
    ele[9][26] != ele[33][26];
    ele[9][26] != ele[34][26];
    ele[9][26] != ele[35][26];
    ele[9][26] != ele[9][27];
    ele[9][26] != ele[9][28];
    ele[9][26] != ele[9][29];
    ele[9][26] != ele[9][30];
    ele[9][26] != ele[9][31];
    ele[9][26] != ele[9][32];
    ele[9][26] != ele[9][33];
    ele[9][26] != ele[9][34];
    ele[9][26] != ele[9][35];
    ele[9][27] != ele[10][24];
    ele[9][27] != ele[10][25];
    ele[9][27] != ele[10][26];
    ele[9][27] != ele[10][27];
    ele[9][27] != ele[10][28];
    ele[9][27] != ele[10][29];
    ele[9][27] != ele[11][24];
    ele[9][27] != ele[11][25];
    ele[9][27] != ele[11][26];
    ele[9][27] != ele[11][27];
    ele[9][27] != ele[11][28];
    ele[9][27] != ele[11][29];
    ele[9][27] != ele[12][27];
    ele[9][27] != ele[13][27];
    ele[9][27] != ele[14][27];
    ele[9][27] != ele[15][27];
    ele[9][27] != ele[16][27];
    ele[9][27] != ele[17][27];
    ele[9][27] != ele[18][27];
    ele[9][27] != ele[19][27];
    ele[9][27] != ele[20][27];
    ele[9][27] != ele[21][27];
    ele[9][27] != ele[22][27];
    ele[9][27] != ele[23][27];
    ele[9][27] != ele[24][27];
    ele[9][27] != ele[25][27];
    ele[9][27] != ele[26][27];
    ele[9][27] != ele[27][27];
    ele[9][27] != ele[28][27];
    ele[9][27] != ele[29][27];
    ele[9][27] != ele[30][27];
    ele[9][27] != ele[31][27];
    ele[9][27] != ele[32][27];
    ele[9][27] != ele[33][27];
    ele[9][27] != ele[34][27];
    ele[9][27] != ele[35][27];
    ele[9][27] != ele[9][28];
    ele[9][27] != ele[9][29];
    ele[9][27] != ele[9][30];
    ele[9][27] != ele[9][31];
    ele[9][27] != ele[9][32];
    ele[9][27] != ele[9][33];
    ele[9][27] != ele[9][34];
    ele[9][27] != ele[9][35];
    ele[9][28] != ele[10][24];
    ele[9][28] != ele[10][25];
    ele[9][28] != ele[10][26];
    ele[9][28] != ele[10][27];
    ele[9][28] != ele[10][28];
    ele[9][28] != ele[10][29];
    ele[9][28] != ele[11][24];
    ele[9][28] != ele[11][25];
    ele[9][28] != ele[11][26];
    ele[9][28] != ele[11][27];
    ele[9][28] != ele[11][28];
    ele[9][28] != ele[11][29];
    ele[9][28] != ele[12][28];
    ele[9][28] != ele[13][28];
    ele[9][28] != ele[14][28];
    ele[9][28] != ele[15][28];
    ele[9][28] != ele[16][28];
    ele[9][28] != ele[17][28];
    ele[9][28] != ele[18][28];
    ele[9][28] != ele[19][28];
    ele[9][28] != ele[20][28];
    ele[9][28] != ele[21][28];
    ele[9][28] != ele[22][28];
    ele[9][28] != ele[23][28];
    ele[9][28] != ele[24][28];
    ele[9][28] != ele[25][28];
    ele[9][28] != ele[26][28];
    ele[9][28] != ele[27][28];
    ele[9][28] != ele[28][28];
    ele[9][28] != ele[29][28];
    ele[9][28] != ele[30][28];
    ele[9][28] != ele[31][28];
    ele[9][28] != ele[32][28];
    ele[9][28] != ele[33][28];
    ele[9][28] != ele[34][28];
    ele[9][28] != ele[35][28];
    ele[9][28] != ele[9][29];
    ele[9][28] != ele[9][30];
    ele[9][28] != ele[9][31];
    ele[9][28] != ele[9][32];
    ele[9][28] != ele[9][33];
    ele[9][28] != ele[9][34];
    ele[9][28] != ele[9][35];
    ele[9][29] != ele[10][24];
    ele[9][29] != ele[10][25];
    ele[9][29] != ele[10][26];
    ele[9][29] != ele[10][27];
    ele[9][29] != ele[10][28];
    ele[9][29] != ele[10][29];
    ele[9][29] != ele[11][24];
    ele[9][29] != ele[11][25];
    ele[9][29] != ele[11][26];
    ele[9][29] != ele[11][27];
    ele[9][29] != ele[11][28];
    ele[9][29] != ele[11][29];
    ele[9][29] != ele[12][29];
    ele[9][29] != ele[13][29];
    ele[9][29] != ele[14][29];
    ele[9][29] != ele[15][29];
    ele[9][29] != ele[16][29];
    ele[9][29] != ele[17][29];
    ele[9][29] != ele[18][29];
    ele[9][29] != ele[19][29];
    ele[9][29] != ele[20][29];
    ele[9][29] != ele[21][29];
    ele[9][29] != ele[22][29];
    ele[9][29] != ele[23][29];
    ele[9][29] != ele[24][29];
    ele[9][29] != ele[25][29];
    ele[9][29] != ele[26][29];
    ele[9][29] != ele[27][29];
    ele[9][29] != ele[28][29];
    ele[9][29] != ele[29][29];
    ele[9][29] != ele[30][29];
    ele[9][29] != ele[31][29];
    ele[9][29] != ele[32][29];
    ele[9][29] != ele[33][29];
    ele[9][29] != ele[34][29];
    ele[9][29] != ele[35][29];
    ele[9][29] != ele[9][30];
    ele[9][29] != ele[9][31];
    ele[9][29] != ele[9][32];
    ele[9][29] != ele[9][33];
    ele[9][29] != ele[9][34];
    ele[9][29] != ele[9][35];
    ele[9][3] != ele[10][0];
    ele[9][3] != ele[10][1];
    ele[9][3] != ele[10][2];
    ele[9][3] != ele[10][3];
    ele[9][3] != ele[10][4];
    ele[9][3] != ele[10][5];
    ele[9][3] != ele[11][0];
    ele[9][3] != ele[11][1];
    ele[9][3] != ele[11][2];
    ele[9][3] != ele[11][3];
    ele[9][3] != ele[11][4];
    ele[9][3] != ele[11][5];
    ele[9][3] != ele[12][3];
    ele[9][3] != ele[13][3];
    ele[9][3] != ele[14][3];
    ele[9][3] != ele[15][3];
    ele[9][3] != ele[16][3];
    ele[9][3] != ele[17][3];
    ele[9][3] != ele[18][3];
    ele[9][3] != ele[19][3];
    ele[9][3] != ele[20][3];
    ele[9][3] != ele[21][3];
    ele[9][3] != ele[22][3];
    ele[9][3] != ele[23][3];
    ele[9][3] != ele[24][3];
    ele[9][3] != ele[25][3];
    ele[9][3] != ele[26][3];
    ele[9][3] != ele[27][3];
    ele[9][3] != ele[28][3];
    ele[9][3] != ele[29][3];
    ele[9][3] != ele[30][3];
    ele[9][3] != ele[31][3];
    ele[9][3] != ele[32][3];
    ele[9][3] != ele[33][3];
    ele[9][3] != ele[34][3];
    ele[9][3] != ele[35][3];
    ele[9][3] != ele[9][10];
    ele[9][3] != ele[9][11];
    ele[9][3] != ele[9][12];
    ele[9][3] != ele[9][13];
    ele[9][3] != ele[9][14];
    ele[9][3] != ele[9][15];
    ele[9][3] != ele[9][16];
    ele[9][3] != ele[9][17];
    ele[9][3] != ele[9][18];
    ele[9][3] != ele[9][19];
    ele[9][3] != ele[9][20];
    ele[9][3] != ele[9][21];
    ele[9][3] != ele[9][22];
    ele[9][3] != ele[9][23];
    ele[9][3] != ele[9][24];
    ele[9][3] != ele[9][25];
    ele[9][3] != ele[9][26];
    ele[9][3] != ele[9][27];
    ele[9][3] != ele[9][28];
    ele[9][3] != ele[9][29];
    ele[9][3] != ele[9][30];
    ele[9][3] != ele[9][31];
    ele[9][3] != ele[9][32];
    ele[9][3] != ele[9][33];
    ele[9][3] != ele[9][34];
    ele[9][3] != ele[9][35];
    ele[9][3] != ele[9][4];
    ele[9][3] != ele[9][5];
    ele[9][3] != ele[9][6];
    ele[9][3] != ele[9][7];
    ele[9][3] != ele[9][8];
    ele[9][3] != ele[9][9];
    ele[9][30] != ele[10][30];
    ele[9][30] != ele[10][31];
    ele[9][30] != ele[10][32];
    ele[9][30] != ele[10][33];
    ele[9][30] != ele[10][34];
    ele[9][30] != ele[10][35];
    ele[9][30] != ele[11][30];
    ele[9][30] != ele[11][31];
    ele[9][30] != ele[11][32];
    ele[9][30] != ele[11][33];
    ele[9][30] != ele[11][34];
    ele[9][30] != ele[11][35];
    ele[9][30] != ele[12][30];
    ele[9][30] != ele[13][30];
    ele[9][30] != ele[14][30];
    ele[9][30] != ele[15][30];
    ele[9][30] != ele[16][30];
    ele[9][30] != ele[17][30];
    ele[9][30] != ele[18][30];
    ele[9][30] != ele[19][30];
    ele[9][30] != ele[20][30];
    ele[9][30] != ele[21][30];
    ele[9][30] != ele[22][30];
    ele[9][30] != ele[23][30];
    ele[9][30] != ele[24][30];
    ele[9][30] != ele[25][30];
    ele[9][30] != ele[26][30];
    ele[9][30] != ele[27][30];
    ele[9][30] != ele[28][30];
    ele[9][30] != ele[29][30];
    ele[9][30] != ele[30][30];
    ele[9][30] != ele[31][30];
    ele[9][30] != ele[32][30];
    ele[9][30] != ele[33][30];
    ele[9][30] != ele[34][30];
    ele[9][30] != ele[35][30];
    ele[9][30] != ele[9][31];
    ele[9][30] != ele[9][32];
    ele[9][30] != ele[9][33];
    ele[9][30] != ele[9][34];
    ele[9][30] != ele[9][35];
    ele[9][31] != ele[10][30];
    ele[9][31] != ele[10][31];
    ele[9][31] != ele[10][32];
    ele[9][31] != ele[10][33];
    ele[9][31] != ele[10][34];
    ele[9][31] != ele[10][35];
    ele[9][31] != ele[11][30];
    ele[9][31] != ele[11][31];
    ele[9][31] != ele[11][32];
    ele[9][31] != ele[11][33];
    ele[9][31] != ele[11][34];
    ele[9][31] != ele[11][35];
    ele[9][31] != ele[12][31];
    ele[9][31] != ele[13][31];
    ele[9][31] != ele[14][31];
    ele[9][31] != ele[15][31];
    ele[9][31] != ele[16][31];
    ele[9][31] != ele[17][31];
    ele[9][31] != ele[18][31];
    ele[9][31] != ele[19][31];
    ele[9][31] != ele[20][31];
    ele[9][31] != ele[21][31];
    ele[9][31] != ele[22][31];
    ele[9][31] != ele[23][31];
    ele[9][31] != ele[24][31];
    ele[9][31] != ele[25][31];
    ele[9][31] != ele[26][31];
    ele[9][31] != ele[27][31];
    ele[9][31] != ele[28][31];
    ele[9][31] != ele[29][31];
    ele[9][31] != ele[30][31];
    ele[9][31] != ele[31][31];
    ele[9][31] != ele[32][31];
    ele[9][31] != ele[33][31];
    ele[9][31] != ele[34][31];
    ele[9][31] != ele[35][31];
    ele[9][31] != ele[9][32];
    ele[9][31] != ele[9][33];
    ele[9][31] != ele[9][34];
    ele[9][31] != ele[9][35];
    ele[9][32] != ele[10][30];
    ele[9][32] != ele[10][31];
    ele[9][32] != ele[10][32];
    ele[9][32] != ele[10][33];
    ele[9][32] != ele[10][34];
    ele[9][32] != ele[10][35];
    ele[9][32] != ele[11][30];
    ele[9][32] != ele[11][31];
    ele[9][32] != ele[11][32];
    ele[9][32] != ele[11][33];
    ele[9][32] != ele[11][34];
    ele[9][32] != ele[11][35];
    ele[9][32] != ele[12][32];
    ele[9][32] != ele[13][32];
    ele[9][32] != ele[14][32];
    ele[9][32] != ele[15][32];
    ele[9][32] != ele[16][32];
    ele[9][32] != ele[17][32];
    ele[9][32] != ele[18][32];
    ele[9][32] != ele[19][32];
    ele[9][32] != ele[20][32];
    ele[9][32] != ele[21][32];
    ele[9][32] != ele[22][32];
    ele[9][32] != ele[23][32];
    ele[9][32] != ele[24][32];
    ele[9][32] != ele[25][32];
    ele[9][32] != ele[26][32];
    ele[9][32] != ele[27][32];
    ele[9][32] != ele[28][32];
    ele[9][32] != ele[29][32];
    ele[9][32] != ele[30][32];
    ele[9][32] != ele[31][32];
    ele[9][32] != ele[32][32];
    ele[9][32] != ele[33][32];
    ele[9][32] != ele[34][32];
    ele[9][32] != ele[35][32];
    ele[9][32] != ele[9][33];
    ele[9][32] != ele[9][34];
    ele[9][32] != ele[9][35];
    ele[9][33] != ele[10][30];
    ele[9][33] != ele[10][31];
    ele[9][33] != ele[10][32];
    ele[9][33] != ele[10][33];
    ele[9][33] != ele[10][34];
    ele[9][33] != ele[10][35];
    ele[9][33] != ele[11][30];
    ele[9][33] != ele[11][31];
    ele[9][33] != ele[11][32];
    ele[9][33] != ele[11][33];
    ele[9][33] != ele[11][34];
    ele[9][33] != ele[11][35];
    ele[9][33] != ele[12][33];
    ele[9][33] != ele[13][33];
    ele[9][33] != ele[14][33];
    ele[9][33] != ele[15][33];
    ele[9][33] != ele[16][33];
    ele[9][33] != ele[17][33];
    ele[9][33] != ele[18][33];
    ele[9][33] != ele[19][33];
    ele[9][33] != ele[20][33];
    ele[9][33] != ele[21][33];
    ele[9][33] != ele[22][33];
    ele[9][33] != ele[23][33];
    ele[9][33] != ele[24][33];
    ele[9][33] != ele[25][33];
    ele[9][33] != ele[26][33];
    ele[9][33] != ele[27][33];
    ele[9][33] != ele[28][33];
    ele[9][33] != ele[29][33];
    ele[9][33] != ele[30][33];
    ele[9][33] != ele[31][33];
    ele[9][33] != ele[32][33];
    ele[9][33] != ele[33][33];
    ele[9][33] != ele[34][33];
    ele[9][33] != ele[35][33];
    ele[9][33] != ele[9][34];
    ele[9][33] != ele[9][35];
    ele[9][34] != ele[10][30];
    ele[9][34] != ele[10][31];
    ele[9][34] != ele[10][32];
    ele[9][34] != ele[10][33];
    ele[9][34] != ele[10][34];
    ele[9][34] != ele[10][35];
    ele[9][34] != ele[11][30];
    ele[9][34] != ele[11][31];
    ele[9][34] != ele[11][32];
    ele[9][34] != ele[11][33];
    ele[9][34] != ele[11][34];
    ele[9][34] != ele[11][35];
    ele[9][34] != ele[12][34];
    ele[9][34] != ele[13][34];
    ele[9][34] != ele[14][34];
    ele[9][34] != ele[15][34];
    ele[9][34] != ele[16][34];
    ele[9][34] != ele[17][34];
    ele[9][34] != ele[18][34];
    ele[9][34] != ele[19][34];
    ele[9][34] != ele[20][34];
    ele[9][34] != ele[21][34];
    ele[9][34] != ele[22][34];
    ele[9][34] != ele[23][34];
    ele[9][34] != ele[24][34];
    ele[9][34] != ele[25][34];
    ele[9][34] != ele[26][34];
    ele[9][34] != ele[27][34];
    ele[9][34] != ele[28][34];
    ele[9][34] != ele[29][34];
    ele[9][34] != ele[30][34];
    ele[9][34] != ele[31][34];
    ele[9][34] != ele[32][34];
    ele[9][34] != ele[33][34];
    ele[9][34] != ele[34][34];
    ele[9][34] != ele[35][34];
    ele[9][34] != ele[9][35];
    ele[9][35] != ele[10][30];
    ele[9][35] != ele[10][31];
    ele[9][35] != ele[10][32];
    ele[9][35] != ele[10][33];
    ele[9][35] != ele[10][34];
    ele[9][35] != ele[10][35];
    ele[9][35] != ele[11][30];
    ele[9][35] != ele[11][31];
    ele[9][35] != ele[11][32];
    ele[9][35] != ele[11][33];
    ele[9][35] != ele[11][34];
    ele[9][35] != ele[11][35];
    ele[9][35] != ele[12][35];
    ele[9][35] != ele[13][35];
    ele[9][35] != ele[14][35];
    ele[9][35] != ele[15][35];
    ele[9][35] != ele[16][35];
    ele[9][35] != ele[17][35];
    ele[9][35] != ele[18][35];
    ele[9][35] != ele[19][35];
    ele[9][35] != ele[20][35];
    ele[9][35] != ele[21][35];
    ele[9][35] != ele[22][35];
    ele[9][35] != ele[23][35];
    ele[9][35] != ele[24][35];
    ele[9][35] != ele[25][35];
    ele[9][35] != ele[26][35];
    ele[9][35] != ele[27][35];
    ele[9][35] != ele[28][35];
    ele[9][35] != ele[29][35];
    ele[9][35] != ele[30][35];
    ele[9][35] != ele[31][35];
    ele[9][35] != ele[32][35];
    ele[9][35] != ele[33][35];
    ele[9][35] != ele[34][35];
    ele[9][35] != ele[35][35];
    ele[9][4] != ele[10][0];
    ele[9][4] != ele[10][1];
    ele[9][4] != ele[10][2];
    ele[9][4] != ele[10][3];
    ele[9][4] != ele[10][4];
    ele[9][4] != ele[10][5];
    ele[9][4] != ele[11][0];
    ele[9][4] != ele[11][1];
    ele[9][4] != ele[11][2];
    ele[9][4] != ele[11][3];
    ele[9][4] != ele[11][4];
    ele[9][4] != ele[11][5];
    ele[9][4] != ele[12][4];
    ele[9][4] != ele[13][4];
    ele[9][4] != ele[14][4];
    ele[9][4] != ele[15][4];
    ele[9][4] != ele[16][4];
    ele[9][4] != ele[17][4];
    ele[9][4] != ele[18][4];
    ele[9][4] != ele[19][4];
    ele[9][4] != ele[20][4];
    ele[9][4] != ele[21][4];
    ele[9][4] != ele[22][4];
    ele[9][4] != ele[23][4];
    ele[9][4] != ele[24][4];
    ele[9][4] != ele[25][4];
    ele[9][4] != ele[26][4];
    ele[9][4] != ele[27][4];
    ele[9][4] != ele[28][4];
    ele[9][4] != ele[29][4];
    ele[9][4] != ele[30][4];
    ele[9][4] != ele[31][4];
    ele[9][4] != ele[32][4];
    ele[9][4] != ele[33][4];
    ele[9][4] != ele[34][4];
    ele[9][4] != ele[35][4];
    ele[9][4] != ele[9][10];
    ele[9][4] != ele[9][11];
    ele[9][4] != ele[9][12];
    ele[9][4] != ele[9][13];
    ele[9][4] != ele[9][14];
    ele[9][4] != ele[9][15];
    ele[9][4] != ele[9][16];
    ele[9][4] != ele[9][17];
    ele[9][4] != ele[9][18];
    ele[9][4] != ele[9][19];
    ele[9][4] != ele[9][20];
    ele[9][4] != ele[9][21];
    ele[9][4] != ele[9][22];
    ele[9][4] != ele[9][23];
    ele[9][4] != ele[9][24];
    ele[9][4] != ele[9][25];
    ele[9][4] != ele[9][26];
    ele[9][4] != ele[9][27];
    ele[9][4] != ele[9][28];
    ele[9][4] != ele[9][29];
    ele[9][4] != ele[9][30];
    ele[9][4] != ele[9][31];
    ele[9][4] != ele[9][32];
    ele[9][4] != ele[9][33];
    ele[9][4] != ele[9][34];
    ele[9][4] != ele[9][35];
    ele[9][4] != ele[9][5];
    ele[9][4] != ele[9][6];
    ele[9][4] != ele[9][7];
    ele[9][4] != ele[9][8];
    ele[9][4] != ele[9][9];
    ele[9][5] != ele[10][0];
    ele[9][5] != ele[10][1];
    ele[9][5] != ele[10][2];
    ele[9][5] != ele[10][3];
    ele[9][5] != ele[10][4];
    ele[9][5] != ele[10][5];
    ele[9][5] != ele[11][0];
    ele[9][5] != ele[11][1];
    ele[9][5] != ele[11][2];
    ele[9][5] != ele[11][3];
    ele[9][5] != ele[11][4];
    ele[9][5] != ele[11][5];
    ele[9][5] != ele[12][5];
    ele[9][5] != ele[13][5];
    ele[9][5] != ele[14][5];
    ele[9][5] != ele[15][5];
    ele[9][5] != ele[16][5];
    ele[9][5] != ele[17][5];
    ele[9][5] != ele[18][5];
    ele[9][5] != ele[19][5];
    ele[9][5] != ele[20][5];
    ele[9][5] != ele[21][5];
    ele[9][5] != ele[22][5];
    ele[9][5] != ele[23][5];
    ele[9][5] != ele[24][5];
    ele[9][5] != ele[25][5];
    ele[9][5] != ele[26][5];
    ele[9][5] != ele[27][5];
    ele[9][5] != ele[28][5];
    ele[9][5] != ele[29][5];
    ele[9][5] != ele[30][5];
    ele[9][5] != ele[31][5];
    ele[9][5] != ele[32][5];
    ele[9][5] != ele[33][5];
    ele[9][5] != ele[34][5];
    ele[9][5] != ele[35][5];
    ele[9][5] != ele[9][10];
    ele[9][5] != ele[9][11];
    ele[9][5] != ele[9][12];
    ele[9][5] != ele[9][13];
    ele[9][5] != ele[9][14];
    ele[9][5] != ele[9][15];
    ele[9][5] != ele[9][16];
    ele[9][5] != ele[9][17];
    ele[9][5] != ele[9][18];
    ele[9][5] != ele[9][19];
    ele[9][5] != ele[9][20];
    ele[9][5] != ele[9][21];
    ele[9][5] != ele[9][22];
    ele[9][5] != ele[9][23];
    ele[9][5] != ele[9][24];
    ele[9][5] != ele[9][25];
    ele[9][5] != ele[9][26];
    ele[9][5] != ele[9][27];
    ele[9][5] != ele[9][28];
    ele[9][5] != ele[9][29];
    ele[9][5] != ele[9][30];
    ele[9][5] != ele[9][31];
    ele[9][5] != ele[9][32];
    ele[9][5] != ele[9][33];
    ele[9][5] != ele[9][34];
    ele[9][5] != ele[9][35];
    ele[9][5] != ele[9][6];
    ele[9][5] != ele[9][7];
    ele[9][5] != ele[9][8];
    ele[9][5] != ele[9][9];
    ele[9][6] != ele[10][10];
    ele[9][6] != ele[10][11];
    ele[9][6] != ele[10][6];
    ele[9][6] != ele[10][7];
    ele[9][6] != ele[10][8];
    ele[9][6] != ele[10][9];
    ele[9][6] != ele[11][10];
    ele[9][6] != ele[11][11];
    ele[9][6] != ele[11][6];
    ele[9][6] != ele[11][7];
    ele[9][6] != ele[11][8];
    ele[9][6] != ele[11][9];
    ele[9][6] != ele[12][6];
    ele[9][6] != ele[13][6];
    ele[9][6] != ele[14][6];
    ele[9][6] != ele[15][6];
    ele[9][6] != ele[16][6];
    ele[9][6] != ele[17][6];
    ele[9][6] != ele[18][6];
    ele[9][6] != ele[19][6];
    ele[9][6] != ele[20][6];
    ele[9][6] != ele[21][6];
    ele[9][6] != ele[22][6];
    ele[9][6] != ele[23][6];
    ele[9][6] != ele[24][6];
    ele[9][6] != ele[25][6];
    ele[9][6] != ele[26][6];
    ele[9][6] != ele[27][6];
    ele[9][6] != ele[28][6];
    ele[9][6] != ele[29][6];
    ele[9][6] != ele[30][6];
    ele[9][6] != ele[31][6];
    ele[9][6] != ele[32][6];
    ele[9][6] != ele[33][6];
    ele[9][6] != ele[34][6];
    ele[9][6] != ele[35][6];
    ele[9][6] != ele[9][10];
    ele[9][6] != ele[9][11];
    ele[9][6] != ele[9][12];
    ele[9][6] != ele[9][13];
    ele[9][6] != ele[9][14];
    ele[9][6] != ele[9][15];
    ele[9][6] != ele[9][16];
    ele[9][6] != ele[9][17];
    ele[9][6] != ele[9][18];
    ele[9][6] != ele[9][19];
    ele[9][6] != ele[9][20];
    ele[9][6] != ele[9][21];
    ele[9][6] != ele[9][22];
    ele[9][6] != ele[9][23];
    ele[9][6] != ele[9][24];
    ele[9][6] != ele[9][25];
    ele[9][6] != ele[9][26];
    ele[9][6] != ele[9][27];
    ele[9][6] != ele[9][28];
    ele[9][6] != ele[9][29];
    ele[9][6] != ele[9][30];
    ele[9][6] != ele[9][31];
    ele[9][6] != ele[9][32];
    ele[9][6] != ele[9][33];
    ele[9][6] != ele[9][34];
    ele[9][6] != ele[9][35];
    ele[9][6] != ele[9][7];
    ele[9][6] != ele[9][8];
    ele[9][6] != ele[9][9];
    ele[9][7] != ele[10][10];
    ele[9][7] != ele[10][11];
    ele[9][7] != ele[10][6];
    ele[9][7] != ele[10][7];
    ele[9][7] != ele[10][8];
    ele[9][7] != ele[10][9];
    ele[9][7] != ele[11][10];
    ele[9][7] != ele[11][11];
    ele[9][7] != ele[11][6];
    ele[9][7] != ele[11][7];
    ele[9][7] != ele[11][8];
    ele[9][7] != ele[11][9];
    ele[9][7] != ele[12][7];
    ele[9][7] != ele[13][7];
    ele[9][7] != ele[14][7];
    ele[9][7] != ele[15][7];
    ele[9][7] != ele[16][7];
    ele[9][7] != ele[17][7];
    ele[9][7] != ele[18][7];
    ele[9][7] != ele[19][7];
    ele[9][7] != ele[20][7];
    ele[9][7] != ele[21][7];
    ele[9][7] != ele[22][7];
    ele[9][7] != ele[23][7];
    ele[9][7] != ele[24][7];
    ele[9][7] != ele[25][7];
    ele[9][7] != ele[26][7];
    ele[9][7] != ele[27][7];
    ele[9][7] != ele[28][7];
    ele[9][7] != ele[29][7];
    ele[9][7] != ele[30][7];
    ele[9][7] != ele[31][7];
    ele[9][7] != ele[32][7];
    ele[9][7] != ele[33][7];
    ele[9][7] != ele[34][7];
    ele[9][7] != ele[35][7];
    ele[9][7] != ele[9][10];
    ele[9][7] != ele[9][11];
    ele[9][7] != ele[9][12];
    ele[9][7] != ele[9][13];
    ele[9][7] != ele[9][14];
    ele[9][7] != ele[9][15];
    ele[9][7] != ele[9][16];
    ele[9][7] != ele[9][17];
    ele[9][7] != ele[9][18];
    ele[9][7] != ele[9][19];
    ele[9][7] != ele[9][20];
    ele[9][7] != ele[9][21];
    ele[9][7] != ele[9][22];
    ele[9][7] != ele[9][23];
    ele[9][7] != ele[9][24];
    ele[9][7] != ele[9][25];
    ele[9][7] != ele[9][26];
    ele[9][7] != ele[9][27];
    ele[9][7] != ele[9][28];
    ele[9][7] != ele[9][29];
    ele[9][7] != ele[9][30];
    ele[9][7] != ele[9][31];
    ele[9][7] != ele[9][32];
    ele[9][7] != ele[9][33];
    ele[9][7] != ele[9][34];
    ele[9][7] != ele[9][35];
    ele[9][7] != ele[9][8];
    ele[9][7] != ele[9][9];
    ele[9][8] != ele[10][10];
    ele[9][8] != ele[10][11];
    ele[9][8] != ele[10][6];
    ele[9][8] != ele[10][7];
    ele[9][8] != ele[10][8];
    ele[9][8] != ele[10][9];
    ele[9][8] != ele[11][10];
    ele[9][8] != ele[11][11];
    ele[9][8] != ele[11][6];
    ele[9][8] != ele[11][7];
    ele[9][8] != ele[11][8];
    ele[9][8] != ele[11][9];
    ele[9][8] != ele[12][8];
    ele[9][8] != ele[13][8];
    ele[9][8] != ele[14][8];
    ele[9][8] != ele[15][8];
    ele[9][8] != ele[16][8];
    ele[9][8] != ele[17][8];
    ele[9][8] != ele[18][8];
    ele[9][8] != ele[19][8];
    ele[9][8] != ele[20][8];
    ele[9][8] != ele[21][8];
    ele[9][8] != ele[22][8];
    ele[9][8] != ele[23][8];
    ele[9][8] != ele[24][8];
    ele[9][8] != ele[25][8];
    ele[9][8] != ele[26][8];
    ele[9][8] != ele[27][8];
    ele[9][8] != ele[28][8];
    ele[9][8] != ele[29][8];
    ele[9][8] != ele[30][8];
    ele[9][8] != ele[31][8];
    ele[9][8] != ele[32][8];
    ele[9][8] != ele[33][8];
    ele[9][8] != ele[34][8];
    ele[9][8] != ele[35][8];
    ele[9][8] != ele[9][10];
    ele[9][8] != ele[9][11];
    ele[9][8] != ele[9][12];
    ele[9][8] != ele[9][13];
    ele[9][8] != ele[9][14];
    ele[9][8] != ele[9][15];
    ele[9][8] != ele[9][16];
    ele[9][8] != ele[9][17];
    ele[9][8] != ele[9][18];
    ele[9][8] != ele[9][19];
    ele[9][8] != ele[9][20];
    ele[9][8] != ele[9][21];
    ele[9][8] != ele[9][22];
    ele[9][8] != ele[9][23];
    ele[9][8] != ele[9][24];
    ele[9][8] != ele[9][25];
    ele[9][8] != ele[9][26];
    ele[9][8] != ele[9][27];
    ele[9][8] != ele[9][28];
    ele[9][8] != ele[9][29];
    ele[9][8] != ele[9][30];
    ele[9][8] != ele[9][31];
    ele[9][8] != ele[9][32];
    ele[9][8] != ele[9][33];
    ele[9][8] != ele[9][34];
    ele[9][8] != ele[9][35];
    ele[9][8] != ele[9][9];
    ele[9][9] != ele[10][10];
    ele[9][9] != ele[10][11];
    ele[9][9] != ele[10][6];
    ele[9][9] != ele[10][7];
    ele[9][9] != ele[10][8];
    ele[9][9] != ele[10][9];
    ele[9][9] != ele[11][10];
    ele[9][9] != ele[11][11];
    ele[9][9] != ele[11][6];
    ele[9][9] != ele[11][7];
    ele[9][9] != ele[11][8];
    ele[9][9] != ele[11][9];
    ele[9][9] != ele[12][9];
    ele[9][9] != ele[13][9];
    ele[9][9] != ele[14][9];
    ele[9][9] != ele[15][9];
    ele[9][9] != ele[16][9];
    ele[9][9] != ele[17][9];
    ele[9][9] != ele[18][9];
    ele[9][9] != ele[19][9];
    ele[9][9] != ele[20][9];
    ele[9][9] != ele[21][9];
    ele[9][9] != ele[22][9];
    ele[9][9] != ele[23][9];
    ele[9][9] != ele[24][9];
    ele[9][9] != ele[25][9];
    ele[9][9] != ele[26][9];
    ele[9][9] != ele[27][9];
    ele[9][9] != ele[28][9];
    ele[9][9] != ele[29][9];
    ele[9][9] != ele[30][9];
    ele[9][9] != ele[31][9];
    ele[9][9] != ele[32][9];
    ele[9][9] != ele[33][9];
    ele[9][9] != ele[34][9];
    ele[9][9] != ele[35][9];
    ele[9][9] != ele[9][10];
    ele[9][9] != ele[9][11];
    ele[9][9] != ele[9][12];
    ele[9][9] != ele[9][13];
    ele[9][9] != ele[9][14];
    ele[9][9] != ele[9][15];
    ele[9][9] != ele[9][16];
    ele[9][9] != ele[9][17];
    ele[9][9] != ele[9][18];
    ele[9][9] != ele[9][19];
    ele[9][9] != ele[9][20];
    ele[9][9] != ele[9][21];
    ele[9][9] != ele[9][22];
    ele[9][9] != ele[9][23];
    ele[9][9] != ele[9][24];
    ele[9][9] != ele[9][25];
    ele[9][9] != ele[9][26];
    ele[9][9] != ele[9][27];
    ele[9][9] != ele[9][28];
    ele[9][9] != ele[9][29];
    ele[9][9] != ele[9][30];
    ele[9][9] != ele[9][31];
    ele[9][9] != ele[9][32];
    ele[9][9] != ele[9][33];
    ele[9][9] != ele[9][34];
    ele[9][9] != ele[9][35];
  // NUMBER OF CONSTRAINTS: 61560
  }
  function new ();
    if (! this.randomize ()) begin
      $display ("ERROR: Randomization failed...!!!");
    end
  endfunction: new
  function show ();
    $display (ele[0][0], ele[0][1], ele[0][2], ele[0][3], ele[0][4], ele[0][5], ele[0][6], ele[0][7], ele[0][8], ele[0][9], ele[0][10], ele[0][11], ele[0][12], ele[0][13], ele[0][14], ele[0][15], ele[0][16], ele[0][17], ele[0][18], ele[0][19], ele[0][20], ele[0][21], ele[0][22], ele[0][23], ele[0][24], ele[0][25], ele[0][26], ele[0][27], ele[0][28], ele[0][29], ele[0][30], ele[0][31], ele[0][32], ele[0][33], ele[0][34], ele[0][35]);
    $display (ele[1][0], ele[1][1], ele[1][2], ele[1][3], ele[1][4], ele[1][5], ele[1][6], ele[1][7], ele[1][8], ele[1][9], ele[1][10], ele[1][11], ele[1][12], ele[1][13], ele[1][14], ele[1][15], ele[1][16], ele[1][17], ele[1][18], ele[1][19], ele[1][20], ele[1][21], ele[1][22], ele[1][23], ele[1][24], ele[1][25], ele[1][26], ele[1][27], ele[1][28], ele[1][29], ele[1][30], ele[1][31], ele[1][32], ele[1][33], ele[1][34], ele[1][35]);
    $display (ele[2][0], ele[2][1], ele[2][2], ele[2][3], ele[2][4], ele[2][5], ele[2][6], ele[2][7], ele[2][8], ele[2][9], ele[2][10], ele[2][11], ele[2][12], ele[2][13], ele[2][14], ele[2][15], ele[2][16], ele[2][17], ele[2][18], ele[2][19], ele[2][20], ele[2][21], ele[2][22], ele[2][23], ele[2][24], ele[2][25], ele[2][26], ele[2][27], ele[2][28], ele[2][29], ele[2][30], ele[2][31], ele[2][32], ele[2][33], ele[2][34], ele[2][35]);
    $display (ele[3][0], ele[3][1], ele[3][2], ele[3][3], ele[3][4], ele[3][5], ele[3][6], ele[3][7], ele[3][8], ele[3][9], ele[3][10], ele[3][11], ele[3][12], ele[3][13], ele[3][14], ele[3][15], ele[3][16], ele[3][17], ele[3][18], ele[3][19], ele[3][20], ele[3][21], ele[3][22], ele[3][23], ele[3][24], ele[3][25], ele[3][26], ele[3][27], ele[3][28], ele[3][29], ele[3][30], ele[3][31], ele[3][32], ele[3][33], ele[3][34], ele[3][35]);
    $display (ele[4][0], ele[4][1], ele[4][2], ele[4][3], ele[4][4], ele[4][5], ele[4][6], ele[4][7], ele[4][8], ele[4][9], ele[4][10], ele[4][11], ele[4][12], ele[4][13], ele[4][14], ele[4][15], ele[4][16], ele[4][17], ele[4][18], ele[4][19], ele[4][20], ele[4][21], ele[4][22], ele[4][23], ele[4][24], ele[4][25], ele[4][26], ele[4][27], ele[4][28], ele[4][29], ele[4][30], ele[4][31], ele[4][32], ele[4][33], ele[4][34], ele[4][35]);
    $display (ele[5][0], ele[5][1], ele[5][2], ele[5][3], ele[5][4], ele[5][5], ele[5][6], ele[5][7], ele[5][8], ele[5][9], ele[5][10], ele[5][11], ele[5][12], ele[5][13], ele[5][14], ele[5][15], ele[5][16], ele[5][17], ele[5][18], ele[5][19], ele[5][20], ele[5][21], ele[5][22], ele[5][23], ele[5][24], ele[5][25], ele[5][26], ele[5][27], ele[5][28], ele[5][29], ele[5][30], ele[5][31], ele[5][32], ele[5][33], ele[5][34], ele[5][35]);
    $display (ele[6][0], ele[6][1], ele[6][2], ele[6][3], ele[6][4], ele[6][5], ele[6][6], ele[6][7], ele[6][8], ele[6][9], ele[6][10], ele[6][11], ele[6][12], ele[6][13], ele[6][14], ele[6][15], ele[6][16], ele[6][17], ele[6][18], ele[6][19], ele[6][20], ele[6][21], ele[6][22], ele[6][23], ele[6][24], ele[6][25], ele[6][26], ele[6][27], ele[6][28], ele[6][29], ele[6][30], ele[6][31], ele[6][32], ele[6][33], ele[6][34], ele[6][35]);
    $display (ele[7][0], ele[7][1], ele[7][2], ele[7][3], ele[7][4], ele[7][5], ele[7][6], ele[7][7], ele[7][8], ele[7][9], ele[7][10], ele[7][11], ele[7][12], ele[7][13], ele[7][14], ele[7][15], ele[7][16], ele[7][17], ele[7][18], ele[7][19], ele[7][20], ele[7][21], ele[7][22], ele[7][23], ele[7][24], ele[7][25], ele[7][26], ele[7][27], ele[7][28], ele[7][29], ele[7][30], ele[7][31], ele[7][32], ele[7][33], ele[7][34], ele[7][35]);
    $display (ele[8][0], ele[8][1], ele[8][2], ele[8][3], ele[8][4], ele[8][5], ele[8][6], ele[8][7], ele[8][8], ele[8][9], ele[8][10], ele[8][11], ele[8][12], ele[8][13], ele[8][14], ele[8][15], ele[8][16], ele[8][17], ele[8][18], ele[8][19], ele[8][20], ele[8][21], ele[8][22], ele[8][23], ele[8][24], ele[8][25], ele[8][26], ele[8][27], ele[8][28], ele[8][29], ele[8][30], ele[8][31], ele[8][32], ele[8][33], ele[8][34], ele[8][35]);
    $display (ele[9][0], ele[9][1], ele[9][2], ele[9][3], ele[9][4], ele[9][5], ele[9][6], ele[9][7], ele[9][8], ele[9][9], ele[9][10], ele[9][11], ele[9][12], ele[9][13], ele[9][14], ele[9][15], ele[9][16], ele[9][17], ele[9][18], ele[9][19], ele[9][20], ele[9][21], ele[9][22], ele[9][23], ele[9][24], ele[9][25], ele[9][26], ele[9][27], ele[9][28], ele[9][29], ele[9][30], ele[9][31], ele[9][32], ele[9][33], ele[9][34], ele[9][35]);
    $display (ele[10][0], ele[10][1], ele[10][2], ele[10][3], ele[10][4], ele[10][5], ele[10][6], ele[10][7], ele[10][8], ele[10][9], ele[10][10], ele[10][11], ele[10][12], ele[10][13], ele[10][14], ele[10][15], ele[10][16], ele[10][17], ele[10][18], ele[10][19], ele[10][20], ele[10][21], ele[10][22], ele[10][23], ele[10][24], ele[10][25], ele[10][26], ele[10][27], ele[10][28], ele[10][29], ele[10][30], ele[10][31], ele[10][32], ele[10][33], ele[10][34], ele[10][35]);
    $display (ele[11][0], ele[11][1], ele[11][2], ele[11][3], ele[11][4], ele[11][5], ele[11][6], ele[11][7], ele[11][8], ele[11][9], ele[11][10], ele[11][11], ele[11][12], ele[11][13], ele[11][14], ele[11][15], ele[11][16], ele[11][17], ele[11][18], ele[11][19], ele[11][20], ele[11][21], ele[11][22], ele[11][23], ele[11][24], ele[11][25], ele[11][26], ele[11][27], ele[11][28], ele[11][29], ele[11][30], ele[11][31], ele[11][32], ele[11][33], ele[11][34], ele[11][35]);
    $display (ele[12][0], ele[12][1], ele[12][2], ele[12][3], ele[12][4], ele[12][5], ele[12][6], ele[12][7], ele[12][8], ele[12][9], ele[12][10], ele[12][11], ele[12][12], ele[12][13], ele[12][14], ele[12][15], ele[12][16], ele[12][17], ele[12][18], ele[12][19], ele[12][20], ele[12][21], ele[12][22], ele[12][23], ele[12][24], ele[12][25], ele[12][26], ele[12][27], ele[12][28], ele[12][29], ele[12][30], ele[12][31], ele[12][32], ele[12][33], ele[12][34], ele[12][35]);
    $display (ele[13][0], ele[13][1], ele[13][2], ele[13][3], ele[13][4], ele[13][5], ele[13][6], ele[13][7], ele[13][8], ele[13][9], ele[13][10], ele[13][11], ele[13][12], ele[13][13], ele[13][14], ele[13][15], ele[13][16], ele[13][17], ele[13][18], ele[13][19], ele[13][20], ele[13][21], ele[13][22], ele[13][23], ele[13][24], ele[13][25], ele[13][26], ele[13][27], ele[13][28], ele[13][29], ele[13][30], ele[13][31], ele[13][32], ele[13][33], ele[13][34], ele[13][35]);
    $display (ele[14][0], ele[14][1], ele[14][2], ele[14][3], ele[14][4], ele[14][5], ele[14][6], ele[14][7], ele[14][8], ele[14][9], ele[14][10], ele[14][11], ele[14][12], ele[14][13], ele[14][14], ele[14][15], ele[14][16], ele[14][17], ele[14][18], ele[14][19], ele[14][20], ele[14][21], ele[14][22], ele[14][23], ele[14][24], ele[14][25], ele[14][26], ele[14][27], ele[14][28], ele[14][29], ele[14][30], ele[14][31], ele[14][32], ele[14][33], ele[14][34], ele[14][35]);
    $display (ele[15][0], ele[15][1], ele[15][2], ele[15][3], ele[15][4], ele[15][5], ele[15][6], ele[15][7], ele[15][8], ele[15][9], ele[15][10], ele[15][11], ele[15][12], ele[15][13], ele[15][14], ele[15][15], ele[15][16], ele[15][17], ele[15][18], ele[15][19], ele[15][20], ele[15][21], ele[15][22], ele[15][23], ele[15][24], ele[15][25], ele[15][26], ele[15][27], ele[15][28], ele[15][29], ele[15][30], ele[15][31], ele[15][32], ele[15][33], ele[15][34], ele[15][35]);
    $display (ele[16][0], ele[16][1], ele[16][2], ele[16][3], ele[16][4], ele[16][5], ele[16][6], ele[16][7], ele[16][8], ele[16][9], ele[16][10], ele[16][11], ele[16][12], ele[16][13], ele[16][14], ele[16][15], ele[16][16], ele[16][17], ele[16][18], ele[16][19], ele[16][20], ele[16][21], ele[16][22], ele[16][23], ele[16][24], ele[16][25], ele[16][26], ele[16][27], ele[16][28], ele[16][29], ele[16][30], ele[16][31], ele[16][32], ele[16][33], ele[16][34], ele[16][35]);
    $display (ele[17][0], ele[17][1], ele[17][2], ele[17][3], ele[17][4], ele[17][5], ele[17][6], ele[17][7], ele[17][8], ele[17][9], ele[17][10], ele[17][11], ele[17][12], ele[17][13], ele[17][14], ele[17][15], ele[17][16], ele[17][17], ele[17][18], ele[17][19], ele[17][20], ele[17][21], ele[17][22], ele[17][23], ele[17][24], ele[17][25], ele[17][26], ele[17][27], ele[17][28], ele[17][29], ele[17][30], ele[17][31], ele[17][32], ele[17][33], ele[17][34], ele[17][35]);
    $display (ele[18][0], ele[18][1], ele[18][2], ele[18][3], ele[18][4], ele[18][5], ele[18][6], ele[18][7], ele[18][8], ele[18][9], ele[18][10], ele[18][11], ele[18][12], ele[18][13], ele[18][14], ele[18][15], ele[18][16], ele[18][17], ele[18][18], ele[18][19], ele[18][20], ele[18][21], ele[18][22], ele[18][23], ele[18][24], ele[18][25], ele[18][26], ele[18][27], ele[18][28], ele[18][29], ele[18][30], ele[18][31], ele[18][32], ele[18][33], ele[18][34], ele[18][35]);
    $display (ele[19][0], ele[19][1], ele[19][2], ele[19][3], ele[19][4], ele[19][5], ele[19][6], ele[19][7], ele[19][8], ele[19][9], ele[19][10], ele[19][11], ele[19][12], ele[19][13], ele[19][14], ele[19][15], ele[19][16], ele[19][17], ele[19][18], ele[19][19], ele[19][20], ele[19][21], ele[19][22], ele[19][23], ele[19][24], ele[19][25], ele[19][26], ele[19][27], ele[19][28], ele[19][29], ele[19][30], ele[19][31], ele[19][32], ele[19][33], ele[19][34], ele[19][35]);
    $display (ele[20][0], ele[20][1], ele[20][2], ele[20][3], ele[20][4], ele[20][5], ele[20][6], ele[20][7], ele[20][8], ele[20][9], ele[20][10], ele[20][11], ele[20][12], ele[20][13], ele[20][14], ele[20][15], ele[20][16], ele[20][17], ele[20][18], ele[20][19], ele[20][20], ele[20][21], ele[20][22], ele[20][23], ele[20][24], ele[20][25], ele[20][26], ele[20][27], ele[20][28], ele[20][29], ele[20][30], ele[20][31], ele[20][32], ele[20][33], ele[20][34], ele[20][35]);
    $display (ele[21][0], ele[21][1], ele[21][2], ele[21][3], ele[21][4], ele[21][5], ele[21][6], ele[21][7], ele[21][8], ele[21][9], ele[21][10], ele[21][11], ele[21][12], ele[21][13], ele[21][14], ele[21][15], ele[21][16], ele[21][17], ele[21][18], ele[21][19], ele[21][20], ele[21][21], ele[21][22], ele[21][23], ele[21][24], ele[21][25], ele[21][26], ele[21][27], ele[21][28], ele[21][29], ele[21][30], ele[21][31], ele[21][32], ele[21][33], ele[21][34], ele[21][35]);
    $display (ele[22][0], ele[22][1], ele[22][2], ele[22][3], ele[22][4], ele[22][5], ele[22][6], ele[22][7], ele[22][8], ele[22][9], ele[22][10], ele[22][11], ele[22][12], ele[22][13], ele[22][14], ele[22][15], ele[22][16], ele[22][17], ele[22][18], ele[22][19], ele[22][20], ele[22][21], ele[22][22], ele[22][23], ele[22][24], ele[22][25], ele[22][26], ele[22][27], ele[22][28], ele[22][29], ele[22][30], ele[22][31], ele[22][32], ele[22][33], ele[22][34], ele[22][35]);
    $display (ele[23][0], ele[23][1], ele[23][2], ele[23][3], ele[23][4], ele[23][5], ele[23][6], ele[23][7], ele[23][8], ele[23][9], ele[23][10], ele[23][11], ele[23][12], ele[23][13], ele[23][14], ele[23][15], ele[23][16], ele[23][17], ele[23][18], ele[23][19], ele[23][20], ele[23][21], ele[23][22], ele[23][23], ele[23][24], ele[23][25], ele[23][26], ele[23][27], ele[23][28], ele[23][29], ele[23][30], ele[23][31], ele[23][32], ele[23][33], ele[23][34], ele[23][35]);
    $display (ele[24][0], ele[24][1], ele[24][2], ele[24][3], ele[24][4], ele[24][5], ele[24][6], ele[24][7], ele[24][8], ele[24][9], ele[24][10], ele[24][11], ele[24][12], ele[24][13], ele[24][14], ele[24][15], ele[24][16], ele[24][17], ele[24][18], ele[24][19], ele[24][20], ele[24][21], ele[24][22], ele[24][23], ele[24][24], ele[24][25], ele[24][26], ele[24][27], ele[24][28], ele[24][29], ele[24][30], ele[24][31], ele[24][32], ele[24][33], ele[24][34], ele[24][35]);
    $display (ele[25][0], ele[25][1], ele[25][2], ele[25][3], ele[25][4], ele[25][5], ele[25][6], ele[25][7], ele[25][8], ele[25][9], ele[25][10], ele[25][11], ele[25][12], ele[25][13], ele[25][14], ele[25][15], ele[25][16], ele[25][17], ele[25][18], ele[25][19], ele[25][20], ele[25][21], ele[25][22], ele[25][23], ele[25][24], ele[25][25], ele[25][26], ele[25][27], ele[25][28], ele[25][29], ele[25][30], ele[25][31], ele[25][32], ele[25][33], ele[25][34], ele[25][35]);
    $display (ele[26][0], ele[26][1], ele[26][2], ele[26][3], ele[26][4], ele[26][5], ele[26][6], ele[26][7], ele[26][8], ele[26][9], ele[26][10], ele[26][11], ele[26][12], ele[26][13], ele[26][14], ele[26][15], ele[26][16], ele[26][17], ele[26][18], ele[26][19], ele[26][20], ele[26][21], ele[26][22], ele[26][23], ele[26][24], ele[26][25], ele[26][26], ele[26][27], ele[26][28], ele[26][29], ele[26][30], ele[26][31], ele[26][32], ele[26][33], ele[26][34], ele[26][35]);
    $display (ele[27][0], ele[27][1], ele[27][2], ele[27][3], ele[27][4], ele[27][5], ele[27][6], ele[27][7], ele[27][8], ele[27][9], ele[27][10], ele[27][11], ele[27][12], ele[27][13], ele[27][14], ele[27][15], ele[27][16], ele[27][17], ele[27][18], ele[27][19], ele[27][20], ele[27][21], ele[27][22], ele[27][23], ele[27][24], ele[27][25], ele[27][26], ele[27][27], ele[27][28], ele[27][29], ele[27][30], ele[27][31], ele[27][32], ele[27][33], ele[27][34], ele[27][35]);
    $display (ele[28][0], ele[28][1], ele[28][2], ele[28][3], ele[28][4], ele[28][5], ele[28][6], ele[28][7], ele[28][8], ele[28][9], ele[28][10], ele[28][11], ele[28][12], ele[28][13], ele[28][14], ele[28][15], ele[28][16], ele[28][17], ele[28][18], ele[28][19], ele[28][20], ele[28][21], ele[28][22], ele[28][23], ele[28][24], ele[28][25], ele[28][26], ele[28][27], ele[28][28], ele[28][29], ele[28][30], ele[28][31], ele[28][32], ele[28][33], ele[28][34], ele[28][35]);
    $display (ele[29][0], ele[29][1], ele[29][2], ele[29][3], ele[29][4], ele[29][5], ele[29][6], ele[29][7], ele[29][8], ele[29][9], ele[29][10], ele[29][11], ele[29][12], ele[29][13], ele[29][14], ele[29][15], ele[29][16], ele[29][17], ele[29][18], ele[29][19], ele[29][20], ele[29][21], ele[29][22], ele[29][23], ele[29][24], ele[29][25], ele[29][26], ele[29][27], ele[29][28], ele[29][29], ele[29][30], ele[29][31], ele[29][32], ele[29][33], ele[29][34], ele[29][35]);
    $display (ele[30][0], ele[30][1], ele[30][2], ele[30][3], ele[30][4], ele[30][5], ele[30][6], ele[30][7], ele[30][8], ele[30][9], ele[30][10], ele[30][11], ele[30][12], ele[30][13], ele[30][14], ele[30][15], ele[30][16], ele[30][17], ele[30][18], ele[30][19], ele[30][20], ele[30][21], ele[30][22], ele[30][23], ele[30][24], ele[30][25], ele[30][26], ele[30][27], ele[30][28], ele[30][29], ele[30][30], ele[30][31], ele[30][32], ele[30][33], ele[30][34], ele[30][35]);
    $display (ele[31][0], ele[31][1], ele[31][2], ele[31][3], ele[31][4], ele[31][5], ele[31][6], ele[31][7], ele[31][8], ele[31][9], ele[31][10], ele[31][11], ele[31][12], ele[31][13], ele[31][14], ele[31][15], ele[31][16], ele[31][17], ele[31][18], ele[31][19], ele[31][20], ele[31][21], ele[31][22], ele[31][23], ele[31][24], ele[31][25], ele[31][26], ele[31][27], ele[31][28], ele[31][29], ele[31][30], ele[31][31], ele[31][32], ele[31][33], ele[31][34], ele[31][35]);
    $display (ele[32][0], ele[32][1], ele[32][2], ele[32][3], ele[32][4], ele[32][5], ele[32][6], ele[32][7], ele[32][8], ele[32][9], ele[32][10], ele[32][11], ele[32][12], ele[32][13], ele[32][14], ele[32][15], ele[32][16], ele[32][17], ele[32][18], ele[32][19], ele[32][20], ele[32][21], ele[32][22], ele[32][23], ele[32][24], ele[32][25], ele[32][26], ele[32][27], ele[32][28], ele[32][29], ele[32][30], ele[32][31], ele[32][32], ele[32][33], ele[32][34], ele[32][35]);
    $display (ele[33][0], ele[33][1], ele[33][2], ele[33][3], ele[33][4], ele[33][5], ele[33][6], ele[33][7], ele[33][8], ele[33][9], ele[33][10], ele[33][11], ele[33][12], ele[33][13], ele[33][14], ele[33][15], ele[33][16], ele[33][17], ele[33][18], ele[33][19], ele[33][20], ele[33][21], ele[33][22], ele[33][23], ele[33][24], ele[33][25], ele[33][26], ele[33][27], ele[33][28], ele[33][29], ele[33][30], ele[33][31], ele[33][32], ele[33][33], ele[33][34], ele[33][35]);
    $display (ele[34][0], ele[34][1], ele[34][2], ele[34][3], ele[34][4], ele[34][5], ele[34][6], ele[34][7], ele[34][8], ele[34][9], ele[34][10], ele[34][11], ele[34][12], ele[34][13], ele[34][14], ele[34][15], ele[34][16], ele[34][17], ele[34][18], ele[34][19], ele[34][20], ele[34][21], ele[34][22], ele[34][23], ele[34][24], ele[34][25], ele[34][26], ele[34][27], ele[34][28], ele[34][29], ele[34][30], ele[34][31], ele[34][32], ele[34][33], ele[34][34], ele[34][35]);
    $display (ele[35][0], ele[35][1], ele[35][2], ele[35][3], ele[35][4], ele[35][5], ele[35][6], ele[35][7], ele[35][8], ele[35][9], ele[35][10], ele[35][11], ele[35][12], ele[35][13], ele[35][14], ele[35][15], ele[35][16], ele[35][17], ele[35][18], ele[35][19], ele[35][20], ele[35][21], ele[35][22], ele[35][23], ele[35][24], ele[35][25], ele[35][26], ele[35][27], ele[35][28], ele[35][29], ele[35][30], ele[35][31], ele[35][32], ele[35][33], ele[35][34], ele[35][35]);
  endfunction: show
endclass: board
